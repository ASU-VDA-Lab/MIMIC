module fake_netlist_6_3529_n_2822 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_397, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_407, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2822);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_397;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_407;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2822;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_491;
wire n_2786;
wire n_1591;
wire n_772;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_2735;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_483;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_433;
wire n_2546;
wire n_792;
wire n_2522;
wire n_476;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1599;
wire n_1068;
wire n_982;
wire n_2674;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_2455;
wire n_558;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2749;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_690;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2810;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_484;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_462;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_2767;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_644;
wire n_682;
wire n_2537;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_536;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_499;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_526;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_552;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_1774;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1475;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2511;
wire n_537;
wire n_2475;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_1141;
wire n_562;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_426;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_2801;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_463;
wire n_1243;
wire n_848;
wire n_2732;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_2627;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2781;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_419;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_2420;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_2756;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1669;
wire n_1403;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_2052;
wire n_1847;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_621;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_2755;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2819;
wire n_466;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_2439;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_1601;
wire n_609;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_1352;
wire n_579;
wire n_2789;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_456;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_654;
wire n_411;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_482;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_420;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_2798;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_523;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_1650;
wire n_706;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2793;
wire n_2715;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_2076;
wire n_2736;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_761;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_611;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_445;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_2265;
wire n_2615;
wire n_414;
wire n_2683;
wire n_1922;
wire n_563;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_2743;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_455;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_2600;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_436;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_2285;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2795;
wire n_2471;
wire n_467;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_1629;
wire n_665;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_2774;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_1322;
wire n_640;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_422;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_396),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_278),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_29),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_92),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_25),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_348),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_371),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_135),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_357),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_183),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_113),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_282),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_8),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_317),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_99),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_323),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_245),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_76),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_244),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_308),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_187),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_195),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_201),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_141),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_235),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_297),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_307),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_123),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_170),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_387),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_128),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_385),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_363),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_82),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_98),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_3),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_285),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_362),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_133),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_279),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_390),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_79),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_130),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_41),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_11),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_15),
.Y(n_455)
);

CKINVDCx14_ASAP7_75t_R g456 ( 
.A(n_231),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_326),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_194),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_78),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_68),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_135),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_331),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_162),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_222),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_281),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_224),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_128),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_378),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_178),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_209),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_157),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_346),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_334),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_333),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_401),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_397),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_19),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_133),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_17),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_263),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_395),
.Y(n_481)
);

BUFx10_ASAP7_75t_L g482 ( 
.A(n_194),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_316),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_306),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_175),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_118),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_188),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_187),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_403),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_312),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_375),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_303),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_167),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_77),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_149),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_199),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_175),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_383),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_264),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_15),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_234),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_343),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_6),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_382),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_27),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_73),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_238),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_81),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_280),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_219),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_70),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_259),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_122),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_246),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_206),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_18),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_95),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_322),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_2),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_49),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_77),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_406),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_223),
.Y(n_523)
);

BUFx8_ASAP7_75t_SL g524 ( 
.A(n_370),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_274),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_112),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_319),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_389),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_353),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_376),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_388),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_65),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_182),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_167),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_399),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_171),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_95),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_394),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_107),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_161),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_145),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_138),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_342),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_125),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_247),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_85),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_153),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_222),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_20),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_339),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_329),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_261),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_155),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_253),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_176),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_294),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_404),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_236),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_29),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_402),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_196),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_212),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_295),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_283),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_391),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_367),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_359),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_407),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_204),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_239),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_1),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_200),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_366),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_225),
.Y(n_574)
);

INVxp67_ASAP7_75t_SL g575 ( 
.A(n_33),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_193),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_286),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_289),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_17),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_168),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_233),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_188),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_405),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_381),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_63),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_384),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_81),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_195),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_44),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_266),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_328),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_54),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_229),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_356),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_210),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_327),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_214),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_9),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_273),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_386),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_372),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_393),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_50),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_231),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_337),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_218),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_309),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_89),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_227),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_110),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_52),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_205),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_25),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_138),
.Y(n_614)
);

BUFx5_ASAP7_75t_L g615 ( 
.A(n_8),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_75),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_216),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_59),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_364),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_98),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_127),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_229),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_16),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_377),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_409),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_321),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_132),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_101),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g629 ( 
.A(n_73),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_250),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_227),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_50),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_80),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_37),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_144),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_139),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_265),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_290),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_111),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_45),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_180),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_109),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_207),
.Y(n_643)
);

INVxp33_ASAP7_75t_R g644 ( 
.A(n_392),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_23),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_68),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_180),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_172),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_9),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_46),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_400),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_116),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_269),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_166),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_96),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_66),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_76),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_215),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_80),
.Y(n_659)
);

BUFx10_ASAP7_75t_L g660 ( 
.A(n_60),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_373),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_212),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_142),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_33),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_132),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_197),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_164),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_254),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_26),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_3),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_96),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_0),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_55),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_325),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_369),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_6),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_152),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_161),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_240),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_0),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_352),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_361),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_237),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_398),
.Y(n_684)
);

BUFx8_ASAP7_75t_SL g685 ( 
.A(n_284),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_7),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_173),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_214),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_248),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_160),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_311),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_305),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_75),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_215),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_69),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_318),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_324),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_344),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_19),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_210),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_276),
.Y(n_701)
);

CKINVDCx14_ASAP7_75t_R g702 ( 
.A(n_191),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_97),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_230),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_131),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_252),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_97),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_408),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_144),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_213),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_163),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_186),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_65),
.Y(n_713)
);

CKINVDCx14_ASAP7_75t_R g714 ( 
.A(n_314),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_90),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_302),
.Y(n_716)
);

BUFx5_ASAP7_75t_L g717 ( 
.A(n_332),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_615),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_456),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_615),
.Y(n_720)
);

INVxp67_ASAP7_75t_SL g721 ( 
.A(n_480),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_615),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_615),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_702),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_418),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_437),
.Y(n_726)
);

BUFx6f_ASAP7_75t_SL g727 ( 
.A(n_556),
.Y(n_727)
);

INVxp67_ASAP7_75t_SL g728 ( 
.A(n_462),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_615),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_615),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_553),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_425),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_412),
.Y(n_733)
);

CKINVDCx16_ASAP7_75t_R g734 ( 
.A(n_551),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_615),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_615),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_491),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_615),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_415),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_553),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_415),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_537),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_426),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_426),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_528),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_419),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_436),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_R g748 ( 
.A(n_714),
.B(n_232),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_436),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_442),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_437),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_422),
.Y(n_752)
);

CKINVDCx16_ASAP7_75t_R g753 ( 
.A(n_551),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_430),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_568),
.Y(n_755)
);

INVxp33_ASAP7_75t_L g756 ( 
.A(n_559),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_601),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_431),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_691),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_442),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_457),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_457),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_432),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_472),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_472),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_438),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_413),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_476),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_462),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_476),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_440),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_481),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_481),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_499),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_443),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_499),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_444),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_501),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_445),
.Y(n_779)
);

INVxp33_ASAP7_75t_SL g780 ( 
.A(n_670),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_451),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_453),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_524),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_417),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_552),
.B(n_1),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_437),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_437),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_501),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_552),
.B(n_2),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_512),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_512),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_577),
.B(n_596),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_461),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_463),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_464),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_530),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_685),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_530),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_437),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_538),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_466),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_538),
.Y(n_802)
);

NOR2xp67_ASAP7_75t_L g803 ( 
.A(n_653),
.B(n_4),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_410),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_560),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_560),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_470),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_564),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_413),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_564),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_471),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_577),
.B(n_4),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_411),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_477),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_416),
.Y(n_815)
);

NOR2xp67_ASAP7_75t_L g816 ( 
.A(n_653),
.B(n_5),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_479),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_485),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_566),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_487),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_566),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_421),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_423),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_496),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_584),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_429),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_584),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_417),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_434),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_435),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_602),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_420),
.B(n_5),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_439),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_602),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_441),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_500),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_420),
.Y(n_837)
);

CKINVDCx20_ASAP7_75t_R g838 ( 
.A(n_446),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_619),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_447),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_619),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_668),
.Y(n_842)
);

INVxp33_ASAP7_75t_SL g843 ( 
.A(n_505),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_668),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_511),
.Y(n_845)
);

CKINVDCx16_ASAP7_75t_R g846 ( 
.A(n_482),
.Y(n_846)
);

CKINVDCx16_ASAP7_75t_R g847 ( 
.A(n_482),
.Y(n_847)
);

BUFx2_ASAP7_75t_L g848 ( 
.A(n_413),
.Y(n_848)
);

CKINVDCx16_ASAP7_75t_R g849 ( 
.A(n_482),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_449),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_596),
.B(n_570),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_513),
.Y(n_852)
);

CKINVDCx16_ASAP7_75t_R g853 ( 
.A(n_482),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_517),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_437),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_478),
.Y(n_856)
);

AND2x6_ASAP7_75t_L g857 ( 
.A(n_718),
.B(n_653),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_751),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_851),
.B(n_539),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_751),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_733),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_803),
.B(n_556),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_804),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_813),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_726),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_815),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_822),
.Y(n_867)
);

AND2x6_ASAP7_75t_L g868 ( 
.A(n_718),
.B(n_653),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_786),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_786),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_787),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_855),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_725),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_767),
.B(n_539),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_855),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_856),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_823),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_792),
.B(n_567),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_767),
.B(n_539),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_787),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_826),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_829),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_732),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_733),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_799),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_856),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_746),
.Y(n_887)
);

CKINVDCx16_ASAP7_75t_R g888 ( 
.A(n_734),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_737),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_739),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_721),
.B(n_809),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_746),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_799),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_741),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_830),
.Y(n_895)
);

NAND2xp33_ASAP7_75t_SL g896 ( 
.A(n_719),
.B(n_459),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_809),
.B(n_576),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_816),
.B(n_556),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_R g899 ( 
.A(n_783),
.B(n_465),
.Y(n_899)
);

CKINVDCx16_ASAP7_75t_R g900 ( 
.A(n_753),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_726),
.B(n_605),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_728),
.B(n_567),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_848),
.B(n_769),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_743),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_744),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_747),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_726),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_843),
.B(n_570),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_833),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_752),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_848),
.B(n_605),
.Y(n_911)
);

AND2x6_ASAP7_75t_L g912 ( 
.A(n_720),
.B(n_428),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_720),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_749),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_722),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_745),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_750),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_835),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_723),
.B(n_605),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_760),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_807),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_761),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_740),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_755),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_727),
.Y(n_925)
);

NAND2x1p5_ASAP7_75t_L g926 ( 
.A(n_785),
.B(n_450),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_729),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_730),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_762),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_735),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_784),
.B(n_576),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_764),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_765),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_757),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_768),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_736),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_828),
.B(n_576),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_770),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_R g939 ( 
.A(n_797),
.B(n_468),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_772),
.B(n_630),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_773),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_738),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_838),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_774),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_759),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_837),
.B(n_776),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_843),
.B(n_630),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_719),
.B(n_473),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_778),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_788),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_840),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_850),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_724),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_724),
.B(n_474),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_752),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_790),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_791),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_796),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_798),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_800),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_754),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_802),
.Y(n_962)
);

NAND2x1p5_ASAP7_75t_L g963 ( 
.A(n_789),
.B(n_514),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_805),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_806),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_754),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_808),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_810),
.B(n_819),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_758),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_846),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_758),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_821),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_825),
.A2(n_535),
.B(n_527),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_827),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_831),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_763),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_834),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_839),
.B(n_527),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_847),
.B(n_478),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_763),
.Y(n_980)
);

INVx4_ASAP7_75t_L g981 ( 
.A(n_930),
.Y(n_981)
);

OAI21xp33_ASAP7_75t_L g982 ( 
.A1(n_878),
.A2(n_812),
.B(n_780),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_870),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_890),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_894),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_869),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_899),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_869),
.Y(n_988)
);

INVx4_ASAP7_75t_L g989 ( 
.A(n_930),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_862),
.B(n_841),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_904),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_905),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_906),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_911),
.B(n_849),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_901),
.B(n_842),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_870),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_862),
.B(n_898),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_914),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_930),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_930),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_930),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_880),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_901),
.B(n_844),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_939),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_870),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_870),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_862),
.B(n_766),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_902),
.B(n_527),
.Y(n_1008)
);

BUFx10_ASAP7_75t_L g1009 ( 
.A(n_953),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_917),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_898),
.B(n_766),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_951),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_920),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_857),
.A2(n_832),
.B1(n_424),
.B2(n_593),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_898),
.B(n_908),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_903),
.B(n_853),
.Y(n_1016)
);

INVx5_ASAP7_75t_L g1017 ( 
.A(n_912),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_901),
.B(n_696),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_880),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_929),
.Y(n_1020)
);

INVx5_ASAP7_75t_L g1021 ( 
.A(n_912),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_932),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_933),
.Y(n_1023)
);

OR2x6_ASAP7_75t_L g1024 ( 
.A(n_961),
.B(n_644),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_922),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_970),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_935),
.Y(n_1027)
);

INVxp67_ASAP7_75t_SL g1028 ( 
.A(n_968),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_870),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_885),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_938),
.Y(n_1031)
);

OR2x2_ASAP7_75t_SL g1032 ( 
.A(n_888),
.B(n_832),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_947),
.B(n_771),
.Y(n_1033)
);

OR2x6_ASAP7_75t_L g1034 ( 
.A(n_884),
.B(n_644),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_941),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_871),
.Y(n_1036)
);

CKINVDCx14_ASAP7_75t_R g1037 ( 
.A(n_970),
.Y(n_1037)
);

AND2x6_ASAP7_75t_L g1038 ( 
.A(n_859),
.B(n_535),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_953),
.Y(n_1039)
);

INVx5_ASAP7_75t_L g1040 ( 
.A(n_912),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_950),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_942),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_885),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_865),
.B(n_771),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_926),
.B(n_535),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_865),
.B(n_915),
.Y(n_1046)
);

INVxp67_ASAP7_75t_SL g1047 ( 
.A(n_919),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_921),
.A2(n_780),
.B1(n_775),
.B2(n_779),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_874),
.Y(n_1049)
);

NOR3xp33_ASAP7_75t_L g1050 ( 
.A(n_923),
.B(n_900),
.C(n_979),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_874),
.B(n_775),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_863),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_913),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_863),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_879),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_942),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_865),
.B(n_777),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_926),
.B(n_581),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_940),
.B(n_696),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_955),
.Y(n_1060)
);

INVx5_ASAP7_75t_L g1061 ( 
.A(n_912),
.Y(n_1061)
);

INVx4_ASAP7_75t_L g1062 ( 
.A(n_942),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_956),
.Y(n_1063)
);

INVx5_ASAP7_75t_L g1064 ( 
.A(n_912),
.Y(n_1064)
);

INVxp67_ASAP7_75t_SL g1065 ( 
.A(n_913),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_957),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_958),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_942),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_942),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_871),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_962),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_940),
.B(n_922),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_857),
.A2(n_424),
.B1(n_593),
.B2(n_494),
.Y(n_1073)
);

INVx4_ASAP7_75t_L g1074 ( 
.A(n_944),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_964),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_963),
.B(n_581),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_891),
.B(n_777),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_907),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_915),
.B(n_779),
.Y(n_1079)
);

AND2x6_ASAP7_75t_L g1080 ( 
.A(n_859),
.B(n_581),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_944),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_896),
.A2(n_781),
.B1(n_793),
.B2(n_782),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_944),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_857),
.A2(n_424),
.B1(n_593),
.B2(n_494),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_965),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_SL g1086 ( 
.A(n_925),
.B(n_455),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_955),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_871),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_927),
.B(n_781),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_967),
.Y(n_1090)
);

AND2x6_ASAP7_75t_L g1091 ( 
.A(n_940),
.B(n_675),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_944),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_972),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_927),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_978),
.B(n_697),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_871),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_928),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_907),
.Y(n_1098)
);

OR2x6_ASAP7_75t_L g1099 ( 
.A(n_887),
.B(n_731),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_948),
.B(n_782),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_871),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_954),
.B(n_793),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_963),
.B(n_794),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_928),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_893),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_936),
.B(n_794),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_978),
.B(n_675),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_944),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_879),
.B(n_795),
.Y(n_1109)
);

INVx4_ASAP7_75t_SL g1110 ( 
.A(n_857),
.Y(n_1110)
);

BUFx4f_ASAP7_75t_L g1111 ( 
.A(n_892),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_864),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_936),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_858),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_860),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_872),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_864),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_978),
.B(n_675),
.Y(n_1118)
);

AO22x2_ASAP7_75t_L g1119 ( 
.A1(n_897),
.A2(n_510),
.B1(n_606),
.B2(n_459),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_875),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_946),
.B(n_428),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_876),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_886),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_949),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_857),
.B(n_868),
.Y(n_1125)
);

INVx8_ASAP7_75t_L g1126 ( 
.A(n_966),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_857),
.B(n_795),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_949),
.Y(n_1128)
);

AO22x2_ASAP7_75t_L g1129 ( 
.A1(n_897),
.A2(n_510),
.B1(n_606),
.B2(n_494),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_931),
.Y(n_1130)
);

OR2x2_ASAP7_75t_L g1131 ( 
.A(n_931),
.B(n_801),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_949),
.B(n_801),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_959),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_946),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_893),
.Y(n_1135)
);

BUFx4f_ASAP7_75t_L g1136 ( 
.A(n_910),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_937),
.B(n_811),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_937),
.B(n_811),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_893),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_959),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_960),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_868),
.B(n_814),
.Y(n_1142)
);

INVx1_ASAP7_75t_SL g1143 ( 
.A(n_951),
.Y(n_1143)
);

OR2x2_ASAP7_75t_L g1144 ( 
.A(n_861),
.B(n_814),
.Y(n_1144)
);

INVxp67_ASAP7_75t_SL g1145 ( 
.A(n_973),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_866),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_960),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_868),
.B(n_817),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_974),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_973),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_982),
.B(n_966),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_1025),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1047),
.B(n_868),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1047),
.B(n_868),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1015),
.B(n_969),
.Y(n_1155)
);

NOR2x2_ASAP7_75t_L g1156 ( 
.A(n_1034),
.B(n_617),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1053),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1028),
.B(n_969),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1008),
.A2(n_868),
.B1(n_623),
.B2(n_648),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_984),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1028),
.B(n_817),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_997),
.B(n_1065),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_985),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_991),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_1099),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_992),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_993),
.Y(n_1167)
);

NAND2x1p5_ASAP7_75t_L g1168 ( 
.A(n_1134),
.B(n_697),
.Y(n_1168)
);

NOR2xp67_ASAP7_75t_L g1169 ( 
.A(n_987),
.B(n_1004),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1077),
.B(n_971),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1014),
.B(n_980),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1077),
.B(n_971),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1065),
.B(n_818),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1014),
.B(n_976),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1145),
.A2(n_912),
.B(n_708),
.Y(n_1175)
);

AND2x6_ASAP7_75t_SL g1176 ( 
.A(n_1034),
.B(n_427),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1053),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1131),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_995),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_998),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1073),
.B(n_980),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1130),
.B(n_976),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_995),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1073),
.B(n_428),
.Y(n_1184)
);

AND2x6_ASAP7_75t_L g1185 ( 
.A(n_1150),
.B(n_1125),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1010),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1008),
.A2(n_623),
.B1(n_648),
.B2(n_617),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1084),
.B(n_428),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1100),
.B(n_818),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1078),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_1025),
.Y(n_1191)
);

INVx4_ASAP7_75t_L g1192 ( 
.A(n_999),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1013),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_995),
.B(n_974),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1046),
.A2(n_977),
.B(n_975),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_1003),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1100),
.B(n_820),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1102),
.B(n_820),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1049),
.B(n_824),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_986),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1102),
.B(n_824),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1038),
.A2(n_623),
.B1(n_648),
.B2(n_617),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1132),
.B(n_836),
.Y(n_1203)
);

NAND2x1_ASAP7_75t_L g1204 ( 
.A(n_983),
.B(n_925),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1078),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1132),
.B(n_836),
.Y(n_1206)
);

INVxp33_ASAP7_75t_L g1207 ( 
.A(n_1109),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1033),
.A2(n_708),
.B(n_701),
.C(n_975),
.Y(n_1208)
);

INVxp67_ASAP7_75t_L g1209 ( 
.A(n_1109),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1038),
.A2(n_672),
.B1(n_703),
.B2(n_666),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1055),
.B(n_1051),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1137),
.A2(n_845),
.B1(n_854),
.B2(n_852),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1038),
.A2(n_672),
.B1(n_703),
.B2(n_666),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1113),
.B(n_845),
.Y(n_1214)
);

INVxp33_ASAP7_75t_SL g1215 ( 
.A(n_987),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1020),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1084),
.B(n_1134),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1127),
.B(n_1142),
.Y(n_1218)
);

NOR3xp33_ASAP7_75t_L g1219 ( 
.A(n_1033),
.B(n_883),
.C(n_867),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1148),
.B(n_428),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1003),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1072),
.B(n_428),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1113),
.B(n_852),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1003),
.B(n_854),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1137),
.B(n_742),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1138),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1124),
.B(n_977),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1016),
.B(n_756),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1022),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1111),
.B(n_866),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1044),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1079),
.B(n_414),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1089),
.B(n_460),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1128),
.B(n_925),
.Y(n_1234)
);

OR2x6_ASAP7_75t_L g1235 ( 
.A(n_1034),
.B(n_664),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1057),
.A2(n_701),
.B(n_692),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_990),
.B(n_748),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_SL g1238 ( 
.A(n_1004),
.B(n_867),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1106),
.B(n_486),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1038),
.B(n_475),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1150),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_994),
.Y(n_1242)
);

NAND2xp33_ASAP7_75t_L g1243 ( 
.A(n_1038),
.B(n_717),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1072),
.B(n_1110),
.Y(n_1244)
);

O2A1O1Ixp5_ASAP7_75t_L g1245 ( 
.A1(n_1145),
.A2(n_1121),
.B(n_1045),
.C(n_1076),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1098),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1023),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1099),
.B(n_877),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1080),
.A2(n_672),
.B1(n_703),
.B2(n_666),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1072),
.B(n_489),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1103),
.A2(n_483),
.B1(n_490),
.B2(n_484),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1027),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1099),
.B(n_877),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1080),
.A2(n_433),
.B1(n_448),
.B2(n_427),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1098),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1110),
.B(n_489),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1007),
.B(n_488),
.Y(n_1257)
);

AND2x6_ASAP7_75t_SL g1258 ( 
.A(n_1024),
.B(n_433),
.Y(n_1258)
);

BUFx8_ASAP7_75t_L g1259 ( 
.A(n_1026),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1111),
.B(n_881),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1011),
.B(n_497),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1110),
.B(n_489),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1080),
.B(n_492),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1080),
.B(n_498),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_986),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1017),
.B(n_1021),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1031),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1035),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_988),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1032),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_1144),
.B(n_881),
.Y(n_1271)
);

NOR2x1p5_ASAP7_75t_L g1272 ( 
.A(n_1052),
.B(n_882),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_SL g1273 ( 
.A(n_1017),
.B(n_489),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1041),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_988),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1080),
.B(n_502),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1002),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1063),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1066),
.Y(n_1279)
);

INVx2_ASAP7_75t_SL g1280 ( 
.A(n_1059),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1129),
.A2(n_452),
.B1(n_454),
.B2(n_448),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1067),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_999),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1071),
.Y(n_1284)
);

AO22x1_ASAP7_75t_L g1285 ( 
.A1(n_1103),
.A2(n_575),
.B1(n_454),
.B2(n_458),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1075),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1086),
.A2(n_895),
.B1(n_909),
.B2(n_882),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_1060),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1085),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1059),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1090),
.Y(n_1291)
);

NAND2xp33_ASAP7_75t_L g1292 ( 
.A(n_1091),
.B(n_717),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1129),
.A2(n_458),
.B1(n_469),
.B2(n_452),
.Y(n_1293)
);

INVx2_ASAP7_75t_SL g1294 ( 
.A(n_1059),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_SL g1295 ( 
.A(n_1136),
.B(n_895),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1114),
.B(n_504),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1115),
.B(n_507),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1017),
.B(n_489),
.Y(n_1298)
);

NAND2x1p5_ASAP7_75t_L g1299 ( 
.A(n_1017),
.B(n_1021),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_999),
.Y(n_1300)
);

OR2x6_ASAP7_75t_L g1301 ( 
.A(n_1126),
.B(n_664),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1093),
.Y(n_1302)
);

AND3x1_ASAP7_75t_L g1303 ( 
.A(n_1050),
.B(n_1048),
.C(n_1082),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1045),
.B(n_613),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1129),
.A2(n_469),
.B1(n_503),
.B2(n_495),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1116),
.B(n_509),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1021),
.B(n_489),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1122),
.B(n_518),
.Y(n_1308)
);

INVx5_ASAP7_75t_L g1309 ( 
.A(n_1091),
.Y(n_1309)
);

NAND2xp33_ASAP7_75t_L g1310 ( 
.A(n_1091),
.B(n_717),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1021),
.B(n_554),
.Y(n_1311)
);

NOR2xp67_ASAP7_75t_SL g1312 ( 
.A(n_1040),
.B(n_554),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1133),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1136),
.B(n_1087),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1002),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1040),
.B(n_554),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1140),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1141),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1147),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1058),
.A2(n_525),
.B1(n_529),
.B2(n_522),
.Y(n_1320)
);

OAI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1058),
.A2(n_634),
.B1(n_546),
.B2(n_664),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1019),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1019),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1076),
.A2(n_543),
.B1(n_545),
.B2(n_531),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1018),
.B(n_550),
.Y(n_1325)
);

AOI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1018),
.A2(n_558),
.B1(n_563),
.B2(n_557),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1018),
.B(n_565),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1091),
.A2(n_578),
.B1(n_583),
.B2(n_573),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1095),
.B(n_713),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1091),
.A2(n_590),
.B1(n_591),
.B2(n_586),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1120),
.B(n_1123),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1149),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1120),
.B(n_594),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1040),
.B(n_554),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1123),
.B(n_599),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1039),
.B(n_909),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1094),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1097),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1030),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1052),
.Y(n_1340)
);

NOR2xp67_ASAP7_75t_L g1341 ( 
.A(n_1054),
.B(n_918),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1121),
.B(n_600),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1095),
.A2(n_624),
.B1(n_625),
.B2(n_607),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1040),
.B(n_554),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1012),
.B(n_1143),
.Y(n_1345)
);

INVx4_ASAP7_75t_L g1346 ( 
.A(n_999),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1095),
.A2(n_637),
.B1(n_638),
.B2(n_626),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1162),
.B(n_1104),
.Y(n_1348)
);

O2A1O1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1217),
.A2(n_1118),
.B(n_1107),
.C(n_1043),
.Y(n_1349)
);

A2O1A1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1170),
.A2(n_503),
.B(n_508),
.C(n_495),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1155),
.B(n_1108),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1215),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1217),
.A2(n_1158),
.B1(n_1174),
.B2(n_1171),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1225),
.B(n_1009),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1225),
.B(n_1009),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1152),
.B(n_1108),
.Y(n_1356)
);

A2O1A1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1170),
.A2(n_516),
.B(n_520),
.C(n_508),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1155),
.B(n_1119),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_1283),
.Y(n_1359)
);

OR2x6_ASAP7_75t_L g1360 ( 
.A(n_1165),
.B(n_1126),
.Y(n_1360)
);

NOR3xp33_ASAP7_75t_SL g1361 ( 
.A(n_1158),
.B(n_1112),
.C(n_1054),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_SL g1362 ( 
.A(n_1172),
.B(n_1117),
.C(n_1112),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1232),
.B(n_1233),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1231),
.A2(n_1118),
.B1(n_1107),
.B2(n_943),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1177),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1345),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1211),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1232),
.B(n_1119),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_SL g1369 ( 
.A1(n_1172),
.A2(n_889),
.B1(n_916),
.B2(n_873),
.Y(n_1369)
);

INVx6_ASAP7_75t_L g1370 ( 
.A(n_1259),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1340),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1207),
.B(n_1126),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1233),
.B(n_1119),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1209),
.B(n_918),
.Y(n_1374)
);

BUFx4f_ASAP7_75t_L g1375 ( 
.A(n_1248),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1331),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1194),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1194),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1336),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1270),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1259),
.Y(n_1381)
);

A2O1A1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1304),
.A2(n_1151),
.B(n_1239),
.C(n_1257),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1309),
.B(n_1061),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1177),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1184),
.A2(n_713),
.B1(n_520),
.B2(n_526),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1283),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1200),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1152),
.B(n_1024),
.Y(n_1388)
);

INVx5_ASAP7_75t_L g1389 ( 
.A(n_1185),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1283),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1191),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1171),
.A2(n_952),
.B1(n_943),
.B2(n_1135),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1239),
.B(n_983),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1200),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1309),
.B(n_1061),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1199),
.Y(n_1396)
);

AOI22x1_ASAP7_75t_L g1397 ( 
.A1(n_1175),
.A2(n_1139),
.B1(n_1135),
.B2(n_1005),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1265),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1161),
.B(n_1203),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1265),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1191),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1275),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1288),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1196),
.B(n_1024),
.Y(n_1404)
);

INVx8_ASAP7_75t_L g1405 ( 
.A(n_1301),
.Y(n_1405)
);

INVxp67_ASAP7_75t_SL g1406 ( 
.A(n_1241),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1275),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1160),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1189),
.B(n_952),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1163),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1164),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1166),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1167),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1283),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1180),
.Y(n_1415)
);

NOR3xp33_ASAP7_75t_SL g1416 ( 
.A(n_1151),
.B(n_1146),
.C(n_1117),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1196),
.B(n_1139),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1206),
.B(n_996),
.Y(n_1418)
);

INVxp67_ASAP7_75t_SL g1419 ( 
.A(n_1241),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1186),
.Y(n_1420)
);

BUFx4f_ASAP7_75t_L g1421 ( 
.A(n_1253),
.Y(n_1421)
);

NAND2xp33_ASAP7_75t_SL g1422 ( 
.A(n_1314),
.B(n_1146),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1193),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1287),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1216),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1157),
.Y(n_1426)
);

INVxp33_ASAP7_75t_L g1427 ( 
.A(n_1228),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1221),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1257),
.B(n_996),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1221),
.B(n_873),
.Y(n_1430)
);

CKINVDCx16_ASAP7_75t_R g1431 ( 
.A(n_1238),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1269),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1261),
.B(n_1005),
.Y(n_1433)
);

BUFx12f_ASAP7_75t_L g1434 ( 
.A(n_1176),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1229),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1277),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1247),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1179),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1280),
.B(n_889),
.Y(n_1439)
);

BUFx12f_ASAP7_75t_L g1440 ( 
.A(n_1258),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1252),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1261),
.B(n_1006),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1226),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1267),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1268),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1230),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1184),
.A2(n_713),
.B1(n_526),
.B2(n_534),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1228),
.B(n_1037),
.Y(n_1448)
);

AOI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1174),
.A2(n_1074),
.B1(n_989),
.B2(n_1001),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1315),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1304),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1260),
.Y(n_1452)
);

INVx5_ASAP7_75t_L g1453 ( 
.A(n_1185),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1173),
.B(n_1006),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1274),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1278),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1279),
.Y(n_1457)
);

BUFx4f_ASAP7_75t_L g1458 ( 
.A(n_1301),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1179),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1290),
.B(n_916),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1212),
.Y(n_1461)
);

INVx4_ASAP7_75t_L g1462 ( 
.A(n_1183),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1156),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1329),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1271),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1183),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1329),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1178),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1197),
.B(n_467),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1182),
.B(n_1037),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1182),
.B(n_924),
.Y(n_1471)
);

AND2x6_ASAP7_75t_L g1472 ( 
.A(n_1153),
.B(n_554),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1282),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1300),
.Y(n_1474)
);

INVx4_ASAP7_75t_L g1475 ( 
.A(n_1300),
.Y(n_1475)
);

NOR3xp33_ASAP7_75t_SL g1476 ( 
.A(n_1321),
.B(n_521),
.C(n_519),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1242),
.B(n_924),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1294),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1284),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1198),
.B(n_1029),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1201),
.B(n_1029),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1235),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1322),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1188),
.A2(n_1187),
.B1(n_1210),
.B2(n_1202),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1235),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1168),
.Y(n_1486)
);

NAND3xp33_ASAP7_75t_SL g1487 ( 
.A(n_1219),
.B(n_945),
.C(n_934),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1309),
.B(n_1061),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1272),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1181),
.A2(n_1074),
.B1(n_989),
.B2(n_1001),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1169),
.B(n_934),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1237),
.B(n_1036),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1286),
.B(n_1036),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1181),
.A2(n_981),
.B1(n_1062),
.B2(n_1042),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1289),
.B(n_945),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1291),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1214),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1302),
.B(n_1070),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_R g1499 ( 
.A(n_1295),
.B(n_493),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1227),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1382),
.A2(n_1210),
.B(n_1213),
.C(n_1202),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1397),
.A2(n_1245),
.B(n_1218),
.Y(n_1502)
);

A2O1A1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1382),
.A2(n_1249),
.B(n_1213),
.C(n_1254),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1363),
.B(n_1223),
.Y(n_1504)
);

AO21x1_ASAP7_75t_L g1505 ( 
.A1(n_1353),
.A2(n_1220),
.B(n_1218),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1349),
.A2(n_1220),
.B(n_1195),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1371),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1365),
.A2(n_1339),
.B(n_1323),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1365),
.A2(n_1205),
.B(n_1190),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1399),
.B(n_1285),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1408),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1354),
.B(n_1341),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1451),
.B(n_1168),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1451),
.B(n_1281),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1367),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1410),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1348),
.A2(n_1309),
.B(n_1154),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1355),
.B(n_1224),
.Y(n_1518)
);

AO31x2_ASAP7_75t_L g1519 ( 
.A1(n_1350),
.A2(n_1208),
.A3(n_1236),
.B(n_1313),
.Y(n_1519)
);

NAND2x1p5_ASAP7_75t_L g1520 ( 
.A(n_1462),
.B(n_1244),
.Y(n_1520)
);

INVx5_ASAP7_75t_L g1521 ( 
.A(n_1359),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1376),
.B(n_1281),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1402),
.A2(n_1492),
.B(n_1418),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1427),
.B(n_1303),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1497),
.B(n_1249),
.Y(n_1525)
);

BUFx12f_ASAP7_75t_L g1526 ( 
.A(n_1370),
.Y(n_1526)
);

AO31x2_ASAP7_75t_L g1527 ( 
.A1(n_1350),
.A2(n_1357),
.A3(n_1358),
.B(n_1368),
.Y(n_1527)
);

OAI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1469),
.A2(n_1235),
.B1(n_1301),
.B2(n_1251),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1402),
.A2(n_1255),
.B(n_1246),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_SL g1530 ( 
.A1(n_1469),
.A2(n_1254),
.B(n_1293),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1406),
.A2(n_1346),
.B(n_1192),
.Y(n_1531)
);

AOI211x1_ASAP7_75t_L g1532 ( 
.A1(n_1373),
.A2(n_1222),
.B(n_1250),
.C(n_1188),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1411),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1406),
.A2(n_1346),
.B(n_1192),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1500),
.B(n_1293),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1430),
.Y(n_1536)
);

O2A1O1Ixp5_ASAP7_75t_L g1537 ( 
.A1(n_1351),
.A2(n_1222),
.B(n_1250),
.C(n_1240),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1484),
.A2(n_1244),
.B1(n_1327),
.B2(n_1325),
.Y(n_1538)
);

AOI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1429),
.A2(n_1264),
.B(n_1263),
.Y(n_1539)
);

OAI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1484),
.A2(n_1185),
.B(n_1276),
.Y(n_1540)
);

AOI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1419),
.A2(n_1454),
.B(n_1299),
.Y(n_1541)
);

AO21x2_ASAP7_75t_L g1542 ( 
.A1(n_1480),
.A2(n_1243),
.B(n_1342),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1449),
.A2(n_1204),
.B(n_1256),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1490),
.A2(n_1262),
.B(n_1256),
.Y(n_1544)
);

A2O1A1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1357),
.A2(n_1305),
.B(n_1187),
.C(n_1159),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1419),
.A2(n_1299),
.B(n_1300),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1384),
.A2(n_1318),
.B(n_1317),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1494),
.A2(n_1262),
.B(n_1319),
.Y(n_1548)
);

OAI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1393),
.A2(n_1185),
.B(n_1159),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1481),
.A2(n_1300),
.B(n_1266),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1387),
.A2(n_1337),
.B(n_1332),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1409),
.B(n_1305),
.Y(n_1552)
);

AO31x2_ASAP7_75t_L g1553 ( 
.A1(n_1433),
.A2(n_1338),
.A3(n_1324),
.B(n_1320),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1439),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1409),
.B(n_1296),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1412),
.B(n_1297),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1394),
.A2(n_1234),
.B(n_1088),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1383),
.A2(n_1266),
.B(n_1042),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1413),
.B(n_1306),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1477),
.B(n_1308),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1398),
.A2(n_1088),
.B(n_1070),
.Y(n_1561)
);

AND2x2_ASAP7_75t_SL g1562 ( 
.A(n_1458),
.B(n_1292),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1400),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1383),
.A2(n_1062),
.B(n_981),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1395),
.A2(n_1488),
.B(n_1442),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1407),
.A2(n_1101),
.B(n_1096),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1395),
.A2(n_1310),
.B(n_1064),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1415),
.B(n_1420),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1488),
.A2(n_1064),
.B(n_1061),
.Y(n_1569)
);

AO31x2_ASAP7_75t_L g1570 ( 
.A1(n_1426),
.A2(n_1335),
.A3(n_1333),
.B(n_1043),
.Y(n_1570)
);

CKINVDCx11_ASAP7_75t_R g1571 ( 
.A(n_1434),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1459),
.B(n_1326),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1430),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_SL g1574 ( 
.A1(n_1486),
.A2(n_1056),
.B(n_1000),
.Y(n_1574)
);

AO31x2_ASAP7_75t_L g1575 ( 
.A1(n_1426),
.A2(n_1030),
.A3(n_534),
.B(n_542),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1423),
.Y(n_1576)
);

AO31x2_ASAP7_75t_L g1577 ( 
.A1(n_1432),
.A2(n_542),
.A3(n_571),
.B(n_516),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1493),
.A2(n_1498),
.B(n_1436),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1425),
.B(n_1185),
.Y(n_1579)
);

AOI21x1_ASAP7_75t_SL g1580 ( 
.A1(n_1417),
.A2(n_1330),
.B(n_1328),
.Y(n_1580)
);

OR2x6_ASAP7_75t_L g1581 ( 
.A(n_1405),
.B(n_1273),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1435),
.B(n_1343),
.Y(n_1582)
);

OAI21x1_ASAP7_75t_L g1583 ( 
.A1(n_1432),
.A2(n_1101),
.B(n_1096),
.Y(n_1583)
);

AND2x6_ASAP7_75t_L g1584 ( 
.A(n_1486),
.B(n_683),
.Y(n_1584)
);

OAI21x1_ASAP7_75t_L g1585 ( 
.A1(n_1436),
.A2(n_1105),
.B(n_1273),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1437),
.B(n_1441),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1444),
.B(n_1347),
.Y(n_1587)
);

OAI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1450),
.A2(n_1307),
.B(n_1298),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1445),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1563),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1504),
.B(n_1367),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1563),
.Y(n_1592)
);

OA21x2_ASAP7_75t_L g1593 ( 
.A1(n_1505),
.A2(n_1483),
.B(n_1450),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1575),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1575),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1502),
.A2(n_1483),
.B(n_1466),
.Y(n_1596)
);

AOI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1530),
.A2(n_1461),
.B1(n_1424),
.B2(n_1427),
.Y(n_1597)
);

OR2x6_ASAP7_75t_L g1598 ( 
.A(n_1574),
.B(n_1532),
.Y(n_1598)
);

OAI21x1_ASAP7_75t_L g1599 ( 
.A1(n_1583),
.A2(n_1466),
.B(n_1459),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1540),
.A2(n_1453),
.B(n_1389),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1583),
.Y(n_1601)
);

INVxp33_ASAP7_75t_L g1602 ( 
.A(n_1554),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1552),
.A2(n_1369),
.B1(n_1431),
.B2(n_1374),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1575),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1575),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1522),
.B(n_1535),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1503),
.A2(n_1447),
.B1(n_1385),
.B2(n_1364),
.Y(n_1607)
);

NAND2x1p5_ASAP7_75t_L g1608 ( 
.A(n_1521),
.B(n_1389),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1511),
.Y(n_1609)
);

AOI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1539),
.A2(n_1417),
.B(n_1455),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1561),
.A2(n_1105),
.B(n_1456),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1518),
.B(n_1476),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1517),
.A2(n_1453),
.B(n_1389),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1524),
.A2(n_1487),
.B1(n_1471),
.B2(n_1470),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1514),
.B(n_1527),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1507),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1516),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1533),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1527),
.B(n_1476),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1557),
.A2(n_1506),
.B(n_1523),
.Y(n_1620)
);

OR2x6_ASAP7_75t_L g1621 ( 
.A(n_1579),
.B(n_1462),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1561),
.A2(n_1473),
.B(n_1457),
.Y(n_1622)
);

INVxp67_ASAP7_75t_SL g1623 ( 
.A(n_1515),
.Y(n_1623)
);

AOI222xp33_ASAP7_75t_L g1624 ( 
.A1(n_1510),
.A2(n_1362),
.B1(n_574),
.B2(n_555),
.C1(n_595),
.C2(n_562),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_SL g1625 ( 
.A(n_1526),
.B(n_1458),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1537),
.A2(n_1472),
.B(n_1392),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1566),
.A2(n_1496),
.B(n_1479),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1508),
.Y(n_1628)
);

INVx3_ASAP7_75t_L g1629 ( 
.A(n_1521),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1515),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1555),
.B(n_1396),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1527),
.B(n_1366),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1576),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1536),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1589),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1509),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_1507),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1526),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1506),
.A2(n_1307),
.B(n_1298),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1536),
.B(n_1428),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1538),
.A2(n_1453),
.B(n_1389),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1523),
.A2(n_1316),
.B(n_1311),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1597),
.A2(n_1374),
.B1(n_1452),
.B2(n_1446),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1619),
.B(n_1527),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_1616),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1597),
.A2(n_1465),
.B1(n_1379),
.B2(n_1372),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1594),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1615),
.B(n_1553),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_1637),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1640),
.B(n_1573),
.Y(n_1650)
);

A2O1A1Ixp33_ASAP7_75t_L g1651 ( 
.A1(n_1612),
.A2(n_1503),
.B(n_1501),
.C(n_1512),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1624),
.A2(n_1448),
.B1(n_1499),
.B2(n_1495),
.Y(n_1652)
);

OAI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1631),
.A2(n_1513),
.B1(n_1375),
.B2(n_1421),
.Y(n_1653)
);

AOI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1603),
.A2(n_1528),
.B1(n_1499),
.B2(n_1422),
.C(n_1372),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1603),
.A2(n_1421),
.B1(n_1375),
.B2(n_1582),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1624),
.A2(n_1495),
.B1(n_1439),
.B2(n_1460),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1590),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1590),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1600),
.A2(n_1501),
.B(n_1549),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1602),
.B(n_1352),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1594),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1591),
.B(n_1556),
.Y(n_1662)
);

AOI221xp5_ASAP7_75t_L g1663 ( 
.A1(n_1607),
.A2(n_1361),
.B1(n_1416),
.B2(n_515),
.C(n_643),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1614),
.A2(n_1587),
.B1(n_1560),
.B2(n_1361),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1609),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1595),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1600),
.A2(n_1541),
.B(n_1537),
.Y(n_1667)
);

OAI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1631),
.A2(n_1416),
.B1(n_1559),
.B2(n_1491),
.C(n_1464),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1595),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1630),
.Y(n_1670)
);

OAI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1596),
.A2(n_1578),
.B(n_1585),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1590),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1612),
.A2(n_1562),
.B1(n_1586),
.B2(n_1568),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1641),
.A2(n_1542),
.B(n_1572),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1619),
.A2(n_1460),
.B1(n_1572),
.B2(n_1573),
.Y(n_1675)
);

OR2x6_ASAP7_75t_L g1676 ( 
.A(n_1598),
.B(n_1565),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1591),
.B(n_1443),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1640),
.B(n_1581),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1609),
.Y(n_1679)
);

CKINVDCx6p67_ASAP7_75t_R g1680 ( 
.A(n_1616),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1592),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1625),
.A2(n_1404),
.B1(n_1388),
.B2(n_1489),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1640),
.B(n_1581),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1623),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1607),
.A2(n_1562),
.B1(n_1404),
.B2(n_1525),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1632),
.A2(n_1525),
.B1(n_1377),
.B2(n_1378),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1630),
.A2(n_1443),
.B1(n_1468),
.B2(n_1478),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1592),
.Y(n_1688)
);

INVx4_ASAP7_75t_L g1689 ( 
.A(n_1629),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1638),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1604),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1632),
.A2(n_1467),
.B1(n_1464),
.B2(n_1380),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1663),
.A2(n_1606),
.B1(n_1615),
.B2(n_1634),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1652),
.A2(n_1616),
.B1(n_1634),
.B2(n_1360),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1656),
.A2(n_1360),
.B1(n_1606),
.B2(n_1617),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1643),
.A2(n_1360),
.B1(n_1618),
.B2(n_1617),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1662),
.A2(n_1545),
.B1(n_1633),
.B2(n_1618),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1644),
.B(n_1604),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1657),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1644),
.B(n_1605),
.Y(n_1700)
);

NAND3xp33_ASAP7_75t_L g1701 ( 
.A(n_1664),
.B(n_1626),
.C(n_1625),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1648),
.B(n_1605),
.Y(n_1702)
);

BUFx12f_ASAP7_75t_L g1703 ( 
.A(n_1690),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1647),
.Y(n_1704)
);

AOI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1668),
.A2(n_655),
.B1(n_662),
.B2(n_639),
.C(n_629),
.Y(n_1705)
);

AOI222xp33_ASAP7_75t_L g1706 ( 
.A1(n_1654),
.A2(n_597),
.B1(n_582),
.B2(n_598),
.C1(n_589),
.C2(n_571),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1667),
.A2(n_1641),
.B(n_1613),
.Y(n_1707)
);

AOI222xp33_ASAP7_75t_L g1708 ( 
.A1(n_1646),
.A2(n_598),
.B1(n_589),
.B2(n_610),
.C1(n_597),
.C2(n_582),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1673),
.A2(n_1598),
.B1(n_1640),
.B2(n_727),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_1678),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_1649),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1675),
.A2(n_1598),
.B1(n_727),
.B2(n_1428),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1648),
.B(n_1593),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1657),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1653),
.A2(n_1598),
.B1(n_1388),
.B2(n_1485),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1647),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1677),
.B(n_1633),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1685),
.A2(n_1545),
.B1(n_1635),
.B2(n_678),
.Y(n_1718)
);

BUFx3_ASAP7_75t_L g1719 ( 
.A(n_1680),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1661),
.B(n_1593),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1655),
.A2(n_1598),
.B1(n_1482),
.B2(n_1626),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1689),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1658),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1670),
.B(n_1635),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1661),
.B(n_1593),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1658),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1692),
.A2(n_673),
.B1(n_532),
.B2(n_533),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1678),
.A2(n_1478),
.B1(n_1467),
.B2(n_660),
.Y(n_1728)
);

NOR2xp67_ASAP7_75t_L g1729 ( 
.A(n_1674),
.B(n_1613),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1666),
.B(n_1593),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1672),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_SL g1732 ( 
.A1(n_1659),
.A2(n_1370),
.B1(n_1440),
.B2(n_1405),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1666),
.Y(n_1733)
);

OAI21x1_ASAP7_75t_L g1734 ( 
.A1(n_1671),
.A2(n_1620),
.B(n_1596),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1672),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1682),
.A2(n_1370),
.B1(n_1581),
.B2(n_1401),
.Y(n_1736)
);

AOI222xp33_ASAP7_75t_L g1737 ( 
.A1(n_1651),
.A2(n_622),
.B1(n_620),
.B2(n_627),
.C1(n_621),
.C2(n_610),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1684),
.B(n_1592),
.Y(n_1738)
);

AOI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1678),
.A2(n_536),
.B1(n_540),
.B2(n_523),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1684),
.A2(n_1447),
.B1(n_1385),
.B2(n_1453),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1669),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1683),
.A2(n_660),
.B1(n_1438),
.B2(n_1621),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1681),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1683),
.A2(n_660),
.B1(n_1438),
.B2(n_1621),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1683),
.A2(n_660),
.B1(n_1621),
.B2(n_1463),
.Y(n_1745)
);

OAI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1680),
.A2(n_1405),
.B1(n_1381),
.B2(n_1621),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1650),
.A2(n_1621),
.B1(n_1584),
.B2(n_1356),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1689),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1689),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1669),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_SL g1751 ( 
.A1(n_1649),
.A2(n_1584),
.B1(n_1544),
.B2(n_621),
.Y(n_1751)
);

OAI21xp33_ASAP7_75t_L g1752 ( 
.A1(n_1686),
.A2(n_544),
.B(n_541),
.Y(n_1752)
);

AO21x2_ASAP7_75t_L g1753 ( 
.A1(n_1671),
.A2(n_1620),
.B(n_1610),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1691),
.B(n_1577),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1650),
.A2(n_1584),
.B1(n_1356),
.B2(n_622),
.Y(n_1755)
);

OAI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1687),
.A2(n_1403),
.B1(n_1401),
.B2(n_1391),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1660),
.A2(n_1391),
.B1(n_1520),
.B2(n_1629),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1691),
.B(n_1577),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1665),
.B(n_1577),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1679),
.A2(n_1645),
.B1(n_1650),
.B2(n_1681),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1676),
.A2(n_1584),
.B1(n_627),
.B2(n_628),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1676),
.A2(n_1584),
.B1(n_628),
.B2(n_632),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1688),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1676),
.A2(n_632),
.B1(n_649),
.B2(n_620),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1676),
.A2(n_656),
.B1(n_676),
.B2(n_649),
.Y(n_1765)
);

OAI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1690),
.A2(n_676),
.B1(n_680),
.B2(n_656),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1645),
.B(n_1577),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1688),
.A2(n_686),
.B1(n_695),
.B2(n_680),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1652),
.A2(n_695),
.B1(n_699),
.B2(n_686),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1648),
.B(n_1570),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1663),
.A2(n_547),
.B1(n_561),
.B2(n_549),
.C(n_548),
.Y(n_1771)
);

A2O1A1Ixp33_ASAP7_75t_L g1772 ( 
.A1(n_1663),
.A2(n_1544),
.B(n_1548),
.C(n_1627),
.Y(n_1772)
);

OAI211xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1663),
.A2(n_709),
.B(n_699),
.C(n_1571),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1670),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1657),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1684),
.Y(n_1776)
);

AOI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1663),
.A2(n_569),
.B1(n_580),
.B2(n_579),
.C(n_572),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1662),
.B(n_1553),
.Y(n_1778)
);

AOI221xp5_ASAP7_75t_L g1779 ( 
.A1(n_1705),
.A2(n_585),
.B1(n_592),
.B2(n_588),
.C(n_587),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1698),
.B(n_1620),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1704),
.Y(n_1781)
);

BUFx3_ASAP7_75t_L g1782 ( 
.A(n_1719),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1776),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1776),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1698),
.B(n_1610),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1774),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1704),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1716),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1716),
.B(n_1596),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1733),
.B(n_1628),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1702),
.B(n_1570),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1733),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1760),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1741),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1741),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1750),
.Y(n_1796)
);

BUFx2_ASAP7_75t_L g1797 ( 
.A(n_1720),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1750),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1720),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1713),
.B(n_1628),
.Y(n_1800)
);

BUFx2_ASAP7_75t_SL g1801 ( 
.A(n_1719),
.Y(n_1801)
);

OR2x6_ASAP7_75t_L g1802 ( 
.A(n_1707),
.B(n_1628),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1700),
.B(n_717),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1700),
.B(n_1713),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1754),
.B(n_717),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1754),
.B(n_717),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1758),
.Y(n_1807)
);

INVxp67_ASAP7_75t_L g1808 ( 
.A(n_1724),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1758),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1725),
.B(n_717),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1702),
.B(n_1570),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1710),
.B(n_1636),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1725),
.B(n_717),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1730),
.B(n_1770),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1730),
.Y(n_1815)
);

BUFx3_ASAP7_75t_L g1816 ( 
.A(n_1710),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1699),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1711),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1759),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1770),
.B(n_1778),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1759),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1737),
.A2(n_709),
.B1(n_604),
.B2(n_608),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1699),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1714),
.Y(n_1824)
);

INVx4_ASAP7_75t_L g1825 ( 
.A(n_1722),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1760),
.Y(n_1826)
);

INVx3_ASAP7_75t_L g1827 ( 
.A(n_1734),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1710),
.B(n_717),
.Y(n_1828)
);

BUFx3_ASAP7_75t_L g1829 ( 
.A(n_1710),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1714),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1710),
.B(n_1553),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1723),
.B(n_1636),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1738),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1767),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1723),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1726),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1726),
.B(n_1553),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1731),
.B(n_1601),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1731),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1735),
.B(n_1601),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1735),
.Y(n_1841)
);

OAI222xp33_ASAP7_75t_L g1842 ( 
.A1(n_1718),
.A2(n_612),
.B1(n_609),
.B2(n_614),
.C1(n_611),
.C2(n_603),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1743),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1743),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1763),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1763),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1775),
.B(n_1721),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1775),
.Y(n_1848)
);

NOR2x1p5_ASAP7_75t_L g1849 ( 
.A(n_1701),
.B(n_1629),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1734),
.Y(n_1850)
);

OAI221xp5_ASAP7_75t_SL g1851 ( 
.A1(n_1706),
.A2(n_631),
.B1(n_633),
.B2(n_618),
.C(n_616),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1753),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1753),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1753),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1697),
.Y(n_1855)
);

AOI33xp33_ASAP7_75t_L g1856 ( 
.A1(n_1766),
.A2(n_11),
.A3(n_13),
.B1(n_7),
.B2(n_10),
.B3(n_12),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1722),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1722),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1697),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1717),
.B(n_1570),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1701),
.B(n_1601),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1748),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1748),
.B(n_1642),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1748),
.B(n_1642),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1693),
.A2(n_1727),
.B1(n_1732),
.B2(n_1715),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1718),
.B(n_635),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1749),
.B(n_1642),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1729),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1737),
.B(n_636),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1749),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1696),
.B(n_640),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1749),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_1711),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1709),
.B(n_1639),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1772),
.B(n_1639),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1695),
.B(n_1636),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1757),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1729),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1740),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1740),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1694),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1764),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1765),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1739),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1746),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1739),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_1703),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1736),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1751),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1712),
.B(n_1639),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1706),
.B(n_1708),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1769),
.Y(n_1892)
);

BUFx2_ASAP7_75t_L g1893 ( 
.A(n_1756),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1708),
.B(n_1727),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_1703),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1761),
.B(n_1622),
.Y(n_1896)
);

INVx3_ASAP7_75t_L g1897 ( 
.A(n_1747),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1769),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1762),
.A2(n_1542),
.B(n_1534),
.Y(n_1899)
);

BUFx6f_ASAP7_75t_L g1900 ( 
.A(n_1742),
.Y(n_1900)
);

BUFx3_ASAP7_75t_L g1901 ( 
.A(n_1744),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1768),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1773),
.B(n_1571),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1745),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1728),
.B(n_1622),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1752),
.B(n_1519),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1752),
.B(n_1627),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1777),
.B(n_641),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1755),
.B(n_478),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1771),
.Y(n_1910)
);

INVx2_ASAP7_75t_SL g1911 ( 
.A(n_1776),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1774),
.B(n_642),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1704),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1776),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1704),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1704),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_1776),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1704),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1698),
.B(n_478),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1704),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1704),
.Y(n_1921)
);

OAI321xp33_ASAP7_75t_L g1922 ( 
.A1(n_1773),
.A2(n_506),
.A3(n_478),
.B1(n_683),
.B2(n_1520),
.C(n_1588),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1704),
.Y(n_1923)
);

INVx2_ASAP7_75t_SL g1924 ( 
.A(n_1776),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1702),
.B(n_1519),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1698),
.B(n_478),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1698),
.B(n_506),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1704),
.Y(n_1928)
);

OA21x2_ASAP7_75t_L g1929 ( 
.A1(n_1852),
.A2(n_1611),
.B(n_1548),
.Y(n_1929)
);

OAI221xp5_ASAP7_75t_L g1930 ( 
.A1(n_1822),
.A2(n_646),
.B1(n_650),
.B2(n_647),
.C(n_645),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1808),
.B(n_652),
.Y(n_1931)
);

AO21x2_ASAP7_75t_L g1932 ( 
.A1(n_1852),
.A2(n_1611),
.B(n_1550),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1781),
.Y(n_1933)
);

CKINVDCx20_ASAP7_75t_R g1934 ( 
.A(n_1873),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1804),
.B(n_506),
.Y(n_1935)
);

INVx2_ASAP7_75t_SL g1936 ( 
.A(n_1895),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1781),
.Y(n_1937)
);

INVx2_ASAP7_75t_SL g1938 ( 
.A(n_1895),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1782),
.Y(n_1939)
);

BUFx3_ASAP7_75t_L g1940 ( 
.A(n_1782),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1804),
.B(n_506),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1786),
.B(n_506),
.Y(n_1942)
);

INVxp67_ASAP7_75t_SL g1943 ( 
.A(n_1854),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1833),
.B(n_654),
.Y(n_1944)
);

NAND2xp33_ASAP7_75t_R g1945 ( 
.A(n_1893),
.B(n_10),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1792),
.Y(n_1946)
);

AOI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1891),
.A2(n_506),
.B1(n_658),
.B2(n_657),
.Y(n_1947)
);

NAND3xp33_ASAP7_75t_L g1948 ( 
.A(n_1866),
.B(n_683),
.C(n_663),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1792),
.Y(n_1949)
);

NAND3xp33_ASAP7_75t_L g1950 ( 
.A(n_1910),
.B(n_683),
.C(n_665),
.Y(n_1950)
);

AND2x4_ASAP7_75t_L g1951 ( 
.A(n_1911),
.B(n_1629),
.Y(n_1951)
);

AO21x2_ASAP7_75t_L g1952 ( 
.A1(n_1854),
.A2(n_1599),
.B(n_1543),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1796),
.Y(n_1953)
);

NAND4xp25_ASAP7_75t_L g1954 ( 
.A(n_1822),
.B(n_667),
.C(n_669),
.D(n_659),
.Y(n_1954)
);

AOI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1922),
.A2(n_1531),
.B(n_1546),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1784),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1796),
.Y(n_1957)
);

OAI222xp33_ASAP7_75t_L g1958 ( 
.A1(n_1894),
.A2(n_690),
.B1(n_715),
.B2(n_712),
.C1(n_711),
.C2(n_710),
.Y(n_1958)
);

AOI22xp33_ASAP7_75t_L g1959 ( 
.A1(n_1910),
.A2(n_677),
.B1(n_687),
.B2(n_671),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1803),
.B(n_1805),
.Y(n_1960)
);

AOI22xp33_ASAP7_75t_L g1961 ( 
.A1(n_1910),
.A2(n_1901),
.B1(n_1900),
.B2(n_1886),
.Y(n_1961)
);

OAI21xp5_ASAP7_75t_SL g1962 ( 
.A1(n_1842),
.A2(n_683),
.B(n_1608),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1911),
.B(n_1599),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1803),
.B(n_688),
.Y(n_1964)
);

CKINVDCx20_ASAP7_75t_R g1965 ( 
.A(n_1818),
.Y(n_1965)
);

AO21x2_ASAP7_75t_L g1966 ( 
.A1(n_1853),
.A2(n_1543),
.B(n_1551),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_R g1967 ( 
.A(n_1887),
.B(n_1885),
.Y(n_1967)
);

AOI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1865),
.A2(n_694),
.B1(n_700),
.B2(n_693),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1798),
.Y(n_1969)
);

NOR2x1_ASAP7_75t_L g1970 ( 
.A(n_1801),
.B(n_683),
.Y(n_1970)
);

AOI221xp5_ASAP7_75t_L g1971 ( 
.A1(n_1851),
.A2(n_1779),
.B1(n_1886),
.B2(n_1884),
.C(n_1871),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1901),
.A2(n_705),
.B1(n_707),
.B2(n_704),
.Y(n_1972)
);

A2O1A1Ixp33_ASAP7_75t_L g1973 ( 
.A1(n_1856),
.A2(n_661),
.B(n_674),
.C(n_651),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1798),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1913),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1784),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1913),
.Y(n_1977)
);

NOR2xp67_ASAP7_75t_L g1978 ( 
.A(n_1912),
.B(n_12),
.Y(n_1978)
);

OAI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1901),
.A2(n_1608),
.B1(n_1521),
.B2(n_681),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1916),
.Y(n_1980)
);

AOI221xp5_ASAP7_75t_L g1981 ( 
.A1(n_1884),
.A2(n_684),
.B1(n_689),
.B2(n_682),
.C(n_679),
.Y(n_1981)
);

INVxp67_ASAP7_75t_L g1982 ( 
.A(n_1783),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1805),
.B(n_13),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1797),
.B(n_1519),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1916),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1924),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1924),
.Y(n_1987)
);

AOI33xp33_ASAP7_75t_L g1988 ( 
.A1(n_1855),
.A2(n_14),
.A3(n_16),
.B1(n_18),
.B2(n_20),
.B3(n_21),
.Y(n_1988)
);

HB1xp67_ASAP7_75t_L g1989 ( 
.A(n_1914),
.Y(n_1989)
);

AOI22xp33_ASAP7_75t_L g1990 ( 
.A1(n_1900),
.A2(n_1472),
.B1(n_1547),
.B2(n_1551),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1900),
.B(n_1521),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1817),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1917),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1817),
.Y(n_1994)
);

OAI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1869),
.A2(n_706),
.B(n_698),
.Y(n_1995)
);

AOI22xp5_ASAP7_75t_L g1996 ( 
.A1(n_1900),
.A2(n_1472),
.B1(n_716),
.B2(n_1608),
.Y(n_1996)
);

OAI33xp33_ASAP7_75t_L g1997 ( 
.A1(n_1908),
.A2(n_14),
.A3(n_21),
.B1(n_22),
.B2(n_23),
.B3(n_24),
.Y(n_1997)
);

AOI22xp33_ASAP7_75t_SL g1998 ( 
.A1(n_1900),
.A2(n_1472),
.B1(n_26),
.B2(n_22),
.Y(n_1998)
);

AOI22xp33_ASAP7_75t_L g1999 ( 
.A1(n_1900),
.A2(n_1472),
.B1(n_28),
.B2(n_24),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1885),
.B(n_27),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1918),
.Y(n_2001)
);

AOI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1903),
.A2(n_1558),
.B1(n_1475),
.B2(n_1564),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1806),
.B(n_1810),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1814),
.B(n_1519),
.Y(n_2004)
);

NAND3xp33_ASAP7_75t_L g2005 ( 
.A(n_1893),
.B(n_1386),
.C(n_1359),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1823),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1814),
.B(n_28),
.Y(n_2007)
);

AO21x2_ASAP7_75t_L g2008 ( 
.A1(n_1853),
.A2(n_1529),
.B(n_1316),
.Y(n_2008)
);

BUFx8_ASAP7_75t_L g2009 ( 
.A(n_1919),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1918),
.Y(n_2010)
);

AOI22xp33_ASAP7_75t_SL g2011 ( 
.A1(n_1904),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_2011)
);

AOI221xp5_ASAP7_75t_L g2012 ( 
.A1(n_1889),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.C(n_34),
.Y(n_2012)
);

OAI21xp33_ASAP7_75t_L g2013 ( 
.A1(n_1855),
.A2(n_1334),
.B(n_1311),
.Y(n_2013)
);

INVx2_ASAP7_75t_SL g2014 ( 
.A(n_1782),
.Y(n_2014)
);

OAI211xp5_ASAP7_75t_L g2015 ( 
.A1(n_1889),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_2015)
);

BUFx2_ASAP7_75t_L g2016 ( 
.A(n_1816),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1816),
.B(n_35),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1806),
.B(n_36),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1816),
.B(n_37),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1920),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1920),
.Y(n_2021)
);

AOI221xp5_ASAP7_75t_L g2022 ( 
.A1(n_1859),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.C(n_41),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1810),
.B(n_38),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1823),
.Y(n_2024)
);

AOI22xp33_ASAP7_75t_SL g2025 ( 
.A1(n_1897),
.A2(n_42),
.B1(n_39),
.B2(n_40),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1823),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_R g2027 ( 
.A(n_1897),
.B(n_42),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1824),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1888),
.B(n_43),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1928),
.Y(n_2030)
);

NAND3xp33_ASAP7_75t_L g2031 ( 
.A(n_1868),
.B(n_1386),
.C(n_1359),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1824),
.Y(n_2032)
);

AOI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_1882),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_2033)
);

AOI22xp33_ASAP7_75t_L g2034 ( 
.A1(n_1882),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1928),
.Y(n_2035)
);

INVx1_ASAP7_75t_SL g2036 ( 
.A(n_1801),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1787),
.Y(n_2037)
);

OAI221xp5_ASAP7_75t_L g2038 ( 
.A1(n_1883),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.C(n_51),
.Y(n_2038)
);

AOI22xp33_ASAP7_75t_L g2039 ( 
.A1(n_1883),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_2039)
);

NAND4xp25_ASAP7_75t_L g2040 ( 
.A(n_1859),
.B(n_55),
.C(n_53),
.D(n_54),
.Y(n_2040)
);

AOI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_1897),
.A2(n_1475),
.B1(n_1386),
.B2(n_1390),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1787),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1824),
.Y(n_2043)
);

INVxp67_ASAP7_75t_L g2044 ( 
.A(n_1793),
.Y(n_2044)
);

OAI33xp33_ASAP7_75t_L g2045 ( 
.A1(n_1902),
.A2(n_56),
.A3(n_57),
.B1(n_58),
.B2(n_59),
.B3(n_60),
.Y(n_2045)
);

BUFx2_ASAP7_75t_L g2046 ( 
.A(n_1829),
.Y(n_2046)
);

INVx4_ASAP7_75t_L g2047 ( 
.A(n_1828),
.Y(n_2047)
);

NAND4xp25_ASAP7_75t_L g2048 ( 
.A(n_1919),
.B(n_58),
.C(n_56),
.D(n_57),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1787),
.Y(n_2049)
);

AO21x2_ASAP7_75t_L g2050 ( 
.A1(n_1850),
.A2(n_1878),
.B(n_1868),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1794),
.Y(n_2051)
);

AOI22xp33_ASAP7_75t_SL g2052 ( 
.A1(n_1897),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1794),
.Y(n_2053)
);

BUFx3_ASAP7_75t_L g2054 ( 
.A(n_1829),
.Y(n_2054)
);

OAI221xp5_ASAP7_75t_L g2055 ( 
.A1(n_1888),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.C(n_66),
.Y(n_2055)
);

BUFx2_ASAP7_75t_L g2056 ( 
.A(n_1829),
.Y(n_2056)
);

OAI31xp33_ASAP7_75t_L g2057 ( 
.A1(n_1849),
.A2(n_69),
.A3(n_64),
.B(n_67),
.Y(n_2057)
);

INVx5_ASAP7_75t_L g2058 ( 
.A(n_1827),
.Y(n_2058)
);

AOI31xp33_ASAP7_75t_L g2059 ( 
.A1(n_1826),
.A2(n_71),
.A3(n_67),
.B(n_70),
.Y(n_2059)
);

OA21x2_ASAP7_75t_L g2060 ( 
.A1(n_1850),
.A2(n_1567),
.B(n_1344),
.Y(n_2060)
);

AOI221xp5_ASAP7_75t_SL g2061 ( 
.A1(n_1926),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.C(n_78),
.Y(n_2061)
);

INVx1_ASAP7_75t_SL g2062 ( 
.A(n_1820),
.Y(n_2062)
);

AOI221xp5_ASAP7_75t_L g2063 ( 
.A1(n_1902),
.A2(n_72),
.B1(n_74),
.B2(n_79),
.C(n_82),
.Y(n_2063)
);

OAI221xp5_ASAP7_75t_L g2064 ( 
.A1(n_1881),
.A2(n_1878),
.B1(n_1877),
.B2(n_1892),
.C(n_1898),
.Y(n_2064)
);

NAND3xp33_ASAP7_75t_L g2065 ( 
.A(n_1881),
.B(n_1386),
.C(n_1359),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_L g2066 ( 
.A1(n_1892),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_2066)
);

OAI221xp5_ASAP7_75t_SL g2067 ( 
.A1(n_1881),
.A2(n_1906),
.B1(n_1909),
.B2(n_1898),
.C(n_1880),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_1799),
.Y(n_2068)
);

AOI221xp5_ASAP7_75t_L g2069 ( 
.A1(n_1834),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.C(n_87),
.Y(n_2069)
);

OAI31xp33_ASAP7_75t_L g2070 ( 
.A1(n_1849),
.A2(n_88),
.A3(n_86),
.B(n_87),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_2062),
.B(n_1799),
.Y(n_2071)
);

INVxp67_ASAP7_75t_SL g2072 ( 
.A(n_2044),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_1989),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1933),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_2016),
.B(n_1797),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1937),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2046),
.B(n_1799),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1946),
.Y(n_2078)
);

INVx1_ASAP7_75t_SL g2079 ( 
.A(n_1967),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2050),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1949),
.Y(n_2081)
);

AND2x4_ASAP7_75t_L g2082 ( 
.A(n_2058),
.B(n_1815),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1953),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_2050),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1957),
.Y(n_2085)
);

HB1xp67_ASAP7_75t_L g2086 ( 
.A(n_1989),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1969),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2044),
.B(n_1813),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_2056),
.B(n_1815),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_2068),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2068),
.B(n_1780),
.Y(n_2091)
);

OAI31xp33_ASAP7_75t_SL g2092 ( 
.A1(n_2000),
.A2(n_1828),
.A3(n_1813),
.B(n_1875),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1956),
.B(n_1780),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1982),
.B(n_1861),
.Y(n_2094)
);

BUFx3_ASAP7_75t_L g2095 ( 
.A(n_1939),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_2037),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_2058),
.B(n_1807),
.Y(n_2097)
);

INVx1_ASAP7_75t_SL g2098 ( 
.A(n_1965),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_1976),
.B(n_1820),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1974),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1975),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1982),
.B(n_1861),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_1993),
.B(n_1807),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1977),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_2042),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_1993),
.B(n_1809),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2003),
.B(n_1877),
.Y(n_2107)
);

INVx3_ASAP7_75t_L g2108 ( 
.A(n_2058),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_1986),
.B(n_1809),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_1987),
.B(n_1819),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_2049),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_2051),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_1960),
.B(n_1819),
.Y(n_2113)
);

NAND4xp25_ASAP7_75t_L g2114 ( 
.A(n_1968),
.B(n_1926),
.C(n_1927),
.D(n_1877),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1980),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_2058),
.B(n_1821),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2004),
.B(n_1821),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_2053),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1985),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2001),
.Y(n_2120)
);

AND2x2_ASAP7_75t_SL g2121 ( 
.A(n_1988),
.B(n_1875),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2006),
.B(n_1800),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2024),
.B(n_1800),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2026),
.B(n_1800),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1961),
.B(n_1785),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2028),
.B(n_2032),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2043),
.B(n_1800),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2010),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1961),
.B(n_1785),
.Y(n_2129)
);

OR2x2_ASAP7_75t_L g2130 ( 
.A(n_1992),
.B(n_1925),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1935),
.B(n_1847),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2020),
.Y(n_2132)
);

AND2x4_ASAP7_75t_L g2133 ( 
.A(n_2054),
.B(n_1794),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_1994),
.B(n_1831),
.Y(n_2134)
);

NOR2xp33_ASAP7_75t_L g2135 ( 
.A(n_1944),
.B(n_1927),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2021),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1941),
.B(n_1847),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1942),
.B(n_1831),
.Y(n_2138)
);

BUFx2_ASAP7_75t_L g2139 ( 
.A(n_1940),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2014),
.B(n_1863),
.Y(n_2140)
);

INVx2_ASAP7_75t_SL g2141 ( 
.A(n_2036),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2030),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2035),
.B(n_1879),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_1963),
.B(n_1863),
.Y(n_2144)
);

OAI33xp33_ASAP7_75t_L g2145 ( 
.A1(n_2040),
.A2(n_1880),
.A3(n_1879),
.B1(n_1860),
.B2(n_1925),
.B3(n_1839),
.Y(n_2145)
);

AOI22xp33_ASAP7_75t_L g2146 ( 
.A1(n_1947),
.A2(n_1898),
.B1(n_1909),
.B2(n_1906),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1943),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_SL g2148 ( 
.A(n_2027),
.B(n_2047),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1943),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_2029),
.B(n_1905),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1984),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_1963),
.B(n_1864),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1952),
.Y(n_2153)
);

AND2x4_ASAP7_75t_SL g2154 ( 
.A(n_2047),
.B(n_1825),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2007),
.B(n_1907),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2064),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_1936),
.B(n_1864),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1951),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1951),
.Y(n_2159)
);

HB1xp67_ASAP7_75t_L g2160 ( 
.A(n_1938),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2017),
.B(n_1867),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2019),
.B(n_1867),
.Y(n_2162)
);

OR2x2_ASAP7_75t_L g2163 ( 
.A(n_1983),
.B(n_1795),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2067),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2067),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2029),
.B(n_1907),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_1952),
.B(n_1795),
.Y(n_2167)
);

OR2x2_ASAP7_75t_SL g2168 ( 
.A(n_1945),
.B(n_1876),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_1966),
.B(n_1795),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_1966),
.B(n_1915),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2018),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2023),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_1929),
.B(n_1915),
.Y(n_2173)
);

NOR2x1_ASAP7_75t_L g2174 ( 
.A(n_1970),
.B(n_1825),
.Y(n_2174)
);

OR2x2_ASAP7_75t_L g2175 ( 
.A(n_1964),
.B(n_1915),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1929),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2000),
.B(n_1905),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_1932),
.B(n_1921),
.Y(n_2178)
);

AND2x4_ASAP7_75t_L g2179 ( 
.A(n_1991),
.B(n_1921),
.Y(n_2179)
);

NOR2xp67_ASAP7_75t_L g2180 ( 
.A(n_1931),
.B(n_1827),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_2008),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_1932),
.B(n_1921),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2008),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2027),
.B(n_1923),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2005),
.B(n_1923),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2060),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2031),
.Y(n_2187)
);

OR2x2_ASAP7_75t_L g2188 ( 
.A(n_2065),
.B(n_1923),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2009),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2009),
.B(n_1788),
.Y(n_2190)
);

BUFx2_ASAP7_75t_L g2191 ( 
.A(n_1934),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_2060),
.B(n_1791),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2041),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1971),
.B(n_1788),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2013),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_1978),
.B(n_1870),
.Y(n_2196)
);

OR2x2_ASAP7_75t_L g2197 ( 
.A(n_2048),
.B(n_1791),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1950),
.Y(n_2198)
);

AND2x4_ASAP7_75t_L g2199 ( 
.A(n_2002),
.B(n_1870),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2059),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2015),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2038),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2055),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_1990),
.B(n_1870),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1948),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2061),
.B(n_1837),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_1990),
.B(n_1811),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2070),
.B(n_1837),
.Y(n_2208)
);

OR2x2_ASAP7_75t_L g2209 ( 
.A(n_2057),
.B(n_1811),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2069),
.B(n_1830),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2128),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2156),
.B(n_1790),
.Y(n_2212)
);

INVx1_ASAP7_75t_SL g2213 ( 
.A(n_2168),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2128),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2097),
.Y(n_2215)
);

NOR2x1_ASAP7_75t_R g2216 ( 
.A(n_2148),
.B(n_2191),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2072),
.B(n_1790),
.Y(n_2217)
);

HB1xp67_ASAP7_75t_L g2218 ( 
.A(n_2073),
.Y(n_2218)
);

OR2x2_ASAP7_75t_L g2219 ( 
.A(n_2099),
.B(n_2088),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2142),
.Y(n_2220)
);

INVx2_ASAP7_75t_SL g2221 ( 
.A(n_2095),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2080),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2080),
.Y(n_2223)
);

OR2x2_ASAP7_75t_L g2224 ( 
.A(n_2094),
.B(n_1876),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2142),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2144),
.B(n_1872),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2164),
.B(n_1790),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2097),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2074),
.Y(n_2229)
);

INVx1_ASAP7_75t_SL g2230 ( 
.A(n_2079),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2076),
.Y(n_2231)
);

OR2x2_ASAP7_75t_L g2232 ( 
.A(n_2102),
.B(n_1830),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_2125),
.B(n_1839),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2165),
.B(n_2147),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2078),
.Y(n_2235)
);

NAND2x1p5_ASAP7_75t_L g2236 ( 
.A(n_2174),
.B(n_1825),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2081),
.Y(n_2237)
);

HB1xp67_ASAP7_75t_L g2238 ( 
.A(n_2086),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2144),
.B(n_1872),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_2152),
.B(n_1872),
.Y(n_2240)
);

AOI21xp5_ASAP7_75t_SL g2241 ( 
.A1(n_2148),
.A2(n_1979),
.B(n_1973),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2083),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2097),
.Y(n_2243)
);

INVx4_ASAP7_75t_L g2244 ( 
.A(n_2196),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2149),
.B(n_1790),
.Y(n_2245)
);

OR2x2_ASAP7_75t_L g2246 ( 
.A(n_2129),
.B(n_1841),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2151),
.B(n_1841),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2152),
.B(n_1812),
.Y(n_2248)
);

AO21x1_ASAP7_75t_L g2249 ( 
.A1(n_2200),
.A2(n_1945),
.B(n_1962),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2161),
.B(n_1812),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2161),
.B(n_1812),
.Y(n_2251)
);

INVx2_ASAP7_75t_SL g2252 ( 
.A(n_2095),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2085),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2138),
.B(n_1843),
.Y(n_2254)
);

INVx3_ASAP7_75t_L g2255 ( 
.A(n_2082),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2087),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_L g2257 ( 
.A(n_2194),
.B(n_1958),
.Y(n_2257)
);

AOI32xp33_ASAP7_75t_L g2258 ( 
.A1(n_2201),
.A2(n_2011),
.A3(n_2025),
.B1(n_2052),
.B2(n_1947),
.Y(n_2258)
);

OR2x2_ASAP7_75t_L g2259 ( 
.A(n_2155),
.B(n_1843),
.Y(n_2259)
);

NOR2x1_ASAP7_75t_L g2260 ( 
.A(n_2180),
.B(n_1979),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2100),
.Y(n_2261)
);

OR2x2_ASAP7_75t_L g2262 ( 
.A(n_2113),
.B(n_1846),
.Y(n_2262)
);

NAND2x1_ASAP7_75t_L g2263 ( 
.A(n_2108),
.B(n_1825),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2162),
.B(n_1812),
.Y(n_2264)
);

INVxp67_ASAP7_75t_L g2265 ( 
.A(n_2184),
.Y(n_2265)
);

AND2x4_ASAP7_75t_L g2266 ( 
.A(n_2196),
.B(n_1857),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2101),
.Y(n_2267)
);

INVx1_ASAP7_75t_SL g2268 ( 
.A(n_2184),
.Y(n_2268)
);

OR2x2_ASAP7_75t_L g2269 ( 
.A(n_2107),
.B(n_1846),
.Y(n_2269)
);

INVx2_ASAP7_75t_SL g2270 ( 
.A(n_2141),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2104),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2115),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2119),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2162),
.B(n_1874),
.Y(n_2274)
);

HB1xp67_ASAP7_75t_L g2275 ( 
.A(n_2167),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2120),
.B(n_1848),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2132),
.Y(n_2277)
);

A2O1A1Ixp33_ASAP7_75t_L g2278 ( 
.A1(n_2202),
.A2(n_2203),
.B(n_2121),
.C(n_2012),
.Y(n_2278)
);

OR2x2_ASAP7_75t_L g2279 ( 
.A(n_2166),
.B(n_2207),
.Y(n_2279)
);

NAND2x1p5_ASAP7_75t_L g2280 ( 
.A(n_2108),
.B(n_1857),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2136),
.Y(n_2281)
);

INVxp67_ASAP7_75t_SL g2282 ( 
.A(n_2084),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2103),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2116),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2171),
.B(n_2172),
.Y(n_2285)
);

INVx1_ASAP7_75t_SL g2286 ( 
.A(n_2185),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2103),
.Y(n_2287)
);

INVx2_ASAP7_75t_SL g2288 ( 
.A(n_2141),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2075),
.B(n_1874),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2075),
.B(n_1858),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2116),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2093),
.B(n_2139),
.Y(n_2292)
);

INVx2_ASAP7_75t_SL g2293 ( 
.A(n_2189),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2106),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2106),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_2207),
.B(n_1848),
.Y(n_2296)
);

INVx3_ASAP7_75t_L g2297 ( 
.A(n_2082),
.Y(n_2297)
);

HB1xp67_ASAP7_75t_L g2298 ( 
.A(n_2167),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2116),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2096),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2093),
.B(n_1858),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2122),
.B(n_1862),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2096),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2122),
.B(n_1862),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2105),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2105),
.Y(n_2306)
);

OR2x2_ASAP7_75t_L g2307 ( 
.A(n_2163),
.B(n_1835),
.Y(n_2307)
);

OR2x2_ASAP7_75t_L g2308 ( 
.A(n_2131),
.B(n_1835),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_2137),
.B(n_1835),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2111),
.Y(n_2310)
);

INVx3_ASAP7_75t_L g2311 ( 
.A(n_2082),
.Y(n_2311)
);

AND2x4_ASAP7_75t_L g2312 ( 
.A(n_2199),
.B(n_1827),
.Y(n_2312)
);

INVx1_ASAP7_75t_SL g2313 ( 
.A(n_2133),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2090),
.B(n_1836),
.Y(n_2314)
);

AND2x4_ASAP7_75t_L g2315 ( 
.A(n_2199),
.B(n_1827),
.Y(n_2315)
);

INVxp67_ASAP7_75t_L g2316 ( 
.A(n_2187),
.Y(n_2316)
);

OR2x2_ASAP7_75t_L g2317 ( 
.A(n_2071),
.B(n_1836),
.Y(n_2317)
);

OR2x2_ASAP7_75t_L g2318 ( 
.A(n_2071),
.B(n_1836),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2111),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2112),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_2084),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2112),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2090),
.B(n_1844),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2118),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2143),
.B(n_1844),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2118),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2123),
.B(n_1890),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2130),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2123),
.B(n_1890),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2130),
.Y(n_2330)
);

OR2x2_ASAP7_75t_L g2331 ( 
.A(n_2213),
.B(n_2177),
.Y(n_2331)
);

OR2x2_ASAP7_75t_L g2332 ( 
.A(n_2213),
.B(n_2175),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2280),
.Y(n_2333)
);

OAI221xp5_ASAP7_75t_L g2334 ( 
.A1(n_2278),
.A2(n_1972),
.B1(n_1959),
.B2(n_1930),
.C(n_2011),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2292),
.B(n_2157),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2229),
.Y(n_2336)
);

AND2x4_ASAP7_75t_L g2337 ( 
.A(n_2244),
.B(n_2108),
.Y(n_2337)
);

INVx1_ASAP7_75t_SL g2338 ( 
.A(n_2230),
.Y(n_2338)
);

OAI211xp5_ASAP7_75t_SL g2339 ( 
.A1(n_2257),
.A2(n_2278),
.B(n_2258),
.C(n_1972),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2280),
.Y(n_2340)
);

NAND2xp33_ASAP7_75t_L g2341 ( 
.A(n_2260),
.B(n_2230),
.Y(n_2341)
);

NAND3xp33_ASAP7_75t_SL g2342 ( 
.A(n_2249),
.B(n_2198),
.C(n_2205),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2268),
.B(n_2157),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2231),
.Y(n_2344)
);

OAI221xp5_ASAP7_75t_L g2345 ( 
.A1(n_2257),
.A2(n_1959),
.B1(n_2146),
.B2(n_2025),
.C(n_2052),
.Y(n_2345)
);

NAND2x1_ASAP7_75t_SL g2346 ( 
.A(n_2244),
.B(n_2160),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2235),
.Y(n_2347)
);

AOI22xp33_ASAP7_75t_L g2348 ( 
.A1(n_2279),
.A2(n_2121),
.B1(n_2150),
.B2(n_2146),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2266),
.Y(n_2349)
);

INVx1_ASAP7_75t_SL g2350 ( 
.A(n_2270),
.Y(n_2350)
);

NAND2xp33_ASAP7_75t_SL g2351 ( 
.A(n_2293),
.B(n_2197),
.Y(n_2351)
);

NAND3xp33_ASAP7_75t_SL g2352 ( 
.A(n_2316),
.B(n_2063),
.C(n_2022),
.Y(n_2352)
);

NOR2x1_ASAP7_75t_SL g2353 ( 
.A(n_2288),
.B(n_2188),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2268),
.B(n_2215),
.Y(n_2354)
);

NOR2xp33_ASAP7_75t_L g2355 ( 
.A(n_2285),
.B(n_2098),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2237),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2316),
.B(n_2150),
.Y(n_2357)
);

AND2x4_ASAP7_75t_L g2358 ( 
.A(n_2265),
.B(n_2199),
.Y(n_2358)
);

NOR2x1_ASAP7_75t_L g2359 ( 
.A(n_2234),
.B(n_2190),
.Y(n_2359)
);

INVx1_ASAP7_75t_SL g2360 ( 
.A(n_2221),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2228),
.B(n_2124),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2286),
.B(n_2195),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2242),
.Y(n_2363)
);

INVxp67_ASAP7_75t_SL g2364 ( 
.A(n_2216),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2243),
.B(n_2124),
.Y(n_2365)
);

HB1xp67_ASAP7_75t_L g2366 ( 
.A(n_2218),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2284),
.B(n_2127),
.Y(n_2367)
);

NOR2xp33_ASAP7_75t_L g2368 ( 
.A(n_2285),
.B(n_2135),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2291),
.B(n_2127),
.Y(n_2369)
);

INVxp67_ASAP7_75t_L g2370 ( 
.A(n_2234),
.Y(n_2370)
);

AOI22xp33_ASAP7_75t_L g2371 ( 
.A1(n_2212),
.A2(n_2145),
.B1(n_1997),
.B2(n_2045),
.Y(n_2371)
);

NAND2xp33_ASAP7_75t_R g2372 ( 
.A(n_2255),
.B(n_2197),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2253),
.Y(n_2373)
);

NAND4xp25_ASAP7_75t_L g2374 ( 
.A(n_2241),
.B(n_2135),
.C(n_2034),
.D(n_2039),
.Y(n_2374)
);

INVx2_ASAP7_75t_SL g2375 ( 
.A(n_2252),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2256),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2299),
.B(n_2140),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2261),
.Y(n_2378)
);

BUFx3_ASAP7_75t_L g2379 ( 
.A(n_2227),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2267),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2271),
.Y(n_2381)
);

NAND2xp33_ASAP7_75t_SL g2382 ( 
.A(n_2263),
.B(n_2206),
.Y(n_2382)
);

NOR4xp25_ASAP7_75t_SL g2383 ( 
.A(n_2282),
.B(n_2193),
.C(n_2092),
.D(n_2159),
.Y(n_2383)
);

NAND2xp33_ASAP7_75t_SL g2384 ( 
.A(n_2218),
.B(n_2209),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2286),
.B(n_2173),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_2265),
.B(n_2140),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_2274),
.B(n_2117),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2272),
.B(n_2173),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2248),
.B(n_2117),
.Y(n_2389)
);

NOR2xp33_ASAP7_75t_L g2390 ( 
.A(n_2227),
.B(n_1958),
.Y(n_2390)
);

OR2x2_ASAP7_75t_L g2391 ( 
.A(n_2212),
.B(n_2209),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2273),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2277),
.Y(n_2393)
);

BUFx2_ASAP7_75t_L g2394 ( 
.A(n_2238),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2266),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2281),
.B(n_2091),
.Y(n_2396)
);

NAND2xp33_ASAP7_75t_R g2397 ( 
.A(n_2255),
.B(n_2210),
.Y(n_2397)
);

NAND3xp33_ASAP7_75t_L g2398 ( 
.A(n_2238),
.B(n_1998),
.C(n_2033),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2328),
.B(n_2091),
.Y(n_2399)
);

OR2x2_ASAP7_75t_L g2400 ( 
.A(n_2219),
.B(n_2208),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2289),
.B(n_2134),
.Y(n_2401)
);

INVx2_ASAP7_75t_SL g2402 ( 
.A(n_2297),
.Y(n_2402)
);

AOI31xp33_ASAP7_75t_L g2403 ( 
.A1(n_2236),
.A2(n_2045),
.A3(n_1997),
.B(n_1998),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2276),
.Y(n_2404)
);

OAI221xp5_ASAP7_75t_L g2405 ( 
.A1(n_2236),
.A2(n_1954),
.B1(n_1995),
.B2(n_2034),
.C(n_2033),
.Y(n_2405)
);

OAI31xp33_ASAP7_75t_SL g2406 ( 
.A1(n_2313),
.A2(n_2114),
.A3(n_2204),
.B(n_2089),
.Y(n_2406)
);

INVxp67_ASAP7_75t_L g2407 ( 
.A(n_2276),
.Y(n_2407)
);

OAI211xp5_ASAP7_75t_L g2408 ( 
.A1(n_2275),
.A2(n_2039),
.B(n_2066),
.C(n_1999),
.Y(n_2408)
);

OR2x2_ASAP7_75t_L g2409 ( 
.A(n_2224),
.B(n_2192),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_2233),
.B(n_2158),
.Y(n_2410)
);

INVx3_ASAP7_75t_L g2411 ( 
.A(n_2297),
.Y(n_2411)
);

OR2x2_ASAP7_75t_L g2412 ( 
.A(n_2246),
.B(n_2134),
.Y(n_2412)
);

AND2x4_ASAP7_75t_SL g2413 ( 
.A(n_2290),
.B(n_2179),
.Y(n_2413)
);

OR2x2_ASAP7_75t_L g2414 ( 
.A(n_2217),
.B(n_2089),
.Y(n_2414)
);

NAND4xp25_ASAP7_75t_L g2415 ( 
.A(n_2217),
.B(n_2066),
.C(n_1999),
.D(n_1981),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2211),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2330),
.B(n_2283),
.Y(n_2417)
);

INVx1_ASAP7_75t_SL g2418 ( 
.A(n_2313),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2250),
.B(n_2154),
.Y(n_2419)
);

INVx2_ASAP7_75t_SL g2420 ( 
.A(n_2311),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2251),
.B(n_2154),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2287),
.B(n_2109),
.Y(n_2422)
);

OR2x2_ASAP7_75t_L g2423 ( 
.A(n_2296),
.B(n_2077),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2311),
.Y(n_2424)
);

NOR2xp33_ASAP7_75t_L g2425 ( 
.A(n_2254),
.B(n_2308),
.Y(n_2425)
);

NAND3xp33_ASAP7_75t_SL g2426 ( 
.A(n_2275),
.B(n_1996),
.C(n_1955),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2294),
.B(n_2109),
.Y(n_2427)
);

HB1xp67_ASAP7_75t_L g2428 ( 
.A(n_2295),
.Y(n_2428)
);

OR2x2_ASAP7_75t_L g2429 ( 
.A(n_2309),
.B(n_2077),
.Y(n_2429)
);

NOR3xp33_ASAP7_75t_L g2430 ( 
.A(n_2282),
.B(n_2153),
.C(n_2204),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2214),
.Y(n_2431)
);

HB1xp67_ASAP7_75t_L g2432 ( 
.A(n_2245),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2264),
.B(n_2110),
.Y(n_2433)
);

NOR2xp33_ASAP7_75t_L g2434 ( 
.A(n_2259),
.B(n_2133),
.Y(n_2434)
);

INVx1_ASAP7_75t_SL g2435 ( 
.A(n_2245),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2226),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2239),
.Y(n_2437)
);

AOI221xp5_ASAP7_75t_L g2438 ( 
.A1(n_2298),
.A2(n_2182),
.B1(n_2178),
.B2(n_2153),
.C(n_2176),
.Y(n_2438)
);

OR2x2_ASAP7_75t_L g2439 ( 
.A(n_2232),
.B(n_2179),
.Y(n_2439)
);

OR2x2_ASAP7_75t_L g2440 ( 
.A(n_2269),
.B(n_2179),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2220),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2225),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2240),
.Y(n_2443)
);

OAI22xp5_ASAP7_75t_L g2444 ( 
.A1(n_2364),
.A2(n_2315),
.B1(n_2312),
.B2(n_2247),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2366),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2366),
.Y(n_2446)
);

A2O1A1Ixp33_ASAP7_75t_L g2447 ( 
.A1(n_2339),
.A2(n_2298),
.B(n_2315),
.C(n_2312),
.Y(n_2447)
);

AOI22xp5_ASAP7_75t_L g2448 ( 
.A1(n_2339),
.A2(n_2178),
.B1(n_2182),
.B2(n_2300),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2336),
.Y(n_2449)
);

AOI32xp33_ASAP7_75t_L g2450 ( 
.A1(n_2341),
.A2(n_2329),
.A3(n_2327),
.B1(n_2326),
.B2(n_2305),
.Y(n_2450)
);

OAI221xp5_ASAP7_75t_SL g2451 ( 
.A1(n_2348),
.A2(n_1802),
.B1(n_2262),
.B2(n_2247),
.C(n_2176),
.Y(n_2451)
);

AND2x4_ASAP7_75t_L g2452 ( 
.A(n_2338),
.B(n_2319),
.Y(n_2452)
);

OAI21xp5_ASAP7_75t_SL g2453 ( 
.A1(n_2342),
.A2(n_2334),
.B(n_2374),
.Y(n_2453)
);

OAI22xp5_ASAP7_75t_L g2454 ( 
.A1(n_2364),
.A2(n_2345),
.B1(n_2398),
.B2(n_2383),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2411),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2390),
.B(n_2302),
.Y(n_2456)
);

AOI221xp5_ASAP7_75t_L g2457 ( 
.A1(n_2342),
.A2(n_2324),
.B1(n_2303),
.B2(n_2322),
.C(n_2306),
.Y(n_2457)
);

OR2x2_ASAP7_75t_L g2458 ( 
.A(n_2331),
.B(n_2307),
.Y(n_2458)
);

OAI322xp33_ASAP7_75t_L g2459 ( 
.A1(n_2370),
.A2(n_2310),
.A3(n_2320),
.B1(n_2325),
.B2(n_2323),
.C1(n_2314),
.C2(n_2222),
.Y(n_2459)
);

AOI21xp33_ASAP7_75t_L g2460 ( 
.A1(n_2397),
.A2(n_2223),
.B(n_2222),
.Y(n_2460)
);

AND2x4_ASAP7_75t_L g2461 ( 
.A(n_2375),
.B(n_2304),
.Y(n_2461)
);

AOI22xp5_ASAP7_75t_L g2462 ( 
.A1(n_2372),
.A2(n_2325),
.B1(n_2133),
.B2(n_2170),
.Y(n_2462)
);

XNOR2xp5_ASAP7_75t_L g2463 ( 
.A(n_2334),
.B(n_88),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2368),
.B(n_2370),
.Y(n_2464)
);

OAI21xp33_ASAP7_75t_SL g2465 ( 
.A1(n_2346),
.A2(n_2314),
.B(n_2323),
.Y(n_2465)
);

AOI22xp5_ASAP7_75t_L g2466 ( 
.A1(n_2352),
.A2(n_1802),
.B1(n_1896),
.B2(n_2169),
.Y(n_2466)
);

INVx1_ASAP7_75t_SL g2467 ( 
.A(n_2351),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2344),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2347),
.Y(n_2469)
);

NAND3x2_ASAP7_75t_L g2470 ( 
.A(n_2394),
.B(n_2332),
.C(n_2391),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2356),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2359),
.B(n_2301),
.Y(n_2472)
);

INVxp67_ASAP7_75t_L g2473 ( 
.A(n_2384),
.Y(n_2473)
);

AOI211xp5_ASAP7_75t_L g2474 ( 
.A1(n_2345),
.A2(n_2223),
.B(n_2321),
.C(n_2186),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2363),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2373),
.Y(n_2476)
);

OAI221xp5_ASAP7_75t_L g2477 ( 
.A1(n_2406),
.A2(n_2321),
.B1(n_2318),
.B2(n_2317),
.C(n_2186),
.Y(n_2477)
);

INVx2_ASAP7_75t_SL g2478 ( 
.A(n_2337),
.Y(n_2478)
);

OAI21xp5_ASAP7_75t_L g2479 ( 
.A1(n_2426),
.A2(n_2352),
.B(n_2382),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_SL g2480 ( 
.A(n_2362),
.B(n_2357),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2376),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2335),
.B(n_2110),
.Y(n_2482)
);

NAND3xp33_ASAP7_75t_SL g2483 ( 
.A(n_2408),
.B(n_2183),
.C(n_2181),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_L g2484 ( 
.A(n_2360),
.B(n_2126),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2378),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2380),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2381),
.Y(n_2487)
);

NAND3xp33_ASAP7_75t_SL g2488 ( 
.A(n_2408),
.B(n_2183),
.C(n_2181),
.Y(n_2488)
);

AOI221xp5_ASAP7_75t_L g2489 ( 
.A1(n_2426),
.A2(n_2170),
.B1(n_2169),
.B2(n_2126),
.C(n_1896),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2357),
.B(n_1844),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2392),
.Y(n_2491)
);

AOI32xp33_ASAP7_75t_L g2492 ( 
.A1(n_2430),
.A2(n_1789),
.A3(n_1845),
.B1(n_1838),
.B2(n_1840),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2379),
.B(n_1845),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2411),
.Y(n_2494)
);

OR2x2_ASAP7_75t_L g2495 ( 
.A(n_2400),
.B(n_1802),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2371),
.B(n_1845),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2393),
.Y(n_2497)
);

OAI21xp33_ASAP7_75t_L g2498 ( 
.A1(n_2403),
.A2(n_1802),
.B(n_1789),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2416),
.Y(n_2499)
);

AOI21xp33_ASAP7_75t_L g2500 ( 
.A1(n_2405),
.A2(n_1802),
.B(n_89),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2362),
.B(n_1789),
.Y(n_2501)
);

NAND2x1p5_ASAP7_75t_L g2502 ( 
.A(n_2337),
.B(n_1789),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2431),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2441),
.Y(n_2504)
);

OAI21xp33_ASAP7_75t_L g2505 ( 
.A1(n_2415),
.A2(n_1840),
.B(n_1838),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2442),
.Y(n_2506)
);

INVx2_ASAP7_75t_SL g2507 ( 
.A(n_2402),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2428),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2417),
.Y(n_2509)
);

OAI22xp33_ASAP7_75t_L g2510 ( 
.A1(n_2405),
.A2(n_1899),
.B1(n_1832),
.B2(n_92),
.Y(n_2510)
);

OA22x2_ASAP7_75t_L g2511 ( 
.A1(n_2350),
.A2(n_1832),
.B1(n_93),
.B2(n_90),
.Y(n_2511)
);

AND2x4_ASAP7_75t_L g2512 ( 
.A(n_2353),
.B(n_1832),
.Y(n_2512)
);

AOI31xp33_ASAP7_75t_L g2513 ( 
.A1(n_2418),
.A2(n_1832),
.A3(n_94),
.B(n_91),
.Y(n_2513)
);

NAND4xp75_ASAP7_75t_SL g2514 ( 
.A(n_2354),
.B(n_1580),
.C(n_1312),
.D(n_94),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_2355),
.B(n_2386),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2417),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2396),
.Y(n_2517)
);

AOI22xp5_ASAP7_75t_L g2518 ( 
.A1(n_2358),
.A2(n_2410),
.B1(n_2435),
.B2(n_2434),
.Y(n_2518)
);

NOR2x1_ASAP7_75t_L g2519 ( 
.A(n_2424),
.B(n_91),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2420),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2396),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2389),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2404),
.Y(n_2523)
);

OAI221xp5_ASAP7_75t_SL g2524 ( 
.A1(n_2438),
.A2(n_2430),
.B1(n_2385),
.B2(n_2407),
.C(n_2409),
.Y(n_2524)
);

AOI22xp5_ASAP7_75t_L g2525 ( 
.A1(n_2358),
.A2(n_1414),
.B1(n_1474),
.B2(n_1390),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2432),
.B(n_93),
.Y(n_2526)
);

AND2x4_ASAP7_75t_L g2527 ( 
.A(n_2349),
.B(n_99),
.Y(n_2527)
);

OAI21xp5_ASAP7_75t_SL g2528 ( 
.A1(n_2438),
.A2(n_100),
.B(n_101),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2361),
.B(n_100),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2399),
.Y(n_2530)
);

INVxp67_ASAP7_75t_L g2531 ( 
.A(n_2385),
.Y(n_2531)
);

OAI22xp5_ASAP7_75t_SL g2532 ( 
.A1(n_2463),
.A2(n_2340),
.B1(n_2333),
.B2(n_2395),
.Y(n_2532)
);

INVx2_ASAP7_75t_SL g2533 ( 
.A(n_2527),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2445),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2446),
.Y(n_2535)
);

INVx2_ASAP7_75t_SL g2536 ( 
.A(n_2527),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2478),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2502),
.Y(n_2538)
);

NOR2xp33_ASAP7_75t_L g2539 ( 
.A(n_2453),
.B(n_2425),
.Y(n_2539)
);

A2O1A1Ixp33_ASAP7_75t_L g2540 ( 
.A1(n_2528),
.A2(n_2407),
.B(n_2343),
.C(n_2388),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2467),
.B(n_2507),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2499),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2503),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2504),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2506),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2454),
.B(n_2365),
.Y(n_2546)
);

OAI22xp5_ASAP7_75t_L g2547 ( 
.A1(n_2470),
.A2(n_2414),
.B1(n_2399),
.B2(n_2413),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2519),
.B(n_2515),
.Y(n_2548)
);

INVx1_ASAP7_75t_SL g2549 ( 
.A(n_2519),
.Y(n_2549)
);

AOI222xp33_ASAP7_75t_L g2550 ( 
.A1(n_2479),
.A2(n_2388),
.B1(n_2427),
.B2(n_2422),
.C1(n_2377),
.C2(n_2436),
.Y(n_2550)
);

O2A1O1Ixp33_ASAP7_75t_SL g2551 ( 
.A1(n_2500),
.A2(n_2422),
.B(n_2427),
.C(n_2439),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2508),
.B(n_2367),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2449),
.Y(n_2553)
);

OAI21xp5_ASAP7_75t_L g2554 ( 
.A1(n_2513),
.A2(n_2440),
.B(n_2369),
.Y(n_2554)
);

INVx1_ASAP7_75t_SL g2555 ( 
.A(n_2511),
.Y(n_2555)
);

OAI221xp5_ASAP7_75t_L g2556 ( 
.A1(n_2474),
.A2(n_2412),
.B1(n_2423),
.B2(n_2429),
.C(n_2443),
.Y(n_2556)
);

HB1xp67_ASAP7_75t_L g2557 ( 
.A(n_2452),
.Y(n_2557)
);

AOI21xp33_ASAP7_75t_SL g2558 ( 
.A1(n_2510),
.A2(n_102),
.B(n_103),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2526),
.B(n_2401),
.Y(n_2559)
);

OR2x2_ASAP7_75t_L g2560 ( 
.A(n_2480),
.B(n_2496),
.Y(n_2560)
);

OAI22xp5_ASAP7_75t_L g2561 ( 
.A1(n_2473),
.A2(n_2437),
.B1(n_2419),
.B2(n_2421),
.Y(n_2561)
);

HB1xp67_ASAP7_75t_L g2562 ( 
.A(n_2452),
.Y(n_2562)
);

INVxp67_ASAP7_75t_L g2563 ( 
.A(n_2520),
.Y(n_2563)
);

INVx1_ASAP7_75t_SL g2564 ( 
.A(n_2529),
.Y(n_2564)
);

NAND3x1_ASAP7_75t_L g2565 ( 
.A(n_2457),
.B(n_2387),
.C(n_2433),
.Y(n_2565)
);

HB1xp67_ASAP7_75t_L g2566 ( 
.A(n_2484),
.Y(n_2566)
);

OAI33xp33_ASAP7_75t_L g2567 ( 
.A1(n_2464),
.A2(n_102),
.A3(n_103),
.B1(n_104),
.B2(n_105),
.B3(n_106),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2468),
.Y(n_2568)
);

HB1xp67_ASAP7_75t_L g2569 ( 
.A(n_2531),
.Y(n_2569)
);

AOI221x1_ASAP7_75t_L g2570 ( 
.A1(n_2483),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.C(n_107),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2469),
.Y(n_2571)
);

NOR2xp67_ASAP7_75t_L g2572 ( 
.A(n_2465),
.B(n_108),
.Y(n_2572)
);

INVx1_ASAP7_75t_SL g2573 ( 
.A(n_2455),
.Y(n_2573)
);

NAND3xp33_ASAP7_75t_L g2574 ( 
.A(n_2524),
.B(n_108),
.C(n_109),
.Y(n_2574)
);

NAND2x1p5_ASAP7_75t_L g2575 ( 
.A(n_2512),
.B(n_110),
.Y(n_2575)
);

OAI22xp5_ASAP7_75t_L g2576 ( 
.A1(n_2447),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2456),
.B(n_2509),
.Y(n_2577)
);

AND2x2_ASAP7_75t_L g2578 ( 
.A(n_2461),
.B(n_114),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2461),
.B(n_114),
.Y(n_2579)
);

AOI22xp5_ASAP7_75t_L g2580 ( 
.A1(n_2488),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2494),
.Y(n_2581)
);

OR2x2_ASAP7_75t_L g2582 ( 
.A(n_2530),
.B(n_2522),
.Y(n_2582)
);

AOI22xp5_ASAP7_75t_L g2583 ( 
.A1(n_2498),
.A2(n_115),
.B1(n_117),
.B2(n_118),
.Y(n_2583)
);

INVx1_ASAP7_75t_SL g2584 ( 
.A(n_2471),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2475),
.Y(n_2585)
);

NAND2x1_ASAP7_75t_L g2586 ( 
.A(n_2512),
.B(n_119),
.Y(n_2586)
);

OAI22xp5_ASAP7_75t_L g2587 ( 
.A1(n_2451),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2476),
.Y(n_2588)
);

AOI31xp33_ASAP7_75t_L g2589 ( 
.A1(n_2460),
.A2(n_120),
.A3(n_121),
.B(n_122),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2481),
.Y(n_2590)
);

AOI221xp5_ASAP7_75t_L g2591 ( 
.A1(n_2489),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.C(n_126),
.Y(n_2591)
);

NOR2xp33_ASAP7_75t_L g2592 ( 
.A(n_2518),
.B(n_124),
.Y(n_2592)
);

AOI221xp5_ASAP7_75t_L g2593 ( 
.A1(n_2465),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.C(n_130),
.Y(n_2593)
);

OAI22xp5_ASAP7_75t_L g2594 ( 
.A1(n_2466),
.A2(n_129),
.B1(n_131),
.B2(n_134),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2516),
.B(n_134),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2485),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2486),
.Y(n_2597)
);

AOI21xp33_ASAP7_75t_L g2598 ( 
.A1(n_2444),
.A2(n_136),
.B(n_137),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2487),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2517),
.B(n_2521),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2482),
.B(n_136),
.Y(n_2601)
);

AND2x4_ASAP7_75t_L g2602 ( 
.A(n_2491),
.B(n_137),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2458),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2497),
.Y(n_2604)
);

INVxp67_ASAP7_75t_SL g2605 ( 
.A(n_2472),
.Y(n_2605)
);

AOI21xp33_ASAP7_75t_L g2606 ( 
.A1(n_2523),
.A2(n_139),
.B(n_140),
.Y(n_2606)
);

INVxp67_ASAP7_75t_SL g2607 ( 
.A(n_2462),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2495),
.Y(n_2608)
);

NAND3xp33_ASAP7_75t_L g2609 ( 
.A(n_2574),
.B(n_2466),
.C(n_2450),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2541),
.B(n_2505),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2555),
.B(n_2448),
.Y(n_2611)
);

AOI21xp33_ASAP7_75t_L g2612 ( 
.A1(n_2539),
.A2(n_2477),
.B(n_2525),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2557),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2533),
.B(n_2501),
.Y(n_2614)
);

AOI32xp33_ASAP7_75t_L g2615 ( 
.A1(n_2549),
.A2(n_2490),
.A3(n_2459),
.B1(n_2493),
.B2(n_2492),
.Y(n_2615)
);

NOR4xp25_ASAP7_75t_SL g2616 ( 
.A(n_2593),
.B(n_2514),
.C(n_141),
.D(n_142),
.Y(n_2616)
);

INVx1_ASAP7_75t_SL g2617 ( 
.A(n_2549),
.Y(n_2617)
);

NOR2xp33_ASAP7_75t_L g2618 ( 
.A(n_2536),
.B(n_140),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2537),
.B(n_143),
.Y(n_2619)
);

NOR2x1_ASAP7_75t_L g2620 ( 
.A(n_2589),
.B(n_2572),
.Y(n_2620)
);

INVx1_ASAP7_75t_SL g2621 ( 
.A(n_2562),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2564),
.B(n_143),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2569),
.Y(n_2623)
);

AOI21xp33_ASAP7_75t_L g2624 ( 
.A1(n_2576),
.A2(n_145),
.B(n_146),
.Y(n_2624)
);

NOR2xp33_ASAP7_75t_R g2625 ( 
.A(n_2592),
.B(n_146),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_SL g2626 ( 
.A(n_2576),
.B(n_147),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2534),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2535),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2575),
.Y(n_2629)
);

AND2x4_ASAP7_75t_L g2630 ( 
.A(n_2573),
.B(n_147),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2603),
.Y(n_2631)
);

NOR2x1_ASAP7_75t_L g2632 ( 
.A(n_2589),
.B(n_148),
.Y(n_2632)
);

OAI21xp33_ASAP7_75t_SL g2633 ( 
.A1(n_2607),
.A2(n_148),
.B(n_149),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2575),
.Y(n_2634)
);

XOR2x2_ASAP7_75t_L g2635 ( 
.A(n_2532),
.B(n_150),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2604),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_SL g2637 ( 
.A(n_2580),
.B(n_150),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2564),
.B(n_151),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2542),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2555),
.B(n_151),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_L g2641 ( 
.A(n_2548),
.B(n_152),
.Y(n_2641)
);

NOR2xp33_ASAP7_75t_R g2642 ( 
.A(n_2595),
.B(n_153),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2543),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2566),
.B(n_154),
.Y(n_2644)
);

INVx2_ASAP7_75t_SL g2645 ( 
.A(n_2586),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2544),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2545),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_L g2648 ( 
.A(n_2573),
.B(n_2563),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2554),
.B(n_154),
.Y(n_2649)
);

NOR2xp33_ASAP7_75t_L g2650 ( 
.A(n_2546),
.B(n_155),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2554),
.B(n_156),
.Y(n_2651)
);

HB1xp67_ASAP7_75t_L g2652 ( 
.A(n_2584),
.Y(n_2652)
);

XNOR2xp5_ASAP7_75t_L g2653 ( 
.A(n_2565),
.B(n_156),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2553),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2568),
.Y(n_2655)
);

O2A1O1Ixp33_ASAP7_75t_L g2656 ( 
.A1(n_2594),
.A2(n_157),
.B(n_158),
.C(n_159),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2605),
.B(n_158),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2571),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2585),
.Y(n_2659)
);

NAND2xp33_ASAP7_75t_SL g2660 ( 
.A(n_2560),
.B(n_159),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2588),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2538),
.Y(n_2662)
);

NOR2xp33_ASAP7_75t_R g2663 ( 
.A(n_2602),
.B(n_160),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2601),
.B(n_162),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2578),
.B(n_163),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2645),
.B(n_2581),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2620),
.B(n_2579),
.Y(n_2667)
);

NOR3xp33_ASAP7_75t_L g2668 ( 
.A(n_2650),
.B(n_2598),
.C(n_2577),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2652),
.Y(n_2669)
);

AOI21xp5_ASAP7_75t_L g2670 ( 
.A1(n_2626),
.A2(n_2551),
.B(n_2587),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2652),
.Y(n_2671)
);

AOI211x1_ASAP7_75t_L g2672 ( 
.A1(n_2626),
.A2(n_2587),
.B(n_2547),
.C(n_2561),
.Y(n_2672)
);

INVx1_ASAP7_75t_SL g2673 ( 
.A(n_2617),
.Y(n_2673)
);

XNOR2x2_ASAP7_75t_L g2674 ( 
.A(n_2635),
.B(n_2591),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2613),
.Y(n_2675)
);

NAND4xp25_ASAP7_75t_L g2676 ( 
.A(n_2650),
.B(n_2570),
.C(n_2550),
.D(n_2583),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2610),
.B(n_2629),
.Y(n_2677)
);

AOI211xp5_ASAP7_75t_L g2678 ( 
.A1(n_2653),
.A2(n_2558),
.B(n_2606),
.C(n_2540),
.Y(n_2678)
);

NOR2xp67_ASAP7_75t_L g2679 ( 
.A(n_2629),
.B(n_2582),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2632),
.B(n_2584),
.Y(n_2680)
);

NOR4xp25_ASAP7_75t_L g2681 ( 
.A(n_2640),
.B(n_2590),
.C(n_2596),
.D(n_2597),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2630),
.Y(n_2682)
);

OR2x2_ASAP7_75t_L g2683 ( 
.A(n_2621),
.B(n_2559),
.Y(n_2683)
);

INVxp67_ASAP7_75t_L g2684 ( 
.A(n_2660),
.Y(n_2684)
);

NOR3xp33_ASAP7_75t_L g2685 ( 
.A(n_2623),
.B(n_2648),
.C(n_2611),
.Y(n_2685)
);

NOR2xp33_ASAP7_75t_L g2686 ( 
.A(n_2634),
.B(n_2644),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2634),
.Y(n_2687)
);

AOI211xp5_ASAP7_75t_L g2688 ( 
.A1(n_2609),
.A2(n_2567),
.B(n_2600),
.C(n_2599),
.Y(n_2688)
);

INVx2_ASAP7_75t_SL g2689 ( 
.A(n_2663),
.Y(n_2689)
);

NAND3xp33_ASAP7_75t_L g2690 ( 
.A(n_2660),
.B(n_2550),
.C(n_2552),
.Y(n_2690)
);

NOR3xp33_ASAP7_75t_SL g2691 ( 
.A(n_2633),
.B(n_2631),
.C(n_2612),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2630),
.Y(n_2692)
);

NOR3xp33_ASAP7_75t_L g2693 ( 
.A(n_2624),
.B(n_2608),
.C(n_2556),
.Y(n_2693)
);

INVxp67_ASAP7_75t_L g2694 ( 
.A(n_2618),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2662),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2649),
.B(n_2602),
.Y(n_2696)
);

NOR2xp67_ASAP7_75t_L g2697 ( 
.A(n_2662),
.B(n_164),
.Y(n_2697)
);

NOR2x1_ASAP7_75t_L g2698 ( 
.A(n_2651),
.B(n_165),
.Y(n_2698)
);

O2A1O1Ixp33_ASAP7_75t_L g2699 ( 
.A1(n_2637),
.A2(n_165),
.B(n_166),
.C(n_168),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2622),
.B(n_169),
.Y(n_2700)
);

XNOR2xp5_ASAP7_75t_L g2701 ( 
.A(n_2664),
.B(n_169),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2638),
.B(n_170),
.Y(n_2702)
);

BUFx4f_ASAP7_75t_SL g2703 ( 
.A(n_2619),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2641),
.B(n_171),
.Y(n_2704)
);

NAND2xp33_ASAP7_75t_SL g2705 ( 
.A(n_2625),
.B(n_172),
.Y(n_2705)
);

NAND3xp33_ASAP7_75t_L g2706 ( 
.A(n_2641),
.B(n_2616),
.C(n_2637),
.Y(n_2706)
);

BUFx6f_ASAP7_75t_L g2707 ( 
.A(n_2618),
.Y(n_2707)
);

AOI211x1_ASAP7_75t_L g2708 ( 
.A1(n_2657),
.A2(n_2614),
.B(n_2636),
.C(n_2628),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2665),
.Y(n_2709)
);

AOI211xp5_ASAP7_75t_SL g2710 ( 
.A1(n_2670),
.A2(n_2627),
.B(n_2661),
.C(n_2659),
.Y(n_2710)
);

NAND3xp33_ASAP7_75t_SL g2711 ( 
.A(n_2678),
.B(n_2625),
.C(n_2656),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2689),
.Y(n_2712)
);

AOI21xp33_ASAP7_75t_SL g2713 ( 
.A1(n_2706),
.A2(n_2684),
.B(n_2680),
.Y(n_2713)
);

NOR2xp33_ASAP7_75t_L g2714 ( 
.A(n_2703),
.B(n_2639),
.Y(n_2714)
);

NAND5xp2_ASAP7_75t_L g2715 ( 
.A(n_2685),
.B(n_2677),
.C(n_2693),
.D(n_2688),
.E(n_2691),
.Y(n_2715)
);

OAI22xp5_ASAP7_75t_L g2716 ( 
.A1(n_2672),
.A2(n_2615),
.B1(n_2658),
.B2(n_2655),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2673),
.B(n_2642),
.Y(n_2717)
);

AOI221xp5_ASAP7_75t_L g2718 ( 
.A1(n_2676),
.A2(n_2690),
.B1(n_2681),
.B2(n_2673),
.C(n_2680),
.Y(n_2718)
);

NOR2xp33_ASAP7_75t_R g2719 ( 
.A(n_2705),
.B(n_2643),
.Y(n_2719)
);

A2O1A1Ixp33_ASAP7_75t_L g2720 ( 
.A1(n_2699),
.A2(n_2654),
.B(n_2647),
.C(n_2646),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2682),
.Y(n_2721)
);

A2O1A1Ixp33_ASAP7_75t_L g2722 ( 
.A1(n_2676),
.A2(n_2642),
.B(n_2663),
.C(n_176),
.Y(n_2722)
);

O2A1O1Ixp33_ASAP7_75t_L g2723 ( 
.A1(n_2669),
.A2(n_173),
.B(n_174),
.C(n_177),
.Y(n_2723)
);

AOI22xp5_ASAP7_75t_L g2724 ( 
.A1(n_2668),
.A2(n_174),
.B1(n_177),
.B2(n_178),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2692),
.Y(n_2725)
);

OAI321xp33_ASAP7_75t_L g2726 ( 
.A1(n_2667),
.A2(n_179),
.A3(n_181),
.B1(n_182),
.B2(n_183),
.C(n_184),
.Y(n_2726)
);

CKINVDCx5p33_ASAP7_75t_R g2727 ( 
.A(n_2701),
.Y(n_2727)
);

AOI21xp33_ASAP7_75t_L g2728 ( 
.A1(n_2671),
.A2(n_179),
.B(n_181),
.Y(n_2728)
);

AOI221xp5_ASAP7_75t_L g2729 ( 
.A1(n_2681),
.A2(n_2708),
.B1(n_2707),
.B2(n_2694),
.C(n_2675),
.Y(n_2729)
);

AOI32xp33_ASAP7_75t_L g2730 ( 
.A1(n_2698),
.A2(n_184),
.A3(n_185),
.B1(n_186),
.B2(n_189),
.Y(n_2730)
);

AOI211xp5_ASAP7_75t_L g2731 ( 
.A1(n_2679),
.A2(n_185),
.B(n_189),
.C(n_190),
.Y(n_2731)
);

AOI221xp5_ASAP7_75t_L g2732 ( 
.A1(n_2707),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.C(n_193),
.Y(n_2732)
);

AOI211x1_ASAP7_75t_L g2733 ( 
.A1(n_2696),
.A2(n_192),
.B(n_196),
.C(n_197),
.Y(n_2733)
);

AOI211xp5_ASAP7_75t_L g2734 ( 
.A1(n_2686),
.A2(n_198),
.B(n_199),
.C(n_200),
.Y(n_2734)
);

AOI222xp33_ASAP7_75t_L g2735 ( 
.A1(n_2707),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.C1(n_203),
.C2(n_204),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2666),
.Y(n_2736)
);

AOI211xp5_ASAP7_75t_L g2737 ( 
.A1(n_2683),
.A2(n_202),
.B(n_203),
.C(n_205),
.Y(n_2737)
);

AOI221xp5_ASAP7_75t_L g2738 ( 
.A1(n_2687),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.C(n_209),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2695),
.Y(n_2739)
);

AOI221xp5_ASAP7_75t_L g2740 ( 
.A1(n_2709),
.A2(n_208),
.B1(n_211),
.B2(n_213),
.C(n_216),
.Y(n_2740)
);

AOI22xp5_ASAP7_75t_L g2741 ( 
.A1(n_2697),
.A2(n_211),
.B1(n_217),
.B2(n_218),
.Y(n_2741)
);

OAI221xp5_ASAP7_75t_L g2742 ( 
.A1(n_2704),
.A2(n_2674),
.B1(n_2702),
.B2(n_2700),
.C(n_221),
.Y(n_2742)
);

O2A1O1Ixp33_ASAP7_75t_L g2743 ( 
.A1(n_2680),
.A2(n_217),
.B(n_219),
.C(n_220),
.Y(n_2743)
);

HB1xp67_ASAP7_75t_L g2744 ( 
.A(n_2719),
.Y(n_2744)
);

AND2x2_ASAP7_75t_L g2745 ( 
.A(n_2736),
.B(n_220),
.Y(n_2745)
);

OAI211xp5_ASAP7_75t_L g2746 ( 
.A1(n_2718),
.A2(n_221),
.B(n_223),
.C(n_224),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2717),
.Y(n_2747)
);

AOI221xp5_ASAP7_75t_L g2748 ( 
.A1(n_2713),
.A2(n_2715),
.B1(n_2716),
.B2(n_2729),
.C(n_2711),
.Y(n_2748)
);

HB1xp67_ASAP7_75t_L g2749 ( 
.A(n_2727),
.Y(n_2749)
);

CKINVDCx5p33_ASAP7_75t_R g2750 ( 
.A(n_2741),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2722),
.B(n_2712),
.Y(n_2751)
);

OAI22xp5_ASAP7_75t_L g2752 ( 
.A1(n_2742),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_2752)
);

NOR2xp33_ASAP7_75t_L g2753 ( 
.A(n_2714),
.B(n_226),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2721),
.B(n_228),
.Y(n_2754)
);

AOI221x1_ASAP7_75t_L g2755 ( 
.A1(n_2725),
.A2(n_230),
.B1(n_1474),
.B2(n_1414),
.C(n_1390),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2733),
.B(n_241),
.Y(n_2756)
);

XNOR2x1_ASAP7_75t_L g2757 ( 
.A(n_2724),
.B(n_242),
.Y(n_2757)
);

AOI221xp5_ASAP7_75t_L g2758 ( 
.A1(n_2720),
.A2(n_1344),
.B1(n_1334),
.B2(n_1390),
.C(n_1474),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2739),
.Y(n_2759)
);

AOI221xp5_ASAP7_75t_L g2760 ( 
.A1(n_2743),
.A2(n_1474),
.B1(n_1414),
.B2(n_251),
.C(n_255),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2723),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2731),
.Y(n_2762)
);

AOI221xp5_ASAP7_75t_L g2763 ( 
.A1(n_2726),
.A2(n_1414),
.B1(n_249),
.B2(n_256),
.C(n_257),
.Y(n_2763)
);

OAI21x1_ASAP7_75t_L g2764 ( 
.A1(n_2738),
.A2(n_1580),
.B(n_1569),
.Y(n_2764)
);

AND2x6_ASAP7_75t_L g2765 ( 
.A(n_2710),
.B(n_243),
.Y(n_2765)
);

OAI22xp5_ASAP7_75t_L g2766 ( 
.A1(n_2748),
.A2(n_2737),
.B1(n_2734),
.B2(n_2730),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2749),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2744),
.B(n_2728),
.Y(n_2768)
);

AND2x4_ASAP7_75t_L g2769 ( 
.A(n_2745),
.B(n_2728),
.Y(n_2769)
);

OAI211xp5_ASAP7_75t_L g2770 ( 
.A1(n_2746),
.A2(n_2761),
.B(n_2751),
.C(n_2755),
.Y(n_2770)
);

NAND4xp75_ASAP7_75t_L g2771 ( 
.A(n_2747),
.B(n_2740),
.C(n_2732),
.D(n_2735),
.Y(n_2771)
);

NAND4xp75_ASAP7_75t_L g2772 ( 
.A(n_2762),
.B(n_258),
.C(n_260),
.D(n_262),
.Y(n_2772)
);

NAND3xp33_ASAP7_75t_L g2773 ( 
.A(n_2752),
.B(n_267),
.C(n_268),
.Y(n_2773)
);

NOR2x1_ASAP7_75t_L g2774 ( 
.A(n_2754),
.B(n_270),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2759),
.Y(n_2775)
);

CKINVDCx5p33_ASAP7_75t_R g2776 ( 
.A(n_2750),
.Y(n_2776)
);

CKINVDCx5p33_ASAP7_75t_R g2777 ( 
.A(n_2753),
.Y(n_2777)
);

NAND3xp33_ASAP7_75t_SL g2778 ( 
.A(n_2763),
.B(n_271),
.C(n_272),
.Y(n_2778)
);

BUFx2_ASAP7_75t_L g2779 ( 
.A(n_2765),
.Y(n_2779)
);

NOR5xp2_ASAP7_75t_L g2780 ( 
.A(n_2765),
.B(n_275),
.C(n_277),
.D(n_287),
.E(n_288),
.Y(n_2780)
);

AND2x2_ASAP7_75t_L g2781 ( 
.A(n_2757),
.B(n_291),
.Y(n_2781)
);

OAI22xp5_ASAP7_75t_L g2782 ( 
.A1(n_2776),
.A2(n_2767),
.B1(n_2777),
.B2(n_2773),
.Y(n_2782)
);

NAND4xp75_ASAP7_75t_L g2783 ( 
.A(n_2768),
.B(n_2758),
.C(n_2760),
.D(n_2756),
.Y(n_2783)
);

NOR3xp33_ASAP7_75t_L g2784 ( 
.A(n_2770),
.B(n_2764),
.C(n_2765),
.Y(n_2784)
);

AOI22xp33_ASAP7_75t_SL g2785 ( 
.A1(n_2779),
.A2(n_2765),
.B1(n_293),
.B2(n_296),
.Y(n_2785)
);

AOI221xp5_ASAP7_75t_L g2786 ( 
.A1(n_2766),
.A2(n_292),
.B1(n_298),
.B2(n_299),
.C(n_300),
.Y(n_2786)
);

OAI211xp5_ASAP7_75t_L g2787 ( 
.A1(n_2775),
.A2(n_301),
.B(n_304),
.C(n_310),
.Y(n_2787)
);

OAI22xp5_ASAP7_75t_L g2788 ( 
.A1(n_2773),
.A2(n_1092),
.B1(n_1083),
.B2(n_1081),
.Y(n_2788)
);

OAI21xp33_ASAP7_75t_L g2789 ( 
.A1(n_2769),
.A2(n_1092),
.B(n_1083),
.Y(n_2789)
);

OR2x6_ASAP7_75t_L g2790 ( 
.A(n_2774),
.B(n_1092),
.Y(n_2790)
);

INVxp33_ASAP7_75t_SL g2791 ( 
.A(n_2771),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_SL g2792 ( 
.A(n_2785),
.B(n_2769),
.Y(n_2792)
);

AOI221xp5_ASAP7_75t_L g2793 ( 
.A1(n_2791),
.A2(n_2778),
.B1(n_2781),
.B2(n_2780),
.C(n_2772),
.Y(n_2793)
);

XNOR2xp5_ASAP7_75t_L g2794 ( 
.A(n_2782),
.B(n_313),
.Y(n_2794)
);

CKINVDCx5p33_ASAP7_75t_R g2795 ( 
.A(n_2790),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2790),
.Y(n_2796)
);

INVx2_ASAP7_75t_SL g2797 ( 
.A(n_2788),
.Y(n_2797)
);

AOI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2784),
.A2(n_1081),
.B1(n_1083),
.B2(n_1092),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2792),
.Y(n_2799)
);

OAI22xp5_ASAP7_75t_L g2800 ( 
.A1(n_2794),
.A2(n_2783),
.B1(n_2786),
.B2(n_2787),
.Y(n_2800)
);

OA22x2_ASAP7_75t_L g2801 ( 
.A1(n_2795),
.A2(n_2789),
.B1(n_320),
.B2(n_330),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2796),
.Y(n_2802)
);

NOR3xp33_ASAP7_75t_L g2803 ( 
.A(n_2793),
.B(n_315),
.C(n_335),
.Y(n_2803)
);

OR3x1_ASAP7_75t_L g2804 ( 
.A(n_2797),
.B(n_336),
.C(n_338),
.Y(n_2804)
);

HB1xp67_ASAP7_75t_L g2805 ( 
.A(n_2804),
.Y(n_2805)
);

XNOR2xp5_ASAP7_75t_L g2806 ( 
.A(n_2800),
.B(n_2798),
.Y(n_2806)
);

OAI22xp5_ASAP7_75t_L g2807 ( 
.A1(n_2799),
.A2(n_1083),
.B1(n_1081),
.B2(n_1069),
.Y(n_2807)
);

OAI22x1_ASAP7_75t_L g2808 ( 
.A1(n_2802),
.A2(n_340),
.B1(n_341),
.B2(n_345),
.Y(n_2808)
);

OAI22xp5_ASAP7_75t_SL g2809 ( 
.A1(n_2801),
.A2(n_347),
.B1(n_349),
.B2(n_350),
.Y(n_2809)
);

CKINVDCx20_ASAP7_75t_R g2810 ( 
.A(n_2805),
.Y(n_2810)
);

AOI22xp33_ASAP7_75t_L g2811 ( 
.A1(n_2809),
.A2(n_2803),
.B1(n_1081),
.B2(n_1069),
.Y(n_2811)
);

AND2x2_ASAP7_75t_L g2812 ( 
.A(n_2806),
.B(n_351),
.Y(n_2812)
);

AOI22xp5_ASAP7_75t_L g2813 ( 
.A1(n_2807),
.A2(n_2808),
.B1(n_1069),
.B2(n_1068),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2805),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_SL g2815 ( 
.A(n_2814),
.B(n_1069),
.Y(n_2815)
);

INVx1_ASAP7_75t_SL g2816 ( 
.A(n_2810),
.Y(n_2816)
);

INVx4_ASAP7_75t_L g2817 ( 
.A(n_2816),
.Y(n_2817)
);

AOI21xp5_ASAP7_75t_L g2818 ( 
.A1(n_2815),
.A2(n_2812),
.B(n_2811),
.Y(n_2818)
);

AOI22xp33_ASAP7_75t_L g2819 ( 
.A1(n_2817),
.A2(n_2813),
.B1(n_1068),
.B2(n_1056),
.Y(n_2819)
);

OAI22xp33_ASAP7_75t_L g2820 ( 
.A1(n_2818),
.A2(n_354),
.B1(n_355),
.B2(n_358),
.Y(n_2820)
);

OAI221xp5_ASAP7_75t_R g2821 ( 
.A1(n_2819),
.A2(n_360),
.B1(n_365),
.B2(n_368),
.C(n_374),
.Y(n_2821)
);

AOI211xp5_ASAP7_75t_L g2822 ( 
.A1(n_2821),
.A2(n_2820),
.B(n_379),
.C(n_380),
.Y(n_2822)
);


endmodule