module fake_jpeg_15884_n_355 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_355);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_29),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_0),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_51),
.Y(n_71)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_0),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_52),
.Y(n_63)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_37),
.B1(n_28),
.B2(n_20),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_55),
.A2(n_43),
.B1(n_53),
.B2(n_50),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_29),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_37),
.B1(n_28),
.B2(n_36),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_35),
.Y(n_102)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_36),
.B1(n_31),
.B2(n_21),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_32),
.Y(n_113)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_71),
.B(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_79),
.B(n_80),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

AO22x2_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_49),
.B1(n_48),
.B2(n_45),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_83),
.A2(n_63),
.B1(n_66),
.B2(n_39),
.Y(n_131)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_69),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_92),
.Y(n_120)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_89),
.B(n_95),
.Y(n_132)
);

AO22x1_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_49),
.B1(n_48),
.B2(n_45),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_110),
.B1(n_57),
.B2(n_74),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_94),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_106),
.B1(n_61),
.B2(n_67),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_62),
.B(n_31),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_99),
.Y(n_138)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_56),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_105),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_102),
.B(n_33),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_34),
.B(n_29),
.C(n_22),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_113),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_72),
.Y(n_105)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_63),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_108),
.Y(n_143)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_109),
.Y(n_119)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_115),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_57),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_124),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_106),
.B1(n_85),
.B2(n_97),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_66),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_127),
.A2(n_131),
.B1(n_43),
.B2(n_104),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_22),
.B(n_25),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_128),
.A2(n_130),
.B(n_145),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_114),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_74),
.B(n_22),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_88),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_136),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_22),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_83),
.B(n_41),
.C(n_38),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_38),
.C(n_112),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_99),
.B1(n_115),
.B2(n_82),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_90),
.B(n_41),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_110),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_83),
.A2(n_25),
.B(n_1),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_147),
.B(n_111),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_148),
.B(n_160),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_152),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_83),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_130),
.C(n_128),
.Y(n_182)
);

BUFx24_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_156),
.A2(n_174),
.B1(n_176),
.B2(n_119),
.Y(n_213)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_161),
.Y(n_206)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_165),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_164),
.A2(n_170),
.B(n_178),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_143),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_86),
.B1(n_91),
.B2(n_107),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_167),
.A2(n_168),
.B1(n_119),
.B2(n_140),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_91),
.B1(n_108),
.B2(n_109),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_0),
.B(n_1),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_L g171 ( 
.A1(n_120),
.A2(n_13),
.B(n_15),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_171),
.A2(n_170),
.B(n_13),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_26),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_179),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_173),
.A2(n_131),
.B1(n_119),
.B2(n_118),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_122),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_177),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

OR2x6_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_33),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_1),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_149),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_180),
.B(n_208),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_181),
.A2(n_203),
.B1(n_178),
.B2(n_131),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_184),
.C(n_187),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_132),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_132),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_120),
.B(n_147),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_189),
.A2(n_195),
.B(n_196),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_152),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_191),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_164),
.A2(n_131),
.B1(n_141),
.B2(n_138),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_193),
.A2(n_212),
.B1(n_179),
.B2(n_176),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_194),
.Y(n_220)
);

XOR2x1_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_126),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_126),
.B(n_138),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_143),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_2),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_125),
.C(n_154),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_210),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_159),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_178),
.A2(n_169),
.B1(n_166),
.B2(n_156),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_10),
.B1(n_12),
.B2(n_7),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_215),
.A2(n_205),
.B1(n_204),
.B2(n_4),
.Y(n_261)
);

AND2x2_ASAP7_75t_SL g217 ( 
.A(n_195),
.B(n_178),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_217),
.A2(n_201),
.B(n_210),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_226),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_221),
.B(n_30),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_172),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_225),
.C(n_228),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_139),
.Y(n_223)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_182),
.A2(n_174),
.B1(n_131),
.B2(n_118),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_224),
.A2(n_231),
.B1(n_241),
.B2(n_205),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_191),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_139),
.C(n_158),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_188),
.C(n_212),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_232),
.C(n_236),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_189),
.B(n_135),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_241),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_183),
.B(n_135),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_33),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_188),
.B(n_32),
.C(n_30),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_209),
.C(n_204),
.Y(n_263)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_238),
.B(n_240),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_181),
.A2(n_32),
.B1(n_30),
.B2(n_19),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_239),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_198),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_185),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_211),
.B(n_8),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_242),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_186),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_246),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_186),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_199),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_254),
.C(n_259),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_248),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_218),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_216),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_266),
.B(n_220),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_193),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_201),
.B(n_192),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_257),
.A2(n_260),
.B(n_264),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_206),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_229),
.A2(n_192),
.B(n_208),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_261),
.A2(n_227),
.B1(n_233),
.B2(n_214),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_224),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_228),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_217),
.A2(n_2),
.B(n_3),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_217),
.A2(n_209),
.B(n_4),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_267),
.B(n_237),
.Y(n_285)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_270),
.A2(n_275),
.B(n_266),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_250),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_271),
.B(n_277),
.Y(n_290)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_272),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_227),
.Y(n_273)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_273),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_236),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_274),
.B(n_276),
.Y(n_296)
);

FAx1_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_231),
.CI(n_221),
.CON(n_275),
.SN(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_214),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_279),
.A2(n_289),
.B(n_262),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_238),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_280),
.B(n_282),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_257),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_255),
.C(n_256),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_243),
.B1(n_265),
.B2(n_263),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_244),
.Y(n_300)
);

XNOR2x2_ASAP7_75t_SL g288 ( 
.A(n_264),
.B(n_225),
.Y(n_288)
);

FAx1_ASAP7_75t_SL g299 ( 
.A(n_288),
.B(n_259),
.CI(n_254),
.CON(n_299),
.SN(n_299)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_260),
.Y(n_289)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_295),
.C(n_303),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_255),
.C(n_247),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_298),
.A2(n_269),
.B1(n_270),
.B2(n_273),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_281),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_301),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_269),
.A2(n_246),
.B(n_267),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_256),
.Y(n_303)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

NOR3xp33_ASAP7_75t_SL g305 ( 
.A(n_288),
.B(n_245),
.C(n_7),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_305),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_19),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_307),
.C(n_285),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_7),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_296),
.B(n_287),
.Y(n_311)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_311),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_297),
.A2(n_279),
.B1(n_278),
.B2(n_275),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_322),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_290),
.B1(n_291),
.B2(n_278),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_315),
.A2(n_319),
.B1(n_299),
.B2(n_4),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_316),
.B(n_321),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_293),
.B(n_275),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_301),
.Y(n_324)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_318),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_280),
.C(n_268),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_3),
.C(n_5),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_277),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_294),
.C(n_300),
.Y(n_328)
);

NAND3xp33_ASAP7_75t_SL g323 ( 
.A(n_309),
.B(n_298),
.C(n_305),
.Y(n_323)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_324),
.B(n_313),
.Y(n_340)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_326),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_308),
.A2(n_306),
.B(n_307),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_327),
.A2(n_328),
.B(n_332),
.Y(n_337)
);

OAI22x1_ASAP7_75t_L g329 ( 
.A1(n_314),
.A2(n_284),
.B1(n_299),
.B2(n_5),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_329),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_310),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_339),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_338),
.A2(n_6),
.B(n_326),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_320),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_340),
.B(n_341),
.Y(n_346)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_333),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_335),
.A2(n_331),
.B(n_325),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_342),
.B(n_343),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_339),
.A2(n_312),
.B(n_328),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_344),
.B(n_332),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_347),
.A2(n_348),
.B(n_346),
.Y(n_350)
);

NOR3xp33_ASAP7_75t_SL g348 ( 
.A(n_345),
.B(n_340),
.C(n_337),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_350),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_349),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_312),
.C(n_336),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_319),
.Y(n_354)
);

AO21x1_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_325),
.B(n_313),
.Y(n_355)
);


endmodule