module fake_aes_733_n_686 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_686);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_686;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_40), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_66), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_46), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_34), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_3), .Y(n_81) );
INVx3_ASAP7_75t_L g82 ( .A(n_76), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_21), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_50), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_21), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_5), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_62), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_52), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_29), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_5), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_28), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_54), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_43), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_14), .Y(n_94) );
CKINVDCx16_ASAP7_75t_R g95 ( .A(n_63), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_64), .Y(n_96) );
INVxp33_ASAP7_75t_L g97 ( .A(n_60), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_72), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_69), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_7), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_67), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_41), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_12), .Y(n_103) );
INVxp33_ASAP7_75t_L g104 ( .A(n_59), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_75), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_73), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_11), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_58), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_9), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_37), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_19), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_45), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_53), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_19), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_22), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_74), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_70), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_25), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_1), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_3), .B(n_36), .Y(n_120) );
INVxp33_ASAP7_75t_L g121 ( .A(n_10), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_38), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_35), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_13), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_85), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_115), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_85), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_95), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g129 ( .A(n_82), .B(n_0), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_85), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_112), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_100), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_112), .Y(n_134) );
CKINVDCx8_ASAP7_75t_R g135 ( .A(n_95), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_82), .B(n_0), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_100), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_100), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_105), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_82), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_105), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_115), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_82), .B(n_1), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_103), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_103), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_110), .B(n_2), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_121), .B(n_2), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_110), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_124), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_84), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_89), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_124), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_124), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_110), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_86), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_117), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_81), .B(n_4), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_77), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_97), .B(n_4), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_108), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_77), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_108), .Y(n_163) );
NOR2xp33_ASAP7_75t_R g164 ( .A(n_79), .B(n_27), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_86), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_79), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_161), .B(n_104), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_136), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_148), .A2(n_114), .B1(n_111), .B2(n_90), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_163), .B(n_116), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_136), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_136), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_136), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_136), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_131), .B(n_116), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_140), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_131), .B(n_80), .Y(n_177) );
BUFx2_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_134), .B(n_80), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_140), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_140), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_135), .B(n_123), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_140), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_140), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_158), .B(n_107), .Y(n_185) );
BUFx2_ASAP7_75t_L g186 ( .A(n_128), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_158), .B(n_107), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_140), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_140), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_155), .Y(n_190) );
NAND2xp33_ASAP7_75t_L g191 ( .A(n_151), .B(n_86), .Y(n_191) );
OAI221xp5_ASAP7_75t_L g192 ( .A1(n_135), .A2(n_114), .B1(n_111), .B2(n_90), .C(n_119), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_148), .A2(n_81), .B1(n_83), .B2(n_119), .Y(n_193) );
INVxp67_ASAP7_75t_SL g194 ( .A(n_148), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_133), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_160), .Y(n_196) );
BUFx2_ASAP7_75t_L g197 ( .A(n_139), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_158), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_133), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_132), .B(n_83), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_149), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_133), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_149), .Y(n_203) );
NAND2x1p5_ASAP7_75t_L g204 ( .A(n_158), .B(n_123), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_160), .B(n_98), .Y(n_205) );
INVxp67_ASAP7_75t_SL g206 ( .A(n_160), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_155), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_133), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_158), .B(n_94), .Y(n_209) );
NOR2x1p5_ASAP7_75t_L g210 ( .A(n_142), .B(n_122), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_165), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_149), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_132), .B(n_94), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_135), .B(n_98), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_165), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_159), .B(n_109), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_155), .Y(n_217) );
AO22x2_ASAP7_75t_L g218 ( .A1(n_129), .A2(n_122), .B1(n_118), .B2(n_113), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_156), .A2(n_109), .B1(n_86), .B2(n_113), .Y(n_219) );
OAI221xp5_ASAP7_75t_L g220 ( .A1(n_159), .A2(n_78), .B1(n_118), .B2(n_106), .C(n_102), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_162), .Y(n_221) );
OR2x2_ASAP7_75t_L g222 ( .A(n_141), .B(n_86), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_152), .B(n_96), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_162), .A2(n_96), .B(n_106), .C(n_102), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_162), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_157), .B(n_92), .Y(n_226) );
BUFx2_ASAP7_75t_L g227 ( .A(n_126), .Y(n_227) );
AND2x4_ASAP7_75t_L g228 ( .A(n_166), .B(n_92), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_221), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_206), .B(n_166), .Y(n_230) );
INVx1_ASAP7_75t_SL g231 ( .A(n_178), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_178), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_194), .B(n_166), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_196), .B(n_137), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_171), .A2(n_137), .B(n_125), .C(n_154), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_196), .A2(n_129), .B1(n_143), .B2(n_147), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_168), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_205), .B(n_164), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_168), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_216), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_192), .A2(n_120), .B1(n_88), .B2(n_91), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_221), .Y(n_242) );
OR2x6_ASAP7_75t_L g243 ( .A(n_204), .B(n_87), .Y(n_243) );
NOR2xp33_ASAP7_75t_R g244 ( .A(n_186), .B(n_87), .Y(n_244) );
INVxp67_ASAP7_75t_SL g245 ( .A(n_204), .Y(n_245) );
NAND2x1p5_ASAP7_75t_L g246 ( .A(n_168), .B(n_88), .Y(n_246) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_186), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_216), .Y(n_248) );
NAND2x1p5_ASAP7_75t_L g249 ( .A(n_213), .B(n_138), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_213), .B(n_164), .Y(n_250) );
INVxp67_ASAP7_75t_L g251 ( .A(n_197), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_213), .B(n_91), .Y(n_252) );
NOR2xp33_ASAP7_75t_R g253 ( .A(n_197), .B(n_93), .Y(n_253) );
AND2x4_ASAP7_75t_SL g254 ( .A(n_213), .B(n_93), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_177), .B(n_144), .Y(n_255) );
OR2x6_ASAP7_75t_L g256 ( .A(n_204), .B(n_99), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_200), .B(n_144), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_225), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_169), .A2(n_99), .B1(n_101), .B2(n_153), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_225), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_200), .B(n_145), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_173), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_227), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_216), .B(n_145), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_185), .B(n_138), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_216), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_227), .Y(n_267) );
NAND2xp33_ASAP7_75t_R g268 ( .A(n_185), .B(n_6), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_175), .B(n_146), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_185), .B(n_101), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_228), .Y(n_271) );
CKINVDCx6p67_ASAP7_75t_R g272 ( .A(n_182), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_228), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_173), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_170), .B(n_146), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_179), .B(n_125), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_185), .B(n_154), .Y(n_277) );
INVx3_ASAP7_75t_L g278 ( .A(n_173), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_198), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_228), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_198), .Y(n_281) );
NOR3xp33_ASAP7_75t_SL g282 ( .A(n_220), .B(n_127), .C(n_130), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_187), .B(n_153), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_210), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_190), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_187), .B(n_209), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_187), .B(n_150), .Y(n_287) );
BUFx4f_ASAP7_75t_L g288 ( .A(n_187), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_209), .B(n_127), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_228), .Y(n_290) );
INVx5_ASAP7_75t_L g291 ( .A(n_198), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_209), .B(n_150), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_190), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_286), .A2(n_171), .B(n_172), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_231), .B(n_169), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_229), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_229), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_242), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_279), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_245), .B(n_209), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_243), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_232), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_249), .B(n_193), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_237), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_279), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_243), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_242), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_232), .B(n_193), .Y(n_308) );
INVx1_ASAP7_75t_SL g309 ( .A(n_247), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_243), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_250), .A2(n_174), .B(n_172), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_249), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_258), .Y(n_313) );
AND2x4_ASAP7_75t_SL g314 ( .A(n_243), .B(n_219), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_281), .A2(n_174), .B(n_198), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_258), .Y(n_316) );
INVx4_ASAP7_75t_L g317 ( .A(n_256), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_260), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_244), .Y(n_319) );
NAND2x1_ASAP7_75t_L g320 ( .A(n_256), .B(n_217), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_256), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_256), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_281), .A2(n_214), .B(n_191), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_285), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_251), .B(n_223), .Y(n_325) );
AOI22xp33_ASAP7_75t_SL g326 ( .A1(n_253), .A2(n_218), .B1(n_226), .B2(n_222), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_254), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_260), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_230), .B(n_210), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_237), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_230), .B(n_190), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_274), .Y(n_332) );
INVx3_ASAP7_75t_SL g333 ( .A(n_263), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_284), .B(n_167), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_274), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_288), .B(n_219), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_237), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_259), .A2(n_218), .B1(n_224), .B2(n_201), .C(n_212), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_254), .B(n_288), .Y(n_339) );
BUFx10_ASAP7_75t_L g340 ( .A(n_265), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_240), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_248), .B(n_222), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_267), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_266), .Y(n_344) );
AOI21x1_ASAP7_75t_L g345 ( .A1(n_311), .A2(n_218), .B(n_189), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_308), .B(n_276), .Y(n_346) );
INVx4_ASAP7_75t_L g347 ( .A(n_306), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_303), .B(n_276), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_317), .A2(n_246), .B1(n_288), .B2(n_218), .Y(n_349) );
OR2x6_ASAP7_75t_L g350 ( .A(n_317), .B(n_246), .Y(n_350) );
OA21x2_ASAP7_75t_L g351 ( .A1(n_315), .A2(n_235), .B(n_189), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_308), .A2(n_265), .B1(n_289), .B2(n_284), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_296), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_300), .B(n_282), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_317), .A2(n_246), .B1(n_235), .B2(n_280), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_295), .A2(n_289), .B1(n_265), .B2(n_263), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_306), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_294), .A2(n_238), .B(n_270), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_295), .A2(n_289), .B1(n_271), .B2(n_273), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_300), .B(n_264), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_309), .B(n_257), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_306), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_317), .A2(n_306), .B1(n_322), .B2(n_321), .Y(n_363) );
NAND2x1_ASAP7_75t_L g364 ( .A(n_306), .B(n_239), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_325), .B(n_261), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_329), .A2(n_275), .B1(n_234), .B2(n_267), .C(n_241), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_300), .B(n_264), .Y(n_367) );
AOI22xp33_ASAP7_75t_SL g368 ( .A1(n_319), .A2(n_268), .B1(n_234), .B2(n_233), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_302), .A2(n_290), .B1(n_278), .B2(n_262), .Y(n_369) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_322), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_300), .B(n_255), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_296), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_312), .B(n_252), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_322), .A2(n_287), .B1(n_283), .B2(n_201), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_314), .A2(n_278), .B1(n_262), .B2(n_239), .Y(n_375) );
OAI21x1_ASAP7_75t_L g376 ( .A1(n_320), .A2(n_184), .B(n_188), .Y(n_376) );
AND2x4_ASAP7_75t_SL g377 ( .A(n_350), .B(n_322), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_346), .B(n_343), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_362), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_368), .A2(n_343), .B1(n_333), .B2(n_326), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_371), .B(n_297), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_356), .A2(n_333), .B1(n_314), .B2(n_301), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_348), .A2(n_301), .B1(n_321), .B2(n_322), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_371), .B(n_297), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_372), .Y(n_385) );
OAI222xp33_ASAP7_75t_L g386 ( .A1(n_349), .A2(n_310), .B1(n_321), .B2(n_320), .C1(n_325), .C2(n_336), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_372), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_346), .A2(n_342), .B1(n_344), .B2(n_341), .Y(n_388) );
OR2x2_ASAP7_75t_L g389 ( .A(n_365), .B(n_298), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_355), .A2(n_298), .B(n_328), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_365), .B(n_341), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_372), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_353), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_366), .A2(n_338), .B1(n_334), .B2(n_269), .C(n_344), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_360), .B(n_307), .Y(n_395) );
BUFx2_ASAP7_75t_L g396 ( .A(n_350), .Y(n_396) );
INVx2_ASAP7_75t_SL g397 ( .A(n_350), .Y(n_397) );
AOI21xp5_ASAP7_75t_SL g398 ( .A1(n_349), .A2(n_310), .B(n_307), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_353), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_359), .A2(n_333), .B1(n_342), .B2(n_130), .C(n_327), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_354), .A2(n_342), .B1(n_313), .B2(n_316), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_361), .Y(n_402) );
OR2x6_ASAP7_75t_L g403 ( .A(n_350), .B(n_313), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_351), .Y(n_404) );
NOR2x1_ASAP7_75t_SL g405 ( .A(n_403), .B(n_350), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_387), .Y(n_406) );
AOI31xp33_ASAP7_75t_L g407 ( .A1(n_380), .A2(n_363), .A3(n_355), .B(n_374), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_385), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_394), .A2(n_352), .B1(n_361), .B2(n_367), .C(n_360), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_394), .B(n_351), .C(n_374), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_388), .A2(n_367), .B1(n_342), .B2(n_369), .C(n_358), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_381), .B(n_316), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_385), .Y(n_413) );
OAI21x1_ASAP7_75t_L g414 ( .A1(n_390), .A2(n_376), .B(n_345), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_381), .B(n_318), .Y(n_415) );
OAI33xp33_ASAP7_75t_L g416 ( .A1(n_402), .A2(n_212), .A3(n_203), .B1(n_363), .B2(n_373), .B3(n_217), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_392), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_387), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_381), .B(n_318), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_378), .A2(n_375), .B1(n_347), .B2(n_357), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_398), .A2(n_328), .B1(n_347), .B2(n_362), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_400), .A2(n_347), .B1(n_357), .B2(n_339), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_403), .A2(n_347), .B1(n_370), .B2(n_362), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_400), .A2(n_357), .B1(n_339), .B2(n_351), .Y(n_424) );
OAI33xp33_ASAP7_75t_L g425 ( .A1(n_399), .A2(n_203), .A3(n_277), .B1(n_292), .B2(n_180), .B3(n_331), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_399), .B(n_351), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_392), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_390), .B(n_364), .C(n_370), .Y(n_428) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_389), .Y(n_429) );
NOR2x1_ASAP7_75t_L g430 ( .A(n_403), .B(n_357), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_403), .Y(n_431) );
OAI33xp33_ASAP7_75t_L g432 ( .A1(n_383), .A2(n_180), .A3(n_335), .B1(n_332), .B2(n_188), .B3(n_184), .Y(n_432) );
AO21x2_ASAP7_75t_L g433 ( .A1(n_404), .A2(n_345), .B(n_376), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_387), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_403), .Y(n_435) );
AOI33xp33_ASAP7_75t_L g436 ( .A1(n_388), .A2(n_236), .A3(n_195), .B1(n_199), .B2(n_188), .B3(n_184), .Y(n_436) );
AOI21xp33_ASAP7_75t_L g437 ( .A1(n_383), .A2(n_364), .B(n_370), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_393), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_393), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_406), .Y(n_440) );
INVx1_ASAP7_75t_SL g441 ( .A(n_406), .Y(n_441) );
INVx2_ASAP7_75t_SL g442 ( .A(n_430), .Y(n_442) );
NAND3xp33_ASAP7_75t_SL g443 ( .A(n_422), .B(n_389), .C(n_382), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_406), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_439), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_408), .B(n_404), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_439), .B(n_393), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_438), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_409), .A2(n_391), .B1(n_395), .B2(n_401), .C(n_386), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_429), .Y(n_450) );
OAI31xp33_ASAP7_75t_SL g451 ( .A1(n_421), .A2(n_384), .A3(n_386), .B(n_395), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_410), .B(n_389), .C(n_401), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_418), .Y(n_453) );
AOI211xp5_ASAP7_75t_SL g454 ( .A1(n_407), .A2(n_384), .B(n_391), .C(n_395), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_421), .B(n_397), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_438), .B(n_403), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_418), .Y(n_457) );
BUFx3_ASAP7_75t_L g458 ( .A(n_439), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_408), .Y(n_459) );
INVx2_ASAP7_75t_SL g460 ( .A(n_430), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_413), .Y(n_461) );
AOI33xp33_ASAP7_75t_L g462 ( .A1(n_420), .A2(n_384), .A3(n_397), .B1(n_377), .B2(n_9), .B3(n_10), .Y(n_462) );
AOI211x1_ASAP7_75t_L g463 ( .A1(n_407), .A2(n_6), .B(n_7), .C(n_8), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_418), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_434), .B(n_396), .Y(n_465) );
NAND4xp25_ASAP7_75t_L g466 ( .A(n_409), .B(n_396), .C(n_165), .D(n_323), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_412), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_434), .B(n_397), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_434), .B(n_377), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_433), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_412), .B(n_377), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_413), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_417), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_415), .B(n_379), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_435), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_433), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_417), .B(n_379), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_415), .B(n_379), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_419), .B(n_272), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_427), .B(n_370), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_419), .Y(n_481) );
AND2x4_ASAP7_75t_SL g482 ( .A(n_431), .B(n_370), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_427), .B(n_370), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_431), .Y(n_484) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_410), .A2(n_165), .B(n_362), .Y(n_485) );
OR2x6_ASAP7_75t_L g486 ( .A(n_435), .B(n_362), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_432), .A2(n_362), .B(n_324), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g488 ( .A1(n_424), .A2(n_304), .B1(n_337), .B2(n_330), .C(n_207), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g489 ( .A1(n_411), .A2(n_304), .B1(n_337), .B2(n_330), .C(n_207), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_467), .B(n_426), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_450), .B(n_431), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_484), .B(n_431), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_484), .B(n_405), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_459), .Y(n_494) );
AND2x4_ASAP7_75t_SL g495 ( .A(n_474), .B(n_405), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_481), .B(n_416), .Y(n_496) );
NOR4xp25_ASAP7_75t_SL g497 ( .A(n_489), .B(n_437), .C(n_411), .D(n_436), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_459), .B(n_426), .Y(n_498) );
AND2x2_ASAP7_75t_SL g499 ( .A(n_451), .B(n_423), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_461), .B(n_423), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_443), .A2(n_425), .B1(n_432), .B2(n_437), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_461), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_472), .B(n_433), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_463), .A2(n_425), .B1(n_428), .B2(n_207), .C(n_176), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_472), .B(n_433), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_451), .B(n_428), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_443), .A2(n_272), .B1(n_337), .B2(n_330), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_473), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_444), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_473), .B(n_8), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_471), .B(n_11), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_471), .B(n_12), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_456), .B(n_13), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_444), .B(n_414), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_456), .B(n_14), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_448), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_474), .B(n_15), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_448), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_445), .B(n_414), .Y(n_519) );
INVx3_ASAP7_75t_L g520 ( .A(n_445), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_484), .B(n_414), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_440), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_447), .B(n_15), .Y(n_523) );
INVx1_ASAP7_75t_SL g524 ( .A(n_478), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_484), .B(n_68), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_478), .B(n_16), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_446), .Y(n_527) );
NAND2xp33_ASAP7_75t_SL g528 ( .A(n_462), .B(n_332), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_446), .Y(n_529) );
INVx1_ASAP7_75t_SL g530 ( .A(n_447), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_477), .B(n_16), .Y(n_531) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_445), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_440), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_440), .Y(n_534) );
OAI31xp33_ASAP7_75t_L g535 ( .A1(n_454), .A2(n_304), .A3(n_18), .B(n_20), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_449), .B(n_17), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g537 ( .A(n_466), .B(n_262), .C(n_239), .Y(n_537) );
INVx3_ASAP7_75t_L g538 ( .A(n_458), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_458), .B(n_17), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_458), .B(n_18), .Y(n_540) );
NAND3xp33_ASAP7_75t_SL g541 ( .A(n_454), .B(n_20), .C(n_22), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_477), .B(n_23), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_449), .B(n_23), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_441), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_480), .B(n_335), .Y(n_545) );
NOR2x1_ASAP7_75t_L g546 ( .A(n_452), .B(n_324), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_535), .A2(n_485), .B(n_455), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_496), .A2(n_479), .B1(n_452), .B2(n_466), .Y(n_548) );
OAI21xp33_ASAP7_75t_L g549 ( .A1(n_499), .A2(n_460), .B(n_442), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_493), .B(n_460), .Y(n_550) );
OAI21xp5_ASAP7_75t_SL g551 ( .A1(n_495), .A2(n_489), .B(n_475), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_524), .B(n_441), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_494), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_530), .B(n_475), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_532), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_527), .B(n_465), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_490), .B(n_457), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_529), .B(n_465), .Y(n_558) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_541), .A2(n_485), .B(n_488), .Y(n_559) );
INVxp67_ASAP7_75t_L g560 ( .A(n_496), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_495), .B(n_469), .Y(n_561) );
OAI32xp33_ASAP7_75t_L g562 ( .A1(n_526), .A2(n_442), .A3(n_460), .B1(n_488), .B2(n_464), .Y(n_562) );
O2A1O1Ixp5_ASAP7_75t_L g563 ( .A1(n_506), .A2(n_476), .B(n_470), .C(n_469), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_499), .B(n_442), .Y(n_564) );
OR3x2_ASAP7_75t_L g565 ( .A(n_513), .B(n_463), .C(n_26), .Y(n_565) );
INVx2_ASAP7_75t_SL g566 ( .A(n_545), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_502), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_508), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_536), .A2(n_468), .B1(n_483), .B2(n_486), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_509), .B(n_464), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_516), .Y(n_571) );
INVxp33_ASAP7_75t_L g572 ( .A(n_517), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_509), .B(n_464), .Y(n_573) );
NOR2xp67_ASAP7_75t_L g574 ( .A(n_520), .B(n_476), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_491), .B(n_453), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_532), .B(n_483), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_518), .B(n_457), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_515), .B(n_457), .Y(n_578) );
OAI22xp33_ASAP7_75t_L g579 ( .A1(n_506), .A2(n_486), .B1(n_453), .B2(n_487), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_539), .B(n_486), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_539), .Y(n_581) );
NAND3xp33_ASAP7_75t_SL g582 ( .A(n_497), .B(n_487), .C(n_470), .Y(n_582) );
O2A1O1Ixp33_ASAP7_75t_L g583 ( .A1(n_543), .A2(n_476), .B(n_470), .C(n_486), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_540), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_540), .B(n_453), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_498), .Y(n_586) );
OAI21xp33_ASAP7_75t_L g587 ( .A1(n_501), .A2(n_486), .B(n_482), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g588 ( .A1(n_510), .A2(n_482), .B1(n_176), .B2(n_181), .C(n_183), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_531), .B(n_482), .Y(n_589) );
O2A1O1Ixp33_ASAP7_75t_L g590 ( .A1(n_511), .A2(n_305), .B(n_299), .C(n_181), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_512), .B(n_520), .Y(n_591) );
AOI322xp5_ASAP7_75t_L g592 ( .A1(n_528), .A2(n_305), .A3(n_299), .B1(n_324), .B2(n_278), .C1(n_291), .C2(n_293), .Y(n_592) );
NAND2x1p5_ASAP7_75t_L g593 ( .A(n_525), .B(n_285), .Y(n_593) );
AOI211xp5_ASAP7_75t_L g594 ( .A1(n_528), .A2(n_24), .B(n_30), .C(n_31), .Y(n_594) );
AND2x4_ASAP7_75t_L g595 ( .A(n_493), .B(n_32), .Y(n_595) );
INVxp67_ASAP7_75t_L g596 ( .A(n_542), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_500), .B(n_33), .Y(n_597) );
NAND3x2_ASAP7_75t_L g598 ( .A(n_591), .B(n_493), .C(n_492), .Y(n_598) );
NOR2xp33_ASAP7_75t_R g599 ( .A(n_582), .B(n_538), .Y(n_599) );
OAI21xp33_ASAP7_75t_L g600 ( .A1(n_560), .A2(n_501), .B(n_505), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_553), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_567), .Y(n_602) );
AOI32xp33_ASAP7_75t_L g603 ( .A1(n_572), .A2(n_546), .A3(n_538), .B1(n_520), .B2(n_525), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_576), .B(n_492), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_561), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_551), .A2(n_523), .B1(n_538), .B2(n_507), .Y(n_606) );
NOR3xp33_ASAP7_75t_SL g607 ( .A(n_549), .B(n_503), .C(n_504), .Y(n_607) );
OAI22xp33_ASAP7_75t_L g608 ( .A1(n_551), .A2(n_544), .B1(n_522), .B2(n_534), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_568), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_586), .B(n_514), .Y(n_610) );
NOR3xp33_ASAP7_75t_SL g611 ( .A(n_564), .B(n_525), .C(n_537), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_580), .B(n_492), .Y(n_612) );
INVxp67_ASAP7_75t_L g613 ( .A(n_566), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_554), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_570), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_550), .B(n_519), .Y(n_616) );
OAI21xp33_ASAP7_75t_L g617 ( .A1(n_587), .A2(n_521), .B(n_514), .Y(n_617) );
INVxp67_ASAP7_75t_L g618 ( .A(n_557), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_596), .A2(n_521), .B1(n_519), .B2(n_544), .C(n_522), .Y(n_619) );
INVxp67_ASAP7_75t_SL g620 ( .A(n_552), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_571), .B(n_534), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_548), .B(n_521), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_556), .B(n_533), .Y(n_623) );
AND2x4_ASAP7_75t_L g624 ( .A(n_550), .B(n_533), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_577), .Y(n_625) );
INVx1_ASAP7_75t_SL g626 ( .A(n_575), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_589), .B(n_39), .Y(n_627) );
XOR2x2_ASAP7_75t_L g628 ( .A(n_594), .B(n_42), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_558), .B(n_581), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_584), .B(n_44), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_578), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_573), .Y(n_632) );
NAND2x1_ASAP7_75t_L g633 ( .A(n_611), .B(n_574), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_611), .A2(n_563), .B(n_594), .C(n_547), .Y(n_634) );
OAI21xp33_ASAP7_75t_L g635 ( .A1(n_622), .A2(n_569), .B(n_559), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g636 ( .A(n_606), .B(n_583), .C(n_592), .D(n_562), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_622), .A2(n_565), .B1(n_555), .B2(n_595), .Y(n_637) );
NAND2xp33_ASAP7_75t_L g638 ( .A(n_603), .B(n_593), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_600), .B(n_555), .Y(n_639) );
AOI21xp33_ASAP7_75t_SL g640 ( .A1(n_608), .A2(n_617), .B(n_613), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_626), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_607), .A2(n_592), .B1(n_593), .B2(n_590), .C(n_585), .Y(n_642) );
BUFx12f_ASAP7_75t_L g643 ( .A(n_630), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_625), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_601), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g646 ( .A1(n_608), .A2(n_579), .B(n_597), .C(n_595), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_SL g647 ( .A1(n_627), .A2(n_588), .B(n_183), .C(n_195), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_602), .Y(n_648) );
AOI211xp5_ASAP7_75t_SL g649 ( .A1(n_619), .A2(n_293), .B(n_48), .C(n_49), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_598), .A2(n_291), .B1(n_293), .B2(n_285), .Y(n_650) );
OAI21xp33_ASAP7_75t_L g651 ( .A1(n_599), .A2(n_199), .B(n_215), .Y(n_651) );
XNOR2x1_ASAP7_75t_L g652 ( .A(n_605), .B(n_47), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_604), .B(n_51), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_637), .A2(n_618), .B1(n_614), .B2(n_620), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_635), .B(n_609), .Y(n_655) );
INVx2_ASAP7_75t_SL g656 ( .A(n_641), .Y(n_656) );
AND2x2_ASAP7_75t_SL g657 ( .A(n_638), .B(n_624), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_645), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_636), .A2(n_631), .B1(n_610), .B2(n_629), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_644), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_648), .B(n_632), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_640), .B(n_615), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_639), .Y(n_663) );
AOI22x1_ASAP7_75t_L g664 ( .A1(n_649), .A2(n_624), .B1(n_615), .B2(n_599), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_639), .Y(n_665) );
OAI311xp33_ASAP7_75t_L g666 ( .A1(n_634), .A2(n_623), .A3(n_621), .B1(n_607), .C1(n_628), .Y(n_666) );
AOI32xp33_ASAP7_75t_L g667 ( .A1(n_650), .A2(n_624), .A3(n_616), .B1(n_612), .B2(n_627), .Y(n_667) );
OAI211xp5_ASAP7_75t_SL g668 ( .A1(n_646), .A2(n_202), .B(n_211), .C(n_208), .Y(n_668) );
OAI211xp5_ASAP7_75t_SL g669 ( .A1(n_642), .A2(n_202), .B(n_211), .C(n_208), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_650), .A2(n_340), .B1(n_291), .B2(n_285), .Y(n_670) );
OAI22xp5_ASAP7_75t_SL g671 ( .A1(n_643), .A2(n_340), .B1(n_56), .B2(n_57), .Y(n_671) );
OAI311xp33_ASAP7_75t_L g672 ( .A1(n_642), .A2(n_55), .A3(n_61), .B1(n_65), .C1(n_71), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_633), .A2(n_291), .B(n_340), .Y(n_673) );
NOR3xp33_ASAP7_75t_L g674 ( .A(n_651), .B(n_340), .C(n_291), .Y(n_674) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_665), .Y(n_675) );
OAI21xp33_ASAP7_75t_L g676 ( .A1(n_662), .A2(n_659), .B(n_657), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_660), .Y(n_677) );
AOI222xp33_ASAP7_75t_L g678 ( .A1(n_655), .A2(n_665), .B1(n_657), .B2(n_663), .C1(n_654), .C2(n_668), .Y(n_678) );
OAI322xp33_ASAP7_75t_L g679 ( .A1(n_675), .A2(n_655), .A3(n_677), .B1(n_656), .B2(n_678), .C1(n_664), .C2(n_666), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_676), .A2(n_669), .B1(n_671), .B2(n_674), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g681 ( .A(n_678), .B(n_667), .C(n_673), .Y(n_681) );
CKINVDCx11_ASAP7_75t_R g682 ( .A(n_679), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_681), .B(n_658), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_682), .A2(n_680), .B1(n_652), .B2(n_658), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_684), .A2(n_683), .B1(n_661), .B2(n_670), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_685), .A2(n_683), .B1(n_672), .B2(n_653), .C(n_647), .Y(n_686) );
endmodule