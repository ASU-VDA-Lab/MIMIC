module real_aes_8209_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_0), .B(n_86), .C(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g123 ( .A(n_0), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_1), .A2(n_151), .B(n_156), .C(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g263 ( .A(n_2), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_3), .A2(n_146), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_4), .B(n_223), .Y(n_472) );
AOI21xp33_ASAP7_75t_L g224 ( .A1(n_5), .A2(n_146), .B(n_225), .Y(n_224) );
AND2x6_ASAP7_75t_L g151 ( .A(n_6), .B(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_7), .A2(n_145), .B(n_153), .Y(n_144) );
INVx1_ASAP7_75t_L g108 ( .A(n_8), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_8), .B(n_40), .Y(n_124) );
INVx1_ASAP7_75t_L g561 ( .A(n_9), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_10), .B(n_195), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_11), .B(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g230 ( .A(n_12), .Y(n_230) );
INVx1_ASAP7_75t_L g143 ( .A(n_13), .Y(n_143) );
INVx1_ASAP7_75t_L g163 ( .A(n_14), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_15), .A2(n_164), .B(n_178), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_16), .B(n_223), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_17), .B(n_180), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_18), .B(n_146), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_19), .B(n_485), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_20), .A2(n_211), .B(n_237), .C(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_21), .B(n_223), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_22), .B(n_195), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g159 ( .A1(n_23), .A2(n_160), .B(n_162), .C(n_164), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_24), .B(n_195), .Y(n_458) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_25), .Y(n_489) );
INVx1_ASAP7_75t_L g457 ( .A(n_26), .Y(n_457) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_27), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_28), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_29), .B(n_195), .Y(n_264) );
INVx1_ASAP7_75t_L g482 ( .A(n_30), .Y(n_482) );
INVx1_ASAP7_75t_L g242 ( .A(n_31), .Y(n_242) );
INVx2_ASAP7_75t_L g149 ( .A(n_32), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_33), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_34), .A2(n_211), .B(n_231), .C(n_470), .Y(n_469) );
INVxp67_ASAP7_75t_L g483 ( .A(n_35), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_36), .A2(n_151), .B(n_156), .C(n_175), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_37), .A2(n_156), .B(n_456), .C(n_461), .Y(n_455) );
CKINVDCx14_ASAP7_75t_R g468 ( .A(n_38), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_39), .A2(n_67), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_39), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_40), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g240 ( .A(n_41), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_42), .A2(n_182), .B(n_228), .C(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_43), .B(n_195), .Y(n_194) );
OAI22xp5_ASAP7_75t_SL g720 ( .A1(n_44), .A2(n_84), .B1(n_721), .B2(n_722), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_44), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_45), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_46), .Y(n_479) );
INVx1_ASAP7_75t_L g527 ( .A(n_47), .Y(n_527) );
CKINVDCx16_ASAP7_75t_R g243 ( .A(n_48), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_49), .B(n_146), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_50), .A2(n_156), .B1(n_237), .B2(n_239), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_51), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_52), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_53), .A2(n_228), .B(n_229), .C(n_231), .Y(n_227) );
CKINVDCx14_ASAP7_75t_R g558 ( .A(n_54), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_55), .Y(n_199) );
INVx1_ASAP7_75t_L g226 ( .A(n_56), .Y(n_226) );
AOI222xp33_ASAP7_75t_SL g126 ( .A1(n_57), .A2(n_127), .B1(n_130), .B2(n_711), .C1(n_712), .C2(n_713), .Y(n_126) );
INVx1_ASAP7_75t_L g152 ( .A(n_58), .Y(n_152) );
INVx1_ASAP7_75t_L g142 ( .A(n_59), .Y(n_142) );
INVx1_ASAP7_75t_SL g471 ( .A(n_60), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_61), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_62), .B(n_223), .Y(n_531) );
INVx1_ASAP7_75t_L g492 ( .A(n_63), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_SL g250 ( .A1(n_64), .A2(n_180), .B(n_231), .C(n_251), .Y(n_250) );
INVxp67_ASAP7_75t_L g252 ( .A(n_65), .Y(n_252) );
INVx1_ASAP7_75t_L g112 ( .A(n_66), .Y(n_112) );
INVx1_ASAP7_75t_L g129 ( .A(n_67), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_68), .A2(n_146), .B(n_557), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_69), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_70), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_71), .A2(n_146), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g190 ( .A(n_72), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_73), .A2(n_145), .B(n_478), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g454 ( .A(n_74), .Y(n_454) );
INVx1_ASAP7_75t_L g519 ( .A(n_75), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_76), .A2(n_151), .B(n_156), .C(n_193), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_77), .A2(n_146), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g522 ( .A(n_78), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_79), .B(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g140 ( .A(n_80), .Y(n_140) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_81), .A2(n_102), .B1(n_113), .B2(n_724), .Y(n_101) );
INVx1_ASAP7_75t_L g511 ( .A(n_82), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_83), .B(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_84), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_85), .A2(n_151), .B(n_156), .C(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g120 ( .A(n_86), .B(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g443 ( .A(n_86), .Y(n_443) );
OR2x2_ASAP7_75t_L g710 ( .A(n_86), .B(n_122), .Y(n_710) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_87), .A2(n_156), .B(n_491), .C(n_495), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_88), .B(n_139), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_89), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_90), .A2(n_151), .B(n_156), .C(n_208), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_91), .Y(n_216) );
INVx1_ASAP7_75t_L g249 ( .A(n_92), .Y(n_249) );
CKINVDCx16_ASAP7_75t_R g154 ( .A(n_93), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_94), .B(n_177), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_95), .B(n_168), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_96), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_97), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_98), .A2(n_146), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g530 ( .A(n_99), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_100), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx6p67_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_105), .Y(n_725) );
CKINVDCx9p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AOI22x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_126), .B1(n_716), .B2(n_718), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g717 ( .A(n_117), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_118), .A2(n_719), .B(n_723), .Y(n_718) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_125), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_120), .Y(n_723) );
NOR2x2_ASAP7_75t_L g715 ( .A(n_121), .B(n_443), .Y(n_715) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g442 ( .A(n_122), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g711 ( .A(n_127), .Y(n_711) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_440), .B1(n_444), .B2(n_708), .Y(n_130) );
INVx2_ASAP7_75t_SL g131 ( .A(n_132), .Y(n_131) );
OAI22xp5_ASAP7_75t_SL g712 ( .A1(n_132), .A2(n_442), .B1(n_445), .B2(n_710), .Y(n_712) );
OR4x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_336), .C(n_395), .D(n_422), .Y(n_132) );
NAND3xp33_ASAP7_75t_SL g133 ( .A(n_134), .B(n_278), .C(n_303), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_201), .B(n_221), .C(n_254), .Y(n_134) );
AOI211xp5_ASAP7_75t_SL g426 ( .A1(n_135), .A2(n_427), .B(n_429), .C(n_432), .Y(n_426) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_170), .Y(n_135) );
INVx1_ASAP7_75t_L g301 ( .A(n_136), .Y(n_301) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g276 ( .A(n_137), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g308 ( .A(n_137), .Y(n_308) );
AND2x2_ASAP7_75t_L g363 ( .A(n_137), .B(n_332), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_137), .B(n_219), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_137), .B(n_220), .Y(n_421) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g282 ( .A(n_138), .Y(n_282) );
AND2x2_ASAP7_75t_L g325 ( .A(n_138), .B(n_188), .Y(n_325) );
AND2x2_ASAP7_75t_L g343 ( .A(n_138), .B(n_220), .Y(n_343) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_144), .B(n_167), .Y(n_138) );
INVx1_ASAP7_75t_L g200 ( .A(n_139), .Y(n_200) );
INVx2_ASAP7_75t_L g205 ( .A(n_139), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g453 ( .A1(n_139), .A2(n_191), .B(n_454), .C(n_455), .Y(n_453) );
OA21x2_ASAP7_75t_L g555 ( .A1(n_139), .A2(n_556), .B(n_562), .Y(n_555) );
AND2x2_ASAP7_75t_SL g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_L g169 ( .A(n_140), .B(n_141), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
NAND2x1p5_ASAP7_75t_L g191 ( .A(n_147), .B(n_151), .Y(n_191) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
INVx1_ASAP7_75t_L g460 ( .A(n_148), .Y(n_460) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
INVx1_ASAP7_75t_L g238 ( .A(n_149), .Y(n_238) );
INVx1_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
INVx3_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
INVx1_ASAP7_75t_L g180 ( .A(n_150), .Y(n_180) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_150), .Y(n_195) );
INVx4_ASAP7_75t_SL g166 ( .A(n_151), .Y(n_166) );
BUFx3_ASAP7_75t_L g461 ( .A(n_151), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_159), .C(n_166), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_155), .A2(n_166), .B(n_226), .C(n_227), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_155), .A2(n_166), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_155), .A2(n_166), .B(n_468), .C(n_469), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_SL g478 ( .A1(n_155), .A2(n_166), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_SL g518 ( .A1(n_155), .A2(n_166), .B(n_519), .C(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_SL g526 ( .A1(n_155), .A2(n_166), .B(n_527), .C(n_528), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_SL g557 ( .A1(n_155), .A2(n_166), .B(n_558), .C(n_559), .Y(n_557) );
INVx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
BUFx3_ASAP7_75t_L g165 ( .A(n_157), .Y(n_165) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_157), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_160), .B(n_163), .Y(n_162) );
OAI22xp33_ASAP7_75t_L g481 ( .A1(n_160), .A2(n_177), .B1(n_482), .B2(n_483), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_160), .B(n_522), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_160), .B(n_530), .Y(n_529) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI22xp5_ASAP7_75t_SL g239 ( .A1(n_161), .A2(n_240), .B1(n_241), .B2(n_242), .Y(n_239) );
INVx2_ASAP7_75t_L g241 ( .A(n_161), .Y(n_241) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g182 ( .A(n_165), .Y(n_182) );
OAI22xp33_ASAP7_75t_L g235 ( .A1(n_166), .A2(n_191), .B1(n_236), .B2(n_243), .Y(n_235) );
INVx1_ASAP7_75t_L g495 ( .A(n_166), .Y(n_495) );
INVx4_ASAP7_75t_L g187 ( .A(n_168), .Y(n_187) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_168), .A2(n_247), .B(n_253), .Y(n_246) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_168), .Y(n_465) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g184 ( .A(n_169), .Y(n_184) );
INVx4_ASAP7_75t_L g275 ( .A(n_170), .Y(n_275) );
OAI21xp5_ASAP7_75t_L g330 ( .A1(n_170), .A2(n_331), .B(n_333), .Y(n_330) );
AND2x2_ASAP7_75t_L g411 ( .A(n_170), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_188), .Y(n_170) );
INVx1_ASAP7_75t_L g218 ( .A(n_171), .Y(n_218) );
AND2x2_ASAP7_75t_L g280 ( .A(n_171), .B(n_220), .Y(n_280) );
OR2x2_ASAP7_75t_L g309 ( .A(n_171), .B(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g323 ( .A(n_171), .Y(n_323) );
INVx3_ASAP7_75t_L g332 ( .A(n_171), .Y(n_332) );
AND2x2_ASAP7_75t_L g342 ( .A(n_171), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g375 ( .A(n_171), .B(n_281), .Y(n_375) );
AND2x2_ASAP7_75t_L g399 ( .A(n_171), .B(n_355), .Y(n_399) );
OR2x6_ASAP7_75t_L g171 ( .A(n_172), .B(n_185), .Y(n_171) );
AOI21xp5_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_174), .B(n_183), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_179), .B(n_181), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_177), .A2(n_263), .B(n_264), .C(n_265), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g456 ( .A1(n_177), .A2(n_457), .B(n_458), .C(n_459), .Y(n_456) );
INVx5_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_178), .B(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_178), .B(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_178), .B(n_561), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_181), .A2(n_194), .B(n_196), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_181), .A2(n_492), .B(n_493), .C(n_494), .Y(n_491) );
O2A1O1Ixp5_ASAP7_75t_L g510 ( .A1(n_181), .A2(n_493), .B(n_511), .C(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g197 ( .A(n_183), .Y(n_197) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_184), .A2(n_235), .B(n_244), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_184), .B(n_245), .Y(n_244) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_184), .A2(n_259), .B(n_266), .Y(n_258) );
NOR2xp33_ASAP7_75t_SL g185 ( .A(n_186), .B(n_187), .Y(n_185) );
INVx3_ASAP7_75t_L g223 ( .A(n_187), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_187), .B(n_463), .Y(n_462) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_187), .A2(n_488), .B(n_496), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_187), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g220 ( .A(n_188), .Y(n_220) );
AND2x2_ASAP7_75t_L g435 ( .A(n_188), .B(n_277), .Y(n_435) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_197), .B(n_198), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_192), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_191), .A2(n_260), .B(n_261), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_191), .A2(n_489), .B(n_490), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_191), .A2(n_508), .B(n_509), .Y(n_507) );
INVx4_ASAP7_75t_L g211 ( .A(n_195), .Y(n_211) );
INVx2_ASAP7_75t_L g228 ( .A(n_195), .Y(n_228) );
INVx1_ASAP7_75t_L g476 ( .A(n_197), .Y(n_476) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_197), .A2(n_501), .B(n_502), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_200), .B(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_200), .B(n_267), .Y(n_266) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_200), .A2(n_507), .B(n_513), .Y(n_506) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_217), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_203), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g355 ( .A(n_203), .B(n_343), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_203), .B(n_332), .Y(n_417) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g277 ( .A(n_204), .Y(n_277) );
AND2x2_ASAP7_75t_L g281 ( .A(n_204), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g322 ( .A(n_204), .B(n_323), .Y(n_322) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_215), .Y(n_204) );
INVx1_ASAP7_75t_L g485 ( .A(n_205), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_205), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_214), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_212), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_211), .B(n_471), .Y(n_470) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx3_ASAP7_75t_L g231 ( .A(n_213), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_217), .B(n_318), .Y(n_340) );
INVx1_ASAP7_75t_L g379 ( .A(n_217), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_217), .B(n_306), .Y(n_423) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
AND2x2_ASAP7_75t_L g286 ( .A(n_218), .B(n_281), .Y(n_286) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_220), .B(n_277), .Y(n_310) );
INVx1_ASAP7_75t_L g389 ( .A(n_220), .Y(n_389) );
AOI322xp5_ASAP7_75t_L g413 ( .A1(n_221), .A2(n_328), .A3(n_388), .B1(n_414), .B2(n_416), .C1(n_418), .C2(n_420), .Y(n_413) );
AND2x2_ASAP7_75t_SL g221 ( .A(n_222), .B(n_233), .Y(n_221) );
AND2x2_ASAP7_75t_L g268 ( .A(n_222), .B(n_246), .Y(n_268) );
INVx1_ASAP7_75t_SL g271 ( .A(n_222), .Y(n_271) );
AND2x2_ASAP7_75t_L g273 ( .A(n_222), .B(n_234), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_222), .B(n_290), .Y(n_296) );
INVx2_ASAP7_75t_L g315 ( .A(n_222), .Y(n_315) );
AND2x2_ASAP7_75t_L g328 ( .A(n_222), .B(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g366 ( .A(n_222), .B(n_290), .Y(n_366) );
BUFx2_ASAP7_75t_L g383 ( .A(n_222), .Y(n_383) );
AND2x2_ASAP7_75t_L g397 ( .A(n_222), .B(n_257), .Y(n_397) );
OA21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_232), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_233), .B(n_285), .Y(n_312) );
AND2x2_ASAP7_75t_L g439 ( .A(n_233), .B(n_315), .Y(n_439) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_246), .Y(n_233) );
OR2x2_ASAP7_75t_L g284 ( .A(n_234), .B(n_285), .Y(n_284) );
INVx3_ASAP7_75t_L g290 ( .A(n_234), .Y(n_290) );
AND2x2_ASAP7_75t_L g335 ( .A(n_234), .B(n_258), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_234), .B(n_383), .Y(n_382) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_234), .Y(n_419) );
INVx2_ASAP7_75t_L g265 ( .A(n_237), .Y(n_265) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g493 ( .A(n_241), .Y(n_493) );
AND2x2_ASAP7_75t_L g270 ( .A(n_246), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g292 ( .A(n_246), .Y(n_292) );
BUFx2_ASAP7_75t_L g298 ( .A(n_246), .Y(n_298) );
AND2x2_ASAP7_75t_L g317 ( .A(n_246), .B(n_290), .Y(n_317) );
INVx3_ASAP7_75t_L g329 ( .A(n_246), .Y(n_329) );
OR2x2_ASAP7_75t_L g339 ( .A(n_246), .B(n_290), .Y(n_339) );
AOI31xp33_ASAP7_75t_SL g254 ( .A1(n_255), .A2(n_269), .A3(n_272), .B(n_274), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_268), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_256), .B(n_291), .Y(n_302) );
OR2x2_ASAP7_75t_L g326 ( .A(n_256), .B(n_296), .Y(n_326) );
INVx1_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_257), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g347 ( .A(n_257), .B(n_339), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_257), .B(n_329), .Y(n_357) );
AND2x2_ASAP7_75t_L g364 ( .A(n_257), .B(n_365), .Y(n_364) );
NAND2x1_ASAP7_75t_L g392 ( .A(n_257), .B(n_328), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_257), .B(n_383), .Y(n_393) );
AND2x2_ASAP7_75t_L g405 ( .A(n_257), .B(n_290), .Y(n_405) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx3_ASAP7_75t_L g285 ( .A(n_258), .Y(n_285) );
INVx1_ASAP7_75t_L g351 ( .A(n_268), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_268), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_270), .B(n_346), .Y(n_380) );
AND2x4_ASAP7_75t_L g291 ( .A(n_271), .B(n_292), .Y(n_291) );
CKINVDCx16_ASAP7_75t_R g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx2_ASAP7_75t_L g370 ( .A(n_276), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_276), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g318 ( .A(n_277), .B(n_308), .Y(n_318) );
AND2x2_ASAP7_75t_L g412 ( .A(n_277), .B(n_282), .Y(n_412) );
INVx1_ASAP7_75t_L g437 ( .A(n_277), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_283), .B1(n_286), .B2(n_287), .C(n_293), .Y(n_278) );
CKINVDCx14_ASAP7_75t_R g299 ( .A(n_279), .Y(n_299) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_280), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_283), .B(n_334), .Y(n_353) );
INVx3_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g402 ( .A(n_284), .B(n_298), .Y(n_402) );
AND2x2_ASAP7_75t_L g316 ( .A(n_285), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g346 ( .A(n_285), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_285), .B(n_329), .Y(n_374) );
NOR3xp33_ASAP7_75t_L g416 ( .A(n_285), .B(n_386), .C(n_417), .Y(n_416) );
AOI211xp5_ASAP7_75t_SL g349 ( .A1(n_286), .A2(n_350), .B(n_352), .C(n_360), .Y(n_349) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_288), .A2(n_339), .B1(n_340), .B2(n_341), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_289), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_289), .B(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g431 ( .A(n_291), .B(n_405), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_299), .B1(n_300), .B2(n_302), .Y(n_293) );
NOR2xp33_ASAP7_75t_SL g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_297), .B(n_346), .Y(n_377) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_300), .A2(n_392), .B1(n_423), .B2(n_430), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_311), .B1(n_313), .B2(n_318), .C(n_319), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVxp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI221xp5_ASAP7_75t_L g319 ( .A1(n_309), .A2(n_320), .B1(n_326), .B2(n_327), .C(n_330), .Y(n_319) );
INVx1_ASAP7_75t_L g362 ( .A(n_310), .Y(n_362) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_SL g334 ( .A(n_315), .Y(n_334) );
OR2x2_ASAP7_75t_L g407 ( .A(n_315), .B(n_339), .Y(n_407) );
AND2x2_ASAP7_75t_L g409 ( .A(n_315), .B(n_317), .Y(n_409) );
INVx1_ASAP7_75t_L g348 ( .A(n_318), .Y(n_348) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_324), .Y(n_320) );
AOI21xp33_ASAP7_75t_SL g378 ( .A1(n_321), .A2(n_379), .B(n_380), .Y(n_378) );
OR2x2_ASAP7_75t_L g385 ( .A(n_321), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g359 ( .A(n_322), .B(n_343), .Y(n_359) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp33_ASAP7_75t_SL g376 ( .A(n_327), .B(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_328), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_329), .B(n_365), .Y(n_428) );
O2A1O1Ixp33_ASAP7_75t_L g344 ( .A1(n_332), .A2(n_345), .B(n_347), .C(n_348), .Y(n_344) );
NAND2x1_ASAP7_75t_SL g369 ( .A(n_332), .B(n_370), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_333), .A2(n_382), .B1(n_384), .B2(n_387), .Y(n_381) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_335), .B(n_425), .Y(n_424) );
NAND5xp2_ASAP7_75t_L g336 ( .A(n_337), .B(n_349), .C(n_367), .D(n_381), .E(n_390), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_344), .Y(n_337) );
INVx1_ASAP7_75t_L g394 ( .A(n_340), .Y(n_394) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_342), .A2(n_361), .B1(n_401), .B2(n_403), .C(n_406), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_343), .B(n_437), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_346), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_346), .B(n_412), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B1(n_356), .B2(n_358), .Y(n_352) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_364), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
AND2x2_ASAP7_75t_L g434 ( .A(n_363), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_371), .B1(n_375), .B2(n_376), .C(n_378), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g418 ( .A(n_373), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g425 ( .A(n_383), .Y(n_425) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI21xp5_ASAP7_75t_SL g390 ( .A1(n_391), .A2(n_393), .B(n_394), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OAI211xp5_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_398), .B(n_400), .C(n_413), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
A2O1A1Ixp33_ASAP7_75t_L g422 ( .A1(n_398), .A2(n_423), .B(n_424), .C(n_426), .Y(n_422) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_402), .B(n_404), .Y(n_403) );
AOI21xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B(n_410), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_436), .B(n_438), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
XOR2xp5_ASAP7_75t_L g719 ( .A(n_445), .B(n_720), .Y(n_719) );
OR3x1_ASAP7_75t_L g445 ( .A(n_446), .B(n_619), .C(n_666), .Y(n_445) );
NAND3xp33_ASAP7_75t_SL g446 ( .A(n_447), .B(n_565), .C(n_590), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_505), .B1(n_532), .B2(n_535), .C(n_543), .Y(n_447) );
OAI21xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_473), .B(n_498), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_450), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_450), .B(n_548), .Y(n_663) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_464), .Y(n_450) );
AND2x2_ASAP7_75t_L g534 ( .A(n_451), .B(n_504), .Y(n_534) );
AND2x2_ASAP7_75t_L g583 ( .A(n_451), .B(n_503), .Y(n_583) );
AND2x2_ASAP7_75t_L g604 ( .A(n_451), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g609 ( .A(n_451), .B(n_576), .Y(n_609) );
OR2x2_ASAP7_75t_L g617 ( .A(n_451), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g689 ( .A(n_451), .B(n_486), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_451), .B(n_638), .Y(n_703) );
INVx3_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g549 ( .A(n_452), .B(n_464), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_452), .B(n_486), .Y(n_550) );
AND2x4_ASAP7_75t_L g571 ( .A(n_452), .B(n_504), .Y(n_571) );
AND2x2_ASAP7_75t_L g601 ( .A(n_452), .B(n_475), .Y(n_601) );
AND2x2_ASAP7_75t_L g610 ( .A(n_452), .B(n_600), .Y(n_610) );
AND2x2_ASAP7_75t_L g626 ( .A(n_452), .B(n_487), .Y(n_626) );
OR2x2_ASAP7_75t_L g635 ( .A(n_452), .B(n_618), .Y(n_635) );
AND2x2_ASAP7_75t_L g641 ( .A(n_452), .B(n_576), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_452), .B(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g655 ( .A(n_452), .B(n_500), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_452), .B(n_545), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_452), .B(n_605), .Y(n_694) );
OR2x6_ASAP7_75t_L g452 ( .A(n_453), .B(n_462), .Y(n_452) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_460), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g504 ( .A(n_464), .Y(n_504) );
AND2x2_ASAP7_75t_L g600 ( .A(n_464), .B(n_486), .Y(n_600) );
AND2x2_ASAP7_75t_L g605 ( .A(n_464), .B(n_487), .Y(n_605) );
INVx1_ASAP7_75t_L g661 ( .A(n_464), .Y(n_661) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B(n_472), .Y(n_464) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_465), .A2(n_517), .B(n_523), .Y(n_516) );
OA21x2_ASAP7_75t_L g524 ( .A1(n_465), .A2(n_525), .B(n_531), .Y(n_524) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g570 ( .A(n_474), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_486), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_475), .B(n_534), .Y(n_533) );
BUFx3_ASAP7_75t_L g548 ( .A(n_475), .Y(n_548) );
OR2x2_ASAP7_75t_L g618 ( .A(n_475), .B(n_486), .Y(n_618) );
OR2x2_ASAP7_75t_L g679 ( .A(n_475), .B(n_586), .Y(n_679) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B(n_484), .Y(n_475) );
INVx1_ASAP7_75t_L g501 ( .A(n_477), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_484), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_486), .B(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g638 ( .A(n_486), .B(n_500), .Y(n_638) );
INVx2_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g577 ( .A(n_487), .Y(n_577) );
INVx1_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_499), .A2(n_683), .B1(n_687), .B2(n_690), .C(n_691), .Y(n_682) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_503), .Y(n_499) );
INVx1_ASAP7_75t_SL g546 ( .A(n_500), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_500), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g677 ( .A(n_500), .B(n_534), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_503), .B(n_548), .Y(n_669) );
AND2x2_ASAP7_75t_L g576 ( .A(n_504), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_SL g580 ( .A(n_505), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_505), .B(n_586), .Y(n_616) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_515), .Y(n_505) );
AND2x2_ASAP7_75t_L g542 ( .A(n_506), .B(n_516), .Y(n_542) );
INVx4_ASAP7_75t_L g554 ( .A(n_506), .Y(n_554) );
BUFx3_ASAP7_75t_L g596 ( .A(n_506), .Y(n_596) );
AND3x2_ASAP7_75t_L g611 ( .A(n_506), .B(n_612), .C(n_613), .Y(n_611) );
AND2x2_ASAP7_75t_L g693 ( .A(n_515), .B(n_607), .Y(n_693) );
AND2x2_ASAP7_75t_L g701 ( .A(n_515), .B(n_586), .Y(n_701) );
INVx1_ASAP7_75t_SL g706 ( .A(n_515), .Y(n_706) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_524), .Y(n_515) );
INVx1_ASAP7_75t_SL g564 ( .A(n_516), .Y(n_564) );
AND2x2_ASAP7_75t_L g587 ( .A(n_516), .B(n_554), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_516), .B(n_538), .Y(n_589) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_516), .Y(n_629) );
OR2x2_ASAP7_75t_L g634 ( .A(n_516), .B(n_554), .Y(n_634) );
INVx2_ASAP7_75t_L g540 ( .A(n_524), .Y(n_540) );
AND2x2_ASAP7_75t_L g574 ( .A(n_524), .B(n_555), .Y(n_574) );
OR2x2_ASAP7_75t_L g594 ( .A(n_524), .B(n_555), .Y(n_594) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_524), .Y(n_614) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
AOI21xp33_ASAP7_75t_L g664 ( .A1(n_533), .A2(n_573), .B(n_665), .Y(n_664) );
AOI322xp5_ASAP7_75t_L g700 ( .A1(n_535), .A2(n_545), .A3(n_571), .B1(n_701), .B2(n_702), .C1(n_704), .C2(n_707), .Y(n_700) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_537), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_538), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g563 ( .A(n_539), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g631 ( .A(n_540), .B(n_554), .Y(n_631) );
AND2x2_ASAP7_75t_L g698 ( .A(n_540), .B(n_555), .Y(n_698) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g639 ( .A(n_542), .B(n_593), .Y(n_639) );
AOI31xp33_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_547), .A3(n_550), .B(n_551), .Y(n_543) );
AND2x2_ASAP7_75t_L g598 ( .A(n_545), .B(n_576), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_545), .B(n_568), .Y(n_680) );
AND2x2_ASAP7_75t_L g699 ( .A(n_545), .B(n_604), .Y(n_699) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_548), .B(n_576), .Y(n_588) );
NAND2x1p5_ASAP7_75t_L g622 ( .A(n_548), .B(n_605), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_548), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_548), .B(n_689), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_549), .B(n_605), .Y(n_637) );
INVx1_ASAP7_75t_L g681 ( .A(n_549), .Y(n_681) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_563), .Y(n_552) );
INVxp67_ASAP7_75t_L g633 ( .A(n_553), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_554), .B(n_564), .Y(n_569) );
INVx1_ASAP7_75t_L g675 ( .A(n_554), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_554), .B(n_652), .Y(n_686) );
BUFx3_ASAP7_75t_L g586 ( .A(n_555), .Y(n_586) );
AND2x2_ASAP7_75t_L g612 ( .A(n_555), .B(n_564), .Y(n_612) );
INVx2_ASAP7_75t_L g652 ( .A(n_555), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_563), .B(n_685), .Y(n_684) );
AOI211xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_570), .B(n_572), .C(n_581), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AOI21xp33_ASAP7_75t_L g615 ( .A1(n_567), .A2(n_616), .B(n_617), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_568), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_568), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g648 ( .A(n_569), .B(n_594), .Y(n_648) );
INVx3_ASAP7_75t_L g579 ( .A(n_571), .Y(n_579) );
OAI22xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_575), .B1(n_578), .B2(n_580), .Y(n_572) );
OAI21xp5_ASAP7_75t_SL g597 ( .A1(n_574), .A2(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g623 ( .A(n_574), .B(n_587), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_574), .B(n_675), .Y(n_674) );
INVxp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g578 ( .A(n_577), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g647 ( .A(n_577), .Y(n_647) );
OAI21xp5_ASAP7_75t_SL g591 ( .A1(n_578), .A2(n_592), .B(n_597), .Y(n_591) );
OAI22xp33_ASAP7_75t_SL g581 ( .A1(n_582), .A2(n_584), .B1(n_588), .B2(n_589), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_583), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g607 ( .A(n_586), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_586), .B(n_629), .Y(n_628) );
NOR3xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_602), .C(n_615), .Y(n_590) );
OAI22xp5_ASAP7_75t_SL g657 ( .A1(n_592), .A2(n_658), .B1(n_662), .B2(n_663), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g662 ( .A(n_594), .B(n_595), .Y(n_662) );
AND2x2_ASAP7_75t_L g670 ( .A(n_595), .B(n_651), .Y(n_670) );
CKINVDCx16_ASAP7_75t_R g595 ( .A(n_596), .Y(n_595) );
O2A1O1Ixp33_ASAP7_75t_SL g678 ( .A1(n_596), .A2(n_679), .B(n_680), .C(n_681), .Y(n_678) );
OR2x2_ASAP7_75t_L g705 ( .A(n_596), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
OAI21xp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_606), .B(n_608), .Y(n_602) );
INVx1_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_604), .A2(n_641), .B(n_642), .C(n_645), .Y(n_640) );
OAI21xp33_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_610), .B(n_611), .Y(n_608) );
AND2x2_ASAP7_75t_L g673 ( .A(n_612), .B(n_631), .Y(n_673) );
INVxp67_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g651 ( .A(n_614), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g656 ( .A(n_616), .Y(n_656) );
NAND3xp33_ASAP7_75t_SL g619 ( .A(n_620), .B(n_640), .C(n_653), .Y(n_619) );
AOI211xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_623), .B(n_624), .C(n_632), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g690 ( .A(n_627), .Y(n_690) );
OR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g650 ( .A(n_629), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_629), .B(n_698), .Y(n_697) );
INVxp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B(n_635), .C(n_636), .Y(n_632) );
INVx2_ASAP7_75t_SL g644 ( .A(n_634), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_635), .A2(n_646), .B1(n_648), .B2(n_649), .Y(n_645) );
OAI21xp33_ASAP7_75t_SL g636 ( .A1(n_637), .A2(n_638), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
AOI211xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_656), .B(n_657), .C(n_664), .Y(n_653) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
INVxp33_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g707 ( .A(n_661), .Y(n_707) );
NAND4xp25_ASAP7_75t_L g666 ( .A(n_667), .B(n_682), .C(n_695), .D(n_700), .Y(n_666) );
AOI211xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_670), .B(n_671), .C(n_678), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_674), .B(n_676), .Y(n_671) );
AOI21xp33_ASAP7_75t_L g691 ( .A1(n_672), .A2(n_692), .B(n_694), .Y(n_691) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_679), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_699), .Y(n_695) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
endmodule