module real_aes_7783_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_1066;
wire n_684;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_635;
wire n_503;
wire n_673;
wire n_386;
wire n_1067;
wire n_518;
wire n_792;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_577;
wire n_580;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_742;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_958;
wire n_677;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_1040;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_1078;
wire n_495;
wire n_892;
wire n_994;
wire n_1072;
wire n_744;
wire n_384;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_532;
wire n_656;
wire n_746;
wire n_1025;
wire n_409;
wire n_860;
wire n_748;
wire n_909;
wire n_523;
wire n_781;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_874;
wire n_796;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_1081;
wire n_973;
wire n_1084;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_1121;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1013;
wire n_737;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_1100;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1103;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_1083;
wire n_727;
wire n_397;
wire n_749;
wire n_385;
wire n_663;
wire n_1056;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1127;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_928;
wire n_637;
wire n_899;
wire n_692;
wire n_789;
wire n_544;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1071;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_1133;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_1114;
wire n_473;
wire n_566;
wire n_719;
wire n_837;
wire n_967;
wire n_871;
wire n_1045;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1097;
wire n_601;
wire n_500;
wire n_1101;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_1119;
wire n_802;
wire n_868;
wire n_877;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g863 ( .A1(n_0), .A2(n_177), .B1(n_601), .B2(n_864), .Y(n_863) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_1), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_2), .B(n_587), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_3), .B(n_692), .Y(n_691) );
XOR2x2_ASAP7_75t_L g825 ( .A(n_4), .B(n_826), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_5), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g1126 ( .A(n_6), .Y(n_1126) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_7), .A2(n_526), .B1(n_570), .B2(n_571), .Y(n_525) );
INVx1_ASAP7_75t_L g571 ( .A(n_7), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_8), .A2(n_287), .B1(n_505), .B2(n_723), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_9), .A2(n_345), .B1(n_743), .B2(n_744), .Y(n_742) );
AOI22xp5_ASAP7_75t_SL g599 ( .A1(n_10), .A2(n_379), .B1(n_600), .B2(n_601), .Y(n_599) );
AO22x2_ASAP7_75t_L g403 ( .A1(n_11), .A2(n_217), .B1(n_404), .B2(n_405), .Y(n_403) );
INVx1_ASAP7_75t_L g1079 ( .A(n_11), .Y(n_1079) );
CKINVDCx20_ASAP7_75t_R g1029 ( .A(n_12), .Y(n_1029) );
AOI22xp5_ASAP7_75t_L g890 ( .A1(n_13), .A2(n_298), .B1(n_433), .B2(n_663), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_14), .A2(n_61), .B1(n_635), .B2(n_918), .Y(n_917) );
AOI22xp5_ASAP7_75t_SL g593 ( .A1(n_15), .A2(n_243), .B1(n_510), .B2(n_594), .Y(n_593) );
AO22x1_ASAP7_75t_L g794 ( .A1(n_16), .A2(n_795), .B1(n_823), .B2(n_824), .Y(n_794) );
INVx1_ASAP7_75t_L g823 ( .A(n_16), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_17), .A2(n_105), .B1(n_701), .B2(n_928), .Y(n_927) );
CKINVDCx20_ASAP7_75t_R g1011 ( .A(n_18), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_19), .A2(n_25), .B1(n_505), .B2(n_751), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_20), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_21), .A2(n_381), .B1(n_617), .B2(n_718), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_22), .A2(n_374), .B1(n_613), .B2(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g949 ( .A(n_23), .Y(n_949) );
AOI22xp5_ASAP7_75t_L g832 ( .A1(n_24), .A2(n_371), .B1(n_470), .B2(n_833), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_26), .A2(n_266), .B1(n_537), .B2(n_780), .Y(n_948) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_27), .A2(n_332), .B1(n_427), .B2(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g841 ( .A(n_28), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_29), .A2(n_88), .B1(n_517), .B2(n_658), .Y(n_1122) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_30), .A2(n_179), .B1(n_590), .B2(n_591), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_31), .A2(n_338), .B1(n_472), .B2(n_716), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_32), .A2(n_93), .B1(n_434), .B2(n_659), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_33), .A2(n_108), .B1(n_546), .B2(n_548), .Y(n_545) );
AOI22xp33_ASAP7_75t_SL g930 ( .A1(n_34), .A2(n_54), .B1(n_475), .B2(n_509), .Y(n_930) );
AO22x2_ASAP7_75t_L g407 ( .A1(n_35), .A2(n_114), .B1(n_404), .B2(n_408), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_36), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_37), .A2(n_201), .B1(n_613), .B2(n_738), .Y(n_1092) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_38), .A2(n_99), .B1(n_635), .B2(n_658), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_39), .Y(n_803) );
AOI22xp33_ASAP7_75t_SL g865 ( .A1(n_40), .A2(n_320), .B1(n_546), .B2(n_680), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_41), .A2(n_223), .B1(n_488), .B2(n_490), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g1048 ( .A(n_42), .Y(n_1048) );
CKINVDCx20_ASAP7_75t_R g1054 ( .A(n_43), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_44), .B(n_665), .Y(n_921) );
AOI22xp33_ASAP7_75t_SL g936 ( .A1(n_45), .A2(n_272), .B1(n_467), .B2(n_597), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_46), .A2(n_227), .B1(n_490), .B2(n_744), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_47), .B(n_767), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_48), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g1051 ( .A(n_49), .Y(n_1051) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_50), .Y(n_812) );
AOI22xp33_ASAP7_75t_SL g854 ( .A1(n_51), .A2(n_196), .B1(n_581), .B2(n_767), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_52), .A2(n_151), .B1(n_478), .B2(n_510), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_53), .A2(n_362), .B1(n_672), .B2(n_926), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_55), .B(n_754), .Y(n_1027) );
AOI22xp33_ASAP7_75t_SL g700 ( .A1(n_56), .A2(n_317), .B1(n_600), .B2(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_SL g450 ( .A1(n_57), .A2(n_326), .B1(n_451), .B2(n_456), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_58), .A2(n_213), .B1(n_616), .B2(n_617), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_59), .A2(n_190), .B1(n_538), .B2(n_613), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_60), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_62), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_63), .A2(n_365), .B1(n_537), .B2(n_883), .Y(n_899) );
AOI22xp33_ASAP7_75t_SL g898 ( .A1(n_64), .A2(n_294), .B1(n_494), .B2(n_780), .Y(n_898) );
AOI22xp5_ASAP7_75t_SL g394 ( .A1(n_65), .A2(n_395), .B1(n_482), .B2(n_483), .Y(n_394) );
CKINVDCx16_ASAP7_75t_R g483 ( .A(n_65), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g1121 ( .A(n_66), .Y(n_1121) );
INVx1_ASAP7_75t_L g605 ( .A(n_67), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_68), .A2(n_109), .B1(n_621), .B2(n_818), .Y(n_817) );
AOI222xp33_ASAP7_75t_L g513 ( .A1(n_69), .A2(n_205), .B1(n_237), .B2(n_514), .C1(n_515), .C2(n_517), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_70), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_71), .Y(n_568) );
AOI22xp33_ASAP7_75t_SL g869 ( .A1(n_72), .A2(n_269), .B1(n_604), .B2(n_833), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_73), .A2(n_279), .B1(n_509), .B2(n_603), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_74), .A2(n_98), .B1(n_604), .B2(n_1089), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_75), .A2(n_254), .B1(n_428), .B2(n_503), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_76), .A2(n_230), .B1(n_488), .B2(n_928), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_77), .A2(n_164), .B1(n_594), .B2(n_601), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_78), .Y(n_530) );
AOI22xp5_ASAP7_75t_SL g595 ( .A1(n_79), .A2(n_251), .B1(n_478), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_SL g922 ( .A1(n_80), .A2(n_224), .B1(n_659), .B2(n_694), .Y(n_922) );
CKINVDCx20_ASAP7_75t_R g996 ( .A(n_81), .Y(n_996) );
AOI22xp33_ASAP7_75t_SL g474 ( .A1(n_82), .A2(n_134), .B1(n_475), .B2(n_478), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_83), .A2(n_120), .B1(n_509), .B2(n_510), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g940 ( .A(n_84), .Y(n_940) );
AO22x2_ASAP7_75t_L g411 ( .A1(n_85), .A2(n_260), .B1(n_404), .B2(n_405), .Y(n_411) );
INVx1_ASAP7_75t_L g1076 ( .A(n_85), .Y(n_1076) );
CKINVDCx20_ASAP7_75t_R g1101 ( .A(n_86), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_87), .A2(n_257), .B1(n_479), .B2(n_1044), .Y(n_1043) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_89), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_90), .A2(n_186), .B1(n_505), .B2(n_694), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_91), .A2(n_283), .B1(n_463), .B2(n_509), .Y(n_1133) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_92), .A2(n_314), .B1(n_671), .B2(n_673), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_94), .A2(n_377), .B1(n_475), .B2(n_668), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_95), .Y(n_533) );
AOI22xp5_ASAP7_75t_SL g602 ( .A1(n_96), .A2(n_210), .B1(n_603), .B2(n_604), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_97), .A2(n_295), .B1(n_475), .B2(n_512), .Y(n_511) );
AOI211xp5_ASAP7_75t_L g674 ( .A1(n_100), .A2(n_594), .B(n_675), .C(n_681), .Y(n_674) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_101), .A2(n_285), .B1(n_662), .B2(n_663), .Y(n_661) );
AOI222xp33_ASAP7_75t_L g884 ( .A1(n_102), .A2(n_229), .B1(n_240), .B2(n_514), .C1(n_517), .C2(n_663), .Y(n_884) );
INVx1_ASAP7_75t_L g1061 ( .A(n_103), .Y(n_1061) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_104), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g979 ( .A(n_106), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_107), .A2(n_197), .B1(n_433), .B2(n_505), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_110), .A2(n_204), .B1(n_692), .B2(n_749), .Y(n_1104) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_111), .A2(n_608), .B1(n_641), .B2(n_642), .Y(n_607) );
INVx1_ASAP7_75t_L g641 ( .A(n_111), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_112), .A2(n_119), .B1(n_515), .B2(n_517), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_113), .A2(n_182), .B1(n_503), .B2(n_558), .Y(n_728) );
INVx1_ASAP7_75t_L g1080 ( .A(n_114), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_115), .A2(n_249), .B1(n_512), .B2(n_718), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_116), .B(n_634), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g1004 ( .A(n_117), .Y(n_1004) );
XOR2xp5_ASAP7_75t_L g873 ( .A(n_118), .B(n_874), .Y(n_873) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_121), .A2(n_328), .B1(n_503), .B2(n_505), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g867 ( .A1(n_122), .A2(n_199), .B1(n_451), .B2(n_868), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_123), .A2(n_354), .B1(n_668), .B2(n_743), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_124), .B(n_499), .Y(n_943) );
CKINVDCx20_ASAP7_75t_R g1047 ( .A(n_125), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_126), .A2(n_191), .B1(n_535), .B2(n_538), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_127), .A2(n_277), .B1(n_451), .B2(n_456), .Y(n_1132) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_128), .A2(n_311), .B1(n_726), .B2(n_837), .Y(n_878) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_129), .A2(n_208), .B1(n_859), .B2(n_860), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_130), .A2(n_239), .B1(n_603), .B2(n_778), .Y(n_777) );
XNOR2xp5_ASAP7_75t_L g1082 ( .A(n_131), .B(n_1083), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_132), .A2(n_148), .B1(n_433), .B2(n_516), .Y(n_1026) );
AOI22xp33_ASAP7_75t_SL g925 ( .A1(n_133), .A2(n_188), .B1(n_539), .B2(n_926), .Y(n_925) );
AOI22xp33_ASAP7_75t_SL g706 ( .A1(n_135), .A2(n_322), .B1(n_478), .B2(n_672), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g1118 ( .A(n_136), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_137), .A2(n_330), .B1(n_475), .B2(n_548), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_138), .A2(n_144), .B1(n_594), .B2(n_672), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_139), .A2(n_241), .B1(n_503), .B2(n_659), .Y(n_895) );
AOI22xp33_ASAP7_75t_SL g1103 ( .A1(n_140), .A2(n_246), .B1(n_662), .B2(n_663), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_141), .A2(n_367), .B1(n_669), .B2(n_786), .Y(n_785) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_142), .A2(n_342), .B1(n_433), .B2(n_581), .Y(n_580) );
AOI22xp33_ASAP7_75t_SL g1093 ( .A1(n_143), .A2(n_206), .B1(n_1044), .B2(n_1094), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_145), .A2(n_192), .B1(n_499), .B2(n_749), .Y(n_748) );
XNOR2x2_ASAP7_75t_L g734 ( .A(n_146), .B(n_735), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_147), .A2(n_160), .B1(n_488), .B2(n_671), .Y(n_1000) );
OA22x2_ASAP7_75t_L g685 ( .A1(n_149), .A2(n_686), .B1(n_687), .B2(n_707), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_149), .Y(n_686) );
INVx1_ASAP7_75t_L g903 ( .A(n_150), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_152), .B(n_587), .Y(n_944) );
AOI22xp33_ASAP7_75t_SL g1130 ( .A1(n_153), .A2(n_250), .B1(n_512), .B2(n_619), .Y(n_1130) );
AND2x6_ASAP7_75t_L g385 ( .A(n_154), .B(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g1073 ( .A(n_154), .Y(n_1073) );
AOI22xp33_ASAP7_75t_SL g1035 ( .A1(n_155), .A2(n_370), .B1(n_600), .B2(n_617), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1057 ( .A(n_156), .B(n_1058), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_157), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g857 ( .A(n_158), .B(n_498), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_159), .Y(n_805) );
AOI22xp33_ASAP7_75t_SL g1036 ( .A1(n_161), .A2(n_348), .B1(n_668), .B2(n_833), .Y(n_1036) );
AOI22xp5_ASAP7_75t_L g828 ( .A1(n_162), .A2(n_194), .B1(n_465), .B2(n_539), .Y(n_828) );
NAND2xp5_ASAP7_75t_SL g856 ( .A(n_163), .B(n_665), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_165), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_166), .A2(n_183), .B1(n_532), .B2(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_167), .B(n_893), .Y(n_920) );
AOI222xp33_ASAP7_75t_L g753 ( .A1(n_168), .A2(n_207), .B1(n_337), .B2(n_567), .C1(n_754), .C2(n_755), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_169), .A2(n_299), .B1(n_488), .B2(n_821), .Y(n_820) );
AOI22xp33_ASAP7_75t_SL g664 ( .A1(n_170), .A2(n_232), .B1(n_499), .B2(n_665), .Y(n_664) );
AO22x2_ASAP7_75t_L g413 ( .A1(n_171), .A2(n_247), .B1(n_404), .B2(n_408), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g1077 ( .A(n_171), .B(n_1078), .Y(n_1077) );
CKINVDCx20_ASAP7_75t_R g1097 ( .A(n_172), .Y(n_1097) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_173), .Y(n_682) );
AOI22xp33_ASAP7_75t_SL g947 ( .A1(n_174), .A2(n_289), .B1(n_452), .B2(n_463), .Y(n_947) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_175), .Y(n_554) );
AOI22xp33_ASAP7_75t_SL g667 ( .A1(n_176), .A2(n_268), .B1(n_668), .B2(n_669), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g977 ( .A(n_178), .Y(n_977) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_180), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g879 ( .A1(n_181), .A2(n_185), .B1(n_427), .B2(n_590), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_184), .A2(n_261), .B1(n_475), .B2(n_537), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_187), .A2(n_313), .B1(n_613), .B2(n_784), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_189), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_193), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g889 ( .A(n_195), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_198), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_200), .B(n_585), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_202), .A2(n_248), .B1(n_537), .B2(n_883), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_203), .A2(n_297), .B1(n_548), .B2(n_619), .Y(n_781) );
XNOR2xp5_ASAP7_75t_L g651 ( .A(n_209), .B(n_652), .Y(n_651) );
AOI22xp33_ASAP7_75t_SL g1032 ( .A1(n_211), .A2(n_238), .B1(n_510), .B2(n_928), .Y(n_1032) );
AOI22xp33_ASAP7_75t_SL g1033 ( .A1(n_212), .A2(n_231), .B1(n_478), .B2(n_620), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_214), .A2(n_333), .B1(n_680), .B2(n_998), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_215), .A2(n_340), .B1(n_619), .B2(n_621), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_216), .A2(n_236), .B1(n_617), .B2(n_672), .Y(n_834) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_218), .B(n_498), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g994 ( .A(n_219), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_220), .A2(n_321), .B1(n_490), .B2(n_539), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_221), .A2(n_353), .B1(n_427), .B2(n_433), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_222), .A2(n_265), .B1(n_472), .B2(n_716), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_225), .B(n_680), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_226), .A2(n_360), .B1(n_461), .B2(n_465), .Y(n_460) );
OA22x2_ASAP7_75t_L g1017 ( .A1(n_228), .A2(n_1018), .B1(n_1019), .B2(n_1020), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_228), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_233), .A2(n_252), .B1(n_492), .B2(n_494), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_234), .A2(n_324), .B1(n_490), .B2(n_738), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g1050 ( .A(n_235), .Y(n_1050) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_242), .Y(n_579) );
INVx2_ASAP7_75t_L g390 ( .A(n_244), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g715 ( .A1(n_245), .A2(n_293), .B1(n_494), .B2(n_716), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_253), .A2(n_282), .B1(n_591), .B2(n_751), .Y(n_1060) );
CKINVDCx14_ASAP7_75t_R g1110 ( .A(n_255), .Y(n_1110) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_255), .A2(n_1110), .B1(n_1114), .B2(n_1115), .Y(n_1113) );
CKINVDCx20_ASAP7_75t_R g1024 ( .A(n_256), .Y(n_1024) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_258), .Y(n_769) );
XNOR2x1_ASAP7_75t_L g912 ( .A(n_259), .B(n_913), .Y(n_912) );
AOI22xp5_ASAP7_75t_L g989 ( .A1(n_262), .A2(n_990), .B1(n_1014), .B2(n_1015), .Y(n_989) );
INVx1_ASAP7_75t_L g1014 ( .A(n_262), .Y(n_1014) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_263), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g1023 ( .A(n_264), .Y(n_1023) );
CKINVDCx20_ASAP7_75t_R g1010 ( .A(n_267), .Y(n_1010) );
CKINVDCx20_ASAP7_75t_R g1007 ( .A(n_270), .Y(n_1007) );
CKINVDCx20_ASAP7_75t_R g1119 ( .A(n_271), .Y(n_1119) );
CKINVDCx20_ASAP7_75t_R g986 ( .A(n_273), .Y(n_986) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_274), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g963 ( .A(n_275), .Y(n_963) );
AOI22x1_ASAP7_75t_L g760 ( .A1(n_276), .A2(n_761), .B1(n_789), .B2(n_790), .Y(n_760) );
INVx1_ASAP7_75t_L g789 ( .A(n_276), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_278), .Y(n_721) );
OA22x2_ASAP7_75t_L g955 ( .A1(n_280), .A2(n_956), .B1(n_957), .B2(n_958), .Y(n_955) );
CKINVDCx16_ASAP7_75t_R g956 ( .A(n_280), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_281), .B(n_498), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_284), .A2(n_350), .B1(n_478), .B2(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g404 ( .A(n_286), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_286), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_288), .A2(n_335), .B1(n_512), .B2(n_818), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_290), .B(n_692), .Y(n_1059) );
AOI22xp33_ASAP7_75t_SL g901 ( .A1(n_291), .A2(n_325), .B1(n_532), .B2(n_620), .Y(n_901) );
AOI22xp33_ASAP7_75t_SL g1087 ( .A1(n_292), .A2(n_368), .B1(n_451), .B2(n_673), .Y(n_1087) );
CKINVDCx20_ASAP7_75t_R g984 ( .A(n_296), .Y(n_984) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_300), .Y(n_798) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_301), .A2(n_383), .B(n_391), .C(n_1081), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_302), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g967 ( .A(n_303), .Y(n_967) );
CKINVDCx20_ASAP7_75t_R g970 ( .A(n_304), .Y(n_970) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_305), .A2(n_849), .B1(n_850), .B2(n_870), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_305), .Y(n_849) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_306), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g971 ( .A(n_307), .Y(n_971) );
CKINVDCx20_ASAP7_75t_R g1099 ( .A(n_308), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_309), .A2(n_358), .B1(n_506), .B2(n_590), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_310), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_312), .Y(n_733) );
INVx1_ASAP7_75t_L g389 ( .A(n_315), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_316), .Y(n_773) );
INVx1_ASAP7_75t_L g386 ( .A(n_318), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g965 ( .A(n_319), .Y(n_965) );
AOI22xp33_ASAP7_75t_SL g469 ( .A1(n_323), .A2(n_366), .B1(n_470), .B2(n_472), .Y(n_469) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_327), .A2(n_336), .B1(n_604), .B2(n_705), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_329), .Y(n_1013) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_331), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_334), .B(n_726), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_339), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_341), .A2(n_373), .B1(n_505), .B2(n_723), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_343), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_344), .B(n_893), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_346), .A2(n_380), .B1(n_726), .B2(n_837), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_347), .Y(n_414) );
AOI22xp33_ASAP7_75t_SL g1055 ( .A1(n_349), .A2(n_356), .B1(n_516), .B2(n_567), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_351), .A2(n_363), .B1(n_604), .B2(n_701), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_352), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_355), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g1030 ( .A(n_357), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_359), .B(n_587), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g1124 ( .A(n_361), .Y(n_1124) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_364), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_369), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_372), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_375), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_376), .B(n_585), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_378), .Y(n_810) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_385), .B(n_387), .Y(n_384) );
HB1xp67_ASAP7_75t_L g1072 ( .A(n_386), .Y(n_1072) );
OA21x2_ASAP7_75t_L g1108 ( .A1(n_387), .A2(n_1071), .B(n_1109), .Y(n_1108) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_646), .B1(n_1066), .B2(n_1067), .C(n_1068), .Y(n_391) );
INVx1_ASAP7_75t_L g1067 ( .A(n_392), .Y(n_1067) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_522), .B1(n_644), .B2(n_645), .Y(n_392) );
INVx1_ASAP7_75t_L g644 ( .A(n_393), .Y(n_644) );
AO22x1_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_484), .B1(n_520), .B2(n_521), .Y(n_393) );
INVx1_ASAP7_75t_L g520 ( .A(n_394), .Y(n_520) );
INVx2_ASAP7_75t_L g482 ( .A(n_395), .Y(n_482) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_448), .Y(n_395) );
NOR3xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_419), .C(n_436), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B1(n_414), .B2(n_415), .Y(n_397) );
INVx1_ASAP7_75t_L g962 ( .A(n_399), .Y(n_962) );
OAI221xp5_ASAP7_75t_SL g1003 ( .A1(n_399), .A2(n_1004), .B1(n_1005), .B2(n_1007), .C(n_1008), .Y(n_1003) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g553 ( .A(n_400), .Y(n_553) );
BUFx3_ASAP7_75t_L g625 ( .A(n_400), .Y(n_625) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_409), .Y(n_400) );
INVx2_ASAP7_75t_L g464 ( .A(n_401), .Y(n_464) );
OR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_407), .Y(n_401) );
AND2x2_ASAP7_75t_L g418 ( .A(n_402), .B(n_407), .Y(n_418) );
AND2x2_ASAP7_75t_L g455 ( .A(n_402), .B(n_431), .Y(n_455) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g422 ( .A(n_403), .B(n_407), .Y(n_422) );
AND2x2_ASAP7_75t_L g432 ( .A(n_403), .B(n_413), .Y(n_432) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_406), .Y(n_408) );
INVx2_ASAP7_75t_L g431 ( .A(n_407), .Y(n_431) );
INVx1_ASAP7_75t_L g481 ( .A(n_407), .Y(n_481) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2x1p5_ASAP7_75t_L g417 ( .A(n_410), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g473 ( .A(n_410), .B(n_455), .Y(n_473) );
AND2x4_ASAP7_75t_L g501 ( .A(n_410), .B(n_464), .Y(n_501) );
AND2x6_ASAP7_75t_L g587 ( .A(n_410), .B(n_418), .Y(n_587) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx1_ASAP7_75t_L g424 ( .A(n_411), .Y(n_424) );
INVx1_ASAP7_75t_L g430 ( .A(n_411), .Y(n_430) );
INVx1_ASAP7_75t_L g447 ( .A(n_411), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_411), .B(n_413), .Y(n_459) );
AND2x2_ASAP7_75t_L g423 ( .A(n_412), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g454 ( .A(n_413), .B(n_447), .Y(n_454) );
OA211x2_ASAP7_75t_L g495 ( .A1(n_415), .A2(n_496), .B(n_497), .C(n_502), .Y(n_495) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g627 ( .A(n_416), .Y(n_627) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx3_ASAP7_75t_L g555 ( .A(n_417), .Y(n_555) );
AND2x4_ASAP7_75t_L g467 ( .A(n_418), .B(n_423), .Y(n_467) );
AND2x2_ASAP7_75t_L g477 ( .A(n_418), .B(n_454), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_418), .B(n_454), .Y(n_678) );
OAI21xp5_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_425), .B(n_426), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_421), .Y(n_514) );
INVx2_ASAP7_75t_L g560 ( .A(n_421), .Y(n_560) );
INVx4_ASAP7_75t_L g578 ( .A(n_421), .Y(n_578) );
BUFx3_ASAP7_75t_L g754 ( .A(n_421), .Y(n_754) );
AND2x6_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g444 ( .A(n_422), .Y(n_444) );
AND2x4_ASAP7_75t_L g506 ( .A(n_422), .B(n_446), .Y(n_506) );
AND2x6_ASAP7_75t_L g463 ( .A(n_423), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g471 ( .A(n_423), .B(n_455), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_427), .Y(n_631) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_428), .Y(n_516) );
BUFx4f_ASAP7_75t_SL g558 ( .A(n_428), .Y(n_558) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_428), .Y(n_659) );
BUFx2_ASAP7_75t_L g755 ( .A(n_428), .Y(n_755) );
AND2x4_ASAP7_75t_L g428 ( .A(n_429), .B(n_432), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g435 ( .A(n_430), .Y(n_435) );
INVx1_ASAP7_75t_L g441 ( .A(n_431), .Y(n_441) );
AND2x4_ASAP7_75t_L g434 ( .A(n_432), .B(n_435), .Y(n_434) );
NAND2x1p5_ASAP7_75t_L g440 ( .A(n_432), .B(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g503 ( .A(n_432), .B(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g518 ( .A(n_433), .Y(n_518) );
BUFx4f_ASAP7_75t_SL g567 ( .A(n_433), .Y(n_567) );
BUFx12f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_434), .Y(n_635) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_434), .Y(n_723) );
INVx1_ASAP7_75t_L g1100 ( .A(n_434), .Y(n_1100) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_442), .B2(n_443), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_438), .A2(n_637), .B1(n_638), .B2(n_639), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_438), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_771) );
INVx3_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g562 ( .A(n_439), .Y(n_562) );
INVx4_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx3_ASAP7_75t_L g811 ( .A(n_440), .Y(n_811) );
OAI22xp33_ASAP7_75t_SL g969 ( .A1(n_440), .A2(n_639), .B1(n_970), .B2(n_971), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_440), .A2(n_443), .B1(n_1029), .B2(n_1030), .Y(n_1028) );
HB1xp67_ASAP7_75t_L g1125 ( .A(n_440), .Y(n_1125) );
AND2x2_ASAP7_75t_L g716 ( .A(n_441), .B(n_458), .Y(n_716) );
BUFx2_ASAP7_75t_L g569 ( .A(n_443), .Y(n_569) );
CKINVDCx16_ASAP7_75t_R g640 ( .A(n_443), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_443), .A2(n_1124), .B1(n_1125), .B2(n_1126), .Y(n_1123) );
OR2x6_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_468), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_460), .Y(n_449) );
BUFx4f_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g745 ( .A(n_452), .Y(n_745) );
BUFx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx3_ASAP7_75t_L g494 ( .A(n_453), .Y(n_494) );
BUFx3_ASAP7_75t_L g539 ( .A(n_453), .Y(n_539) );
BUFx3_ASAP7_75t_L g600 ( .A(n_453), .Y(n_600) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_454), .B(n_455), .Y(n_982) );
AND2x4_ASAP7_75t_L g457 ( .A(n_455), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g995 ( .A(n_456), .Y(n_995) );
BUFx2_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g490 ( .A(n_457), .Y(n_490) );
INVx1_ASAP7_75t_L g543 ( .A(n_457), .Y(n_543) );
BUFx2_ASAP7_75t_L g601 ( .A(n_457), .Y(n_601) );
BUFx3_ASAP7_75t_L g617 ( .A(n_457), .Y(n_617) );
BUFx3_ASAP7_75t_L g780 ( .A(n_457), .Y(n_780) );
BUFx2_ASAP7_75t_SL g926 ( .A(n_457), .Y(n_926) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x6_ASAP7_75t_L g480 ( .A(n_459), .B(n_481), .Y(n_480) );
INVx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_SL g603 ( .A(n_462), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_462), .B(n_682), .Y(n_681) );
INVx4_ASAP7_75t_L g833 ( .A(n_462), .Y(n_833) );
INVx11_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx11_ASAP7_75t_L g489 ( .A(n_463), .Y(n_489) );
INVx2_ASAP7_75t_L g978 ( .A(n_465), .Y(n_978) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g509 ( .A(n_466), .Y(n_509) );
INVx2_ASAP7_75t_L g604 ( .A(n_466), .Y(n_604) );
INVx2_ASAP7_75t_L g821 ( .A(n_466), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g1046 ( .A1(n_466), .A2(n_489), .B1(n_1047), .B2(n_1048), .Y(n_1046) );
INVx6_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx3_ASAP7_75t_L g532 ( .A(n_467), .Y(n_532) );
BUFx3_ASAP7_75t_L g668 ( .A(n_467), .Y(n_668) );
BUFx3_ASAP7_75t_L g788 ( .A(n_467), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_474), .Y(n_468) );
BUFx2_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g493 ( .A(n_471), .Y(n_493) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_471), .Y(n_537) );
BUFx2_ASAP7_75t_SL g594 ( .A(n_471), .Y(n_594) );
INVx4_ASAP7_75t_L g739 ( .A(n_472), .Y(n_739) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g510 ( .A(n_473), .Y(n_510) );
INVx2_ASAP7_75t_L g541 ( .A(n_473), .Y(n_541) );
BUFx3_ASAP7_75t_L g672 ( .A(n_473), .Y(n_672) );
BUFx3_ASAP7_75t_L g718 ( .A(n_473), .Y(n_718) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx3_ASAP7_75t_L g547 ( .A(n_476), .Y(n_547) );
INVx4_ASAP7_75t_L g597 ( .A(n_476), .Y(n_597) );
INVx5_ASAP7_75t_L g620 ( .A(n_476), .Y(n_620) );
INVx1_ASAP7_75t_L g705 ( .A(n_476), .Y(n_705) );
INVx2_ASAP7_75t_L g830 ( .A(n_476), .Y(n_830) );
INVx8_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g512 ( .A(n_479), .Y(n_512) );
BUFx4f_ASAP7_75t_SL g621 ( .A(n_479), .Y(n_621) );
INVx6_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g548 ( .A(n_480), .Y(n_548) );
INVx1_ASAP7_75t_SL g680 ( .A(n_480), .Y(n_680) );
INVx1_ASAP7_75t_SL g1094 ( .A(n_480), .Y(n_1094) );
INVx1_ASAP7_75t_L g504 ( .A(n_481), .Y(n_504) );
INVx1_ASAP7_75t_L g521 ( .A(n_484), .Y(n_521) );
XNOR2x2_ASAP7_75t_L g573 ( .A(n_484), .B(n_574), .Y(n_573) );
XOR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_519), .Y(n_484) );
NAND4xp75_ASAP7_75t_L g485 ( .A(n_486), .B(n_495), .C(n_507), .D(n_513), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_491), .Y(n_486) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_489), .Y(n_529) );
INVx4_ASAP7_75t_L g701 ( .A(n_489), .Y(n_701) );
INVx2_ASAP7_75t_SL g731 ( .A(n_489), .Y(n_731) );
INVx5_ASAP7_75t_SL g883 ( .A(n_489), .Y(n_883) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx3_ASAP7_75t_L g928 ( .A(n_493), .Y(n_928) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx5_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g692 ( .A(n_500), .Y(n_692) );
INVx2_ASAP7_75t_L g726 ( .A(n_500), .Y(n_726) );
INVx2_ASAP7_75t_L g893 ( .A(n_500), .Y(n_893) );
INVx4_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx3_ASAP7_75t_L g590 ( .A(n_503), .Y(n_590) );
BUFx2_ASAP7_75t_L g662 ( .A(n_503), .Y(n_662) );
BUFx2_ASAP7_75t_L g694 ( .A(n_503), .Y(n_694) );
INVx1_ASAP7_75t_L g752 ( .A(n_503), .Y(n_752) );
INVx1_ASAP7_75t_SL g861 ( .A(n_505), .Y(n_861) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_SL g591 ( .A(n_506), .Y(n_591) );
BUFx3_ASAP7_75t_L g663 ( .A(n_506), .Y(n_663) );
BUFx2_ASAP7_75t_SL g918 ( .A(n_506), .Y(n_918) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_511), .Y(n_507) );
INVx1_ASAP7_75t_L g985 ( .A(n_510), .Y(n_985) );
INVx2_ASAP7_75t_L g655 ( .A(n_514), .Y(n_655) );
INVx2_ASAP7_75t_SL g804 ( .A(n_514), .Y(n_804) );
BUFx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx4_ASAP7_75t_L g582 ( .A(n_516), .Y(n_582) );
INVx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g645 ( .A(n_522), .Y(n_645) );
OAI22xp5_ASAP7_75t_SL g522 ( .A1(n_523), .A2(n_524), .B1(n_607), .B2(n_643), .Y(n_522) );
INVx2_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_572), .B1(n_573), .B2(n_606), .Y(n_524) );
INVx2_ASAP7_75t_L g606 ( .A(n_525), .Y(n_606) );
INVx1_ASAP7_75t_L g570 ( .A(n_526), .Y(n_570) );
AND2x2_ASAP7_75t_SL g526 ( .A(n_527), .B(n_549), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_528), .B(n_540), .Y(n_527) );
OAI221xp5_ASAP7_75t_SL g528 ( .A1(n_529), .A2(n_530), .B1(n_531), .B2(n_533), .C(n_534), .Y(n_528) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_536), .A2(n_980), .B1(n_1050), .B2(n_1051), .Y(n_1049) );
INVx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx3_ASAP7_75t_L g613 ( .A(n_537), .Y(n_613) );
BUFx3_ASAP7_75t_L g743 ( .A(n_537), .Y(n_743) );
BUFx6f_ASAP7_75t_L g868 ( .A(n_537), .Y(n_868) );
BUFx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI221xp5_ASAP7_75t_SL g540 ( .A1(n_541), .A2(n_542), .B1(n_543), .B2(n_544), .C(n_545), .Y(n_540) );
INVx2_ASAP7_75t_L g616 ( .A(n_541), .Y(n_616) );
INVx1_ASAP7_75t_L g816 ( .A(n_541), .Y(n_816) );
INVx1_ASAP7_75t_L g673 ( .A(n_543), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g983 ( .A1(n_543), .A2(n_984), .B1(n_985), .B2(n_986), .Y(n_983) );
INVx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NOR3xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_556), .C(n_564), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_552), .B1(n_554), .B2(n_555), .Y(n_550) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g799 ( .A(n_553), .Y(n_799) );
BUFx3_ASAP7_75t_L g964 ( .A(n_555), .Y(n_964) );
INVx2_ASAP7_75t_L g1006 ( .A(n_555), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_555), .A2(n_625), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
OAI222xp33_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_559), .B1(n_560), .B2(n_561), .C1(n_562), .C2(n_563), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g1098 ( .A(n_558), .Y(n_1098) );
OAI221xp5_ASAP7_75t_L g763 ( .A1(n_560), .A2(n_631), .B1(n_764), .B2(n_765), .C(n_766), .Y(n_763) );
OAI21xp5_ASAP7_75t_L g888 ( .A1(n_560), .A2(n_889), .B(n_890), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .B1(n_568), .B2(n_569), .Y(n_564) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
XOR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_605), .Y(n_574) );
NAND3x1_ASAP7_75t_L g575 ( .A(n_576), .B(n_592), .C(n_598), .Y(n_575) );
NOR2x1_ASAP7_75t_L g576 ( .A(n_577), .B(n_583), .Y(n_576) );
OAI21xp5_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_579), .B(n_580), .Y(n_577) );
BUFx2_ASAP7_75t_L g629 ( .A(n_578), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g720 ( .A1(n_578), .A2(n_721), .B(n_722), .Y(n_720) );
OAI21xp5_ASAP7_75t_SL g915 ( .A1(n_578), .A2(n_916), .B(n_917), .Y(n_915) );
OAI21xp5_ASAP7_75t_L g939 ( .A1(n_578), .A2(n_940), .B(n_941), .Y(n_939) );
OAI21xp5_ASAP7_75t_SL g1053 ( .A1(n_578), .A2(n_1054), .B(n_1055), .Y(n_1053) );
INVx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_588), .C(n_589), .Y(n_583) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_SL g749 ( .A(n_586), .Y(n_749) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
BUFx2_ASAP7_75t_L g665 ( .A(n_587), .Y(n_665) );
BUFx4f_ASAP7_75t_L g837 ( .A(n_587), .Y(n_837) );
BUFx2_ASAP7_75t_L g1058 ( .A(n_587), .Y(n_1058) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
BUFx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx6f_ASAP7_75t_L g818 ( .A(n_597), .Y(n_818) );
INVx2_ASAP7_75t_L g1045 ( .A(n_597), .Y(n_1045) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .Y(n_598) );
BUFx2_ASAP7_75t_L g669 ( .A(n_600), .Y(n_669) );
INVx1_ASAP7_75t_L g643 ( .A(n_607), .Y(n_643) );
INVx1_ASAP7_75t_SL g642 ( .A(n_608), .Y(n_642) );
AND2x2_ASAP7_75t_SL g608 ( .A(n_609), .B(n_622), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_614), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_618), .Y(n_614) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_628), .C(n_636), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B1(n_626), .B2(n_627), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_625), .A2(n_627), .B1(n_769), .B2(n_770), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_627), .A2(n_798), .B1(n_799), .B2(n_800), .Y(n_797) );
OAI221xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_631), .B2(n_632), .C(n_633), .Y(n_628) );
OAI21xp5_ASAP7_75t_SL g695 ( .A1(n_629), .A2(n_696), .B(n_697), .Y(n_695) );
OAI21xp5_ASAP7_75t_SL g1120 ( .A1(n_629), .A2(n_1121), .B(n_1122), .Y(n_1120) );
OAI222xp33_ASAP7_75t_L g1009 ( .A1(n_631), .A2(n_804), .B1(n_1010), .B2(n_1011), .C1(n_1012), .C2(n_1013), .Y(n_1009) );
INVxp67_ASAP7_75t_L g1012 ( .A(n_634), .Y(n_1012) );
BUFx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx3_ASAP7_75t_L g807 ( .A(n_635), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_639), .A2(n_810), .B1(n_811), .B2(n_812), .Y(n_809) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g774 ( .A(n_640), .Y(n_774) );
INVx1_ASAP7_75t_L g1066 ( .A(n_646), .Y(n_1066) );
XOR2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_909), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B1(n_759), .B2(n_908), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_709), .B1(n_757), .B2(n_758), .Y(n_649) );
INVx1_ASAP7_75t_L g757 ( .A(n_650), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_683), .B1(n_684), .B2(n_708), .Y(n_650) );
INVx1_ASAP7_75t_L g708 ( .A(n_651), .Y(n_708) );
NAND3x1_ASAP7_75t_L g652 ( .A(n_653), .B(n_666), .C(n_674), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_660), .Y(n_653) );
OAI21xp5_ASAP7_75t_SL g654 ( .A1(n_655), .A2(n_656), .B(n_657), .Y(n_654) );
OAI21xp5_ASAP7_75t_SL g852 ( .A1(n_655), .A2(n_853), .B(n_854), .Y(n_852) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_664), .Y(n_660) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_670), .Y(n_666) );
BUFx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI21xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B(n_679), .Y(n_675) );
BUFx2_ASAP7_75t_R g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_SL g707 ( .A(n_687), .Y(n_707) );
NAND2x1p5_ASAP7_75t_L g687 ( .A(n_688), .B(n_698), .Y(n_687) );
NOR2xp67_ASAP7_75t_SL g688 ( .A(n_689), .B(n_695), .Y(n_688) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .C(n_693), .Y(n_689) );
NOR2x1_ASAP7_75t_L g698 ( .A(n_699), .B(n_703), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_706), .Y(n_703) );
INVx1_ASAP7_75t_L g758 ( .A(n_709), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B1(n_734), .B2(n_756), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
XOR2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_733), .Y(n_712) );
NAND3x1_ASAP7_75t_L g713 ( .A(n_714), .B(n_719), .C(n_729), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_717), .Y(n_714) );
BUFx2_ASAP7_75t_L g784 ( .A(n_718), .Y(n_784) );
NOR2x1_ASAP7_75t_L g719 ( .A(n_720), .B(n_724), .Y(n_719) );
BUFx4f_ASAP7_75t_L g767 ( .A(n_723), .Y(n_767) );
NAND3xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_727), .C(n_728), .Y(n_724) );
AND2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
INVx2_ASAP7_75t_L g756 ( .A(n_734), .Y(n_756) );
NAND4xp75_ASAP7_75t_L g735 ( .A(n_736), .B(n_741), .C(n_747), .D(n_753), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_740), .Y(n_736) );
INVx4_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx3_ASAP7_75t_L g864 ( .A(n_739), .Y(n_864) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_746), .Y(n_741) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_SL g747 ( .A(n_748), .B(n_750), .Y(n_747) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g859 ( .A(n_752), .Y(n_859) );
INVx3_ASAP7_75t_L g840 ( .A(n_754), .Y(n_840) );
INVx1_ASAP7_75t_L g802 ( .A(n_755), .Y(n_802) );
INVx1_ASAP7_75t_L g908 ( .A(n_759), .Y(n_908) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_791), .B1(n_906), .B2(n_907), .Y(n_759) );
INVx1_ASAP7_75t_L g906 ( .A(n_760), .Y(n_906) );
INVx2_ASAP7_75t_SL g790 ( .A(n_761), .Y(n_790) );
AND2x4_ASAP7_75t_L g761 ( .A(n_762), .B(n_775), .Y(n_761) );
NOR3xp33_ASAP7_75t_SL g762 ( .A(n_763), .B(n_768), .C(n_771), .Y(n_762) );
NOR2x1_ASAP7_75t_L g775 ( .A(n_776), .B(n_782), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_781), .Y(n_776) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_785), .Y(n_782) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g907 ( .A(n_791), .Y(n_907) );
XOR2xp5_ASAP7_75t_L g791 ( .A(n_792), .B(n_844), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B1(n_825), .B2(n_843), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_SL g824 ( .A(n_795), .Y(n_824) );
AND2x2_ASAP7_75t_L g795 ( .A(n_796), .B(n_813), .Y(n_795) );
NOR3xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_801), .C(n_809), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g1117 ( .A1(n_799), .A2(n_964), .B1(n_1118), .B2(n_1119), .Y(n_1117) );
OAI222xp33_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_803), .B1(n_804), .B2(n_805), .C1(n_806), .C2(n_808), .Y(n_801) );
OAI222xp33_ASAP7_75t_L g1096 ( .A1(n_804), .A2(n_1097), .B1(n_1098), .B2(n_1099), .C1(n_1100), .C2(n_1101), .Y(n_1096) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_819), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_817), .Y(n_814) );
NAND2xp5_ASAP7_75t_SL g819 ( .A(n_820), .B(n_822), .Y(n_819) );
INVx1_ASAP7_75t_SL g843 ( .A(n_825), .Y(n_843) );
NOR4xp75_ASAP7_75t_L g826 ( .A(n_827), .B(n_831), .C(n_835), .D(n_839), .Y(n_826) );
NAND2xp5_ASAP7_75t_SL g827 ( .A(n_828), .B(n_829), .Y(n_827) );
HB1xp67_ASAP7_75t_L g998 ( .A(n_830), .Y(n_998) );
NAND2xp5_ASAP7_75t_SL g831 ( .A(n_832), .B(n_834), .Y(n_831) );
NAND2xp5_ASAP7_75t_SL g835 ( .A(n_836), .B(n_838), .Y(n_835) );
OAI21xp5_ASAP7_75t_SL g839 ( .A1(n_840), .A2(n_841), .B(n_842), .Y(n_839) );
OAI21xp33_ASAP7_75t_SL g966 ( .A1(n_840), .A2(n_967), .B(n_968), .Y(n_966) );
AOI22xp5_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_846), .B1(n_871), .B2(n_872), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
BUFx2_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g870 ( .A(n_850), .Y(n_870) );
NAND3x1_ASAP7_75t_L g850 ( .A(n_851), .B(n_862), .C(n_866), .Y(n_850) );
NOR2x1_ASAP7_75t_L g851 ( .A(n_852), .B(n_855), .Y(n_851) );
NAND3xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_857), .C(n_858), .Y(n_855) );
INVx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
AND2x2_ASAP7_75t_L g862 ( .A(n_863), .B(n_865), .Y(n_862) );
AND2x2_ASAP7_75t_L g866 ( .A(n_867), .B(n_869), .Y(n_866) );
INVx1_ASAP7_75t_SL g871 ( .A(n_872), .Y(n_871) );
AO22x2_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_885), .B1(n_904), .B2(n_905), .Y(n_872) );
INVx1_ASAP7_75t_L g904 ( .A(n_873), .Y(n_904) );
NAND5xp2_ASAP7_75t_SL g874 ( .A(n_875), .B(n_876), .C(n_877), .D(n_880), .E(n_884), .Y(n_874) );
AND2x2_ASAP7_75t_SL g877 ( .A(n_878), .B(n_879), .Y(n_877) );
AND2x2_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
INVx1_ASAP7_75t_L g1090 ( .A(n_883), .Y(n_1090) );
INVx2_ASAP7_75t_L g905 ( .A(n_885), .Y(n_905) );
XOR2x2_ASAP7_75t_L g885 ( .A(n_886), .B(n_903), .Y(n_885) );
NAND2x1p5_ASAP7_75t_L g886 ( .A(n_887), .B(n_896), .Y(n_886) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_888), .B(n_891), .Y(n_887) );
NAND3xp33_ASAP7_75t_L g891 ( .A(n_892), .B(n_894), .C(n_895), .Y(n_891) );
NOR2x1_ASAP7_75t_L g896 ( .A(n_897), .B(n_900), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_901), .B(n_902), .Y(n_900) );
AOI22xp5_ASAP7_75t_L g909 ( .A1(n_910), .A2(n_911), .B1(n_951), .B2(n_1065), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
OAI22x1_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_932), .B1(n_933), .B2(n_950), .Y(n_911) );
INVx2_ASAP7_75t_L g950 ( .A(n_912), .Y(n_950) );
AND2x4_ASAP7_75t_L g913 ( .A(n_914), .B(n_923), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g914 ( .A(n_915), .B(n_919), .Y(n_914) );
NAND3xp33_ASAP7_75t_L g919 ( .A(n_920), .B(n_921), .C(n_922), .Y(n_919) );
NOR2x1_ASAP7_75t_L g923 ( .A(n_924), .B(n_929), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g924 ( .A(n_925), .B(n_927), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_930), .B(n_931), .Y(n_929) );
OA22x2_ASAP7_75t_L g1037 ( .A1(n_932), .A2(n_933), .B1(n_1038), .B2(n_1062), .Y(n_1037) );
INVx3_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
XOR2x2_ASAP7_75t_L g933 ( .A(n_934), .B(n_949), .Y(n_933) );
NAND3x1_ASAP7_75t_SL g934 ( .A(n_935), .B(n_938), .C(n_946), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_936), .B(n_937), .Y(n_935) );
NOR2x1_ASAP7_75t_L g938 ( .A(n_939), .B(n_942), .Y(n_938) );
NAND3xp33_ASAP7_75t_L g942 ( .A(n_943), .B(n_944), .C(n_945), .Y(n_942) );
AND2x2_ASAP7_75t_L g946 ( .A(n_947), .B(n_948), .Y(n_946) );
INVx1_ASAP7_75t_L g1065 ( .A(n_951), .Y(n_1065) );
XNOR2xp5_ASAP7_75t_SL g951 ( .A(n_952), .B(n_1016), .Y(n_951) );
AOI22xp5_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_954), .B1(n_987), .B2(n_988), .Y(n_952) );
INVx2_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
HB1xp67_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx2_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_959), .B(n_972), .Y(n_958) );
NOR3xp33_ASAP7_75t_L g959 ( .A(n_960), .B(n_966), .C(n_969), .Y(n_959) );
OAI22xp5_ASAP7_75t_SL g960 ( .A1(n_961), .A2(n_963), .B1(n_964), .B2(n_965), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
NOR3xp33_ASAP7_75t_L g972 ( .A(n_973), .B(n_976), .C(n_983), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_974), .B(n_975), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_977), .A2(n_978), .B1(n_979), .B2(n_980), .Y(n_976) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
INVx1_ASAP7_75t_L g993 ( .A(n_981), .Y(n_993) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx2_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g1015 ( .A(n_990), .Y(n_1015) );
AND2x2_ASAP7_75t_SL g990 ( .A(n_991), .B(n_1002), .Y(n_990) );
NOR2xp33_ASAP7_75t_L g991 ( .A(n_992), .B(n_999), .Y(n_991) );
OAI221xp5_ASAP7_75t_SL g992 ( .A1(n_993), .A2(n_994), .B1(n_995), .B2(n_996), .C(n_997), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1001), .Y(n_999) );
NOR2xp33_ASAP7_75t_SL g1002 ( .A(n_1003), .B(n_1009), .Y(n_1002) );
INVx2_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g1016 ( .A1(n_1017), .A2(n_1037), .B1(n_1063), .B2(n_1064), .Y(n_1016) );
INVx2_ASAP7_75t_SL g1063 ( .A(n_1017), .Y(n_1063) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
AND3x1_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1031), .C(n_1034), .Y(n_1020) );
NOR3xp33_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1025), .C(n_1028), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1027), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1033), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .Y(n_1034) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1037), .Y(n_1064) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1038), .Y(n_1062) );
XOR2x2_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1061), .Y(n_1038) );
AND2x2_ASAP7_75t_SL g1039 ( .A(n_1040), .B(n_1052), .Y(n_1039) );
NOR3xp33_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1046), .C(n_1049), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1043), .Y(n_1041) );
INVx3_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
NOR2xp33_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1056), .Y(n_1052) );
NAND3xp33_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1059), .C(n_1060), .Y(n_1056) );
INVx1_ASAP7_75t_SL g1068 ( .A(n_1069), .Y(n_1068) );
NOR2x1_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1074), .Y(n_1069) );
OR2x2_ASAP7_75t_SL g1134 ( .A(n_1070), .B(n_1075), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1073), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
OAI322xp33_ASAP7_75t_L g1081 ( .A1(n_1072), .A2(n_1082), .A3(n_1105), .B1(n_1108), .B2(n_1110), .C1(n_1111), .C2(n_1134), .Y(n_1081) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1072), .B(n_1107), .Y(n_1109) );
CKINVDCx16_ASAP7_75t_R g1107 ( .A(n_1073), .Y(n_1107) );
CKINVDCx20_ASAP7_75t_R g1074 ( .A(n_1075), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1077), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1080), .Y(n_1078) );
HB1xp67_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
NAND2xp5_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1095), .Y(n_1084) );
NOR2xp33_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1091), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1087), .B(n_1088), .Y(n_1086) );
INVx2_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1093), .Y(n_1091) );
NOR2xp33_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1102), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1104), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
HB1xp67_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1127), .Y(n_1115) );
NOR3xp33_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1120), .C(n_1123), .Y(n_1116) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1131), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1129), .B(n_1130), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1133), .Y(n_1131) );
endmodule