module fake_netlist_5_568_n_1689 (n_137, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1689);

input n_137;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1689;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_60),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_78),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_59),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_115),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_28),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_28),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_125),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_52),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_146),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_50),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_63),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_20),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_69),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_119),
.Y(n_183)
);

BUFx8_ASAP7_75t_SL g184 ( 
.A(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_0),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_91),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_51),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_29),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_19),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_57),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_38),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_45),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_150),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_98),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_32),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_27),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_132),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_74),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_106),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_39),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_23),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_56),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_67),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_62),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_54),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_72),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_38),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_37),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_109),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_22),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_134),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_58),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_158),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_127),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_14),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_116),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_143),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_110),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_103),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_133),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_21),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_104),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_111),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_122),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_59),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_7),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_142),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_50),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_88),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_13),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_105),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_11),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_40),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_97),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_161),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_33),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_32),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_9),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_64),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_45),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_165),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_53),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_95),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_14),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_89),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_5),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_0),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_10),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_65),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_41),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_6),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_15),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_144),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_13),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_1),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_163),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_6),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_34),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_81),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_3),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_18),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_85),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_20),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_57),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_118),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_131),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_66),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_49),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_124),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_159),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_33),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_153),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_77),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_112),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_2),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_126),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_92),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_79),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_47),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_41),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_53),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_51),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_164),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_80),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_99),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_148),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_52),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_25),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_46),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_73),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_36),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_36),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_43),
.Y(n_298)
);

BUFx2_ASAP7_75t_SL g299 ( 
.A(n_34),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_19),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_100),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_68),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_93),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_8),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_2),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_58),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_30),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_84),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_1),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_87),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_47),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_15),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_156),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_120),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_46),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_8),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_147),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_24),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_154),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_83),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_160),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_141),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_3),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_61),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_35),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_136),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_71),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_48),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_35),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_137),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_40),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_172),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_194),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_275),
.B(n_4),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_184),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_194),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_183),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_210),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_233),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_275),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_210),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_233),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_168),
.B(n_4),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_167),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_252),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_172),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_170),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_174),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_252),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_322),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_219),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_213),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_176),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_285),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_322),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_213),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_227),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_285),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_178),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_197),
.B(n_5),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_297),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_258),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_297),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_279),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_197),
.B(n_7),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_180),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_309),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_182),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_186),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_168),
.B(n_9),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_237),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_302),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_280),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_195),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_171),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_237),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_305),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_324),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_299),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_189),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_299),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_201),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_305),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_203),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_237),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_211),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_214),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_216),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_218),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_318),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_222),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_318),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_173),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_173),
.Y(n_397)
);

NOR2xp67_ASAP7_75t_L g398 ( 
.A(n_181),
.B(n_10),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_177),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_R g400 ( 
.A(n_223),
.B(n_166),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_225),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_175),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_228),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_232),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_221),
.B(n_11),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_177),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_185),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_236),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_185),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_187),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_192),
.B(n_12),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_239),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_187),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_334),
.B(n_196),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_345),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_345),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_378),
.B(n_192),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_344),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_370),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_370),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_381),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_347),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_333),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_402),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_402),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_333),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_336),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_348),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_337),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_396),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_397),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_353),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_336),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_359),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_R g436 ( 
.A(n_335),
.B(n_383),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_368),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_332),
.B(n_169),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_398),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_378),
.B(n_221),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_384),
.B(n_200),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_384),
.B(n_224),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_397),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_385),
.B(n_200),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_369),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_399),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_375),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_332),
.A2(n_306),
.B1(n_329),
.B2(n_198),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_398),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_340),
.B(n_246),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_351),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_339),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_399),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_385),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_339),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_392),
.B(n_224),
.Y(n_456)
);

INVx6_ASAP7_75t_L g457 ( 
.A(n_372),
.Y(n_457)
);

OAI21x1_ASAP7_75t_L g458 ( 
.A1(n_360),
.A2(n_330),
.B(n_254),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_342),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_342),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_366),
.B(n_261),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_349),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_388),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_389),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_406),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_390),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_L g467 ( 
.A(n_380),
.B(n_254),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_357),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_406),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_362),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_392),
.B(n_204),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_349),
.Y(n_472)
);

OA21x2_ASAP7_75t_L g473 ( 
.A1(n_365),
.A2(n_208),
.B(n_204),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_391),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_407),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_393),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_346),
.B(n_169),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_401),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_404),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_354),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_394),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_R g482 ( 
.A(n_386),
.B(n_240),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_412),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_354),
.Y(n_484)
);

CKINVDCx11_ASAP7_75t_R g485 ( 
.A(n_364),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_376),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_407),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_394),
.Y(n_488)
);

OR2x6_ASAP7_75t_L g489 ( 
.A(n_457),
.B(n_181),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_454),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_428),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_414),
.B(n_346),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_440),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_417),
.B(n_395),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_461),
.B(n_395),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_415),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_454),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_414),
.B(n_450),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_454),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_417),
.B(n_382),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_473),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_428),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_417),
.B(n_358),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_450),
.B(n_244),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_423),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_415),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_481),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_481),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_451),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_423),
.Y(n_510)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_428),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_448),
.B(n_373),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_441),
.B(n_208),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_421),
.Y(n_514)
);

NAND3xp33_ASAP7_75t_L g515 ( 
.A(n_439),
.B(n_449),
.C(n_356),
.Y(n_515)
);

OR2x6_ASAP7_75t_L g516 ( 
.A(n_457),
.B(n_405),
.Y(n_516)
);

AND2x6_ASAP7_75t_L g517 ( 
.A(n_441),
.B(n_188),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_473),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_L g519 ( 
.A(n_439),
.B(n_188),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_431),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_473),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_415),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_431),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_432),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_482),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_449),
.B(n_264),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_428),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_432),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_421),
.B(n_350),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_473),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_441),
.B(n_267),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_440),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_443),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_418),
.B(n_350),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_428),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_428),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_426),
.B(n_355),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_446),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_440),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_428),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_455),
.Y(n_542)
);

AND2x2_ASAP7_75t_SL g543 ( 
.A(n_473),
.B(n_355),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_446),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_440),
.Y(n_545)
);

OR2x2_ASAP7_75t_SL g546 ( 
.A(n_486),
.B(n_372),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_422),
.B(n_403),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_444),
.B(n_270),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_455),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_426),
.B(n_377),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_429),
.B(n_408),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_455),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_433),
.B(n_377),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_444),
.B(n_358),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_425),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_486),
.Y(n_556)
);

BUFx8_ASAP7_75t_SL g557 ( 
.A(n_468),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_453),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_453),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_442),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_444),
.B(n_361),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_455),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_471),
.B(n_272),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_465),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_442),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_471),
.B(n_277),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_471),
.B(n_278),
.Y(n_567)
);

AND2x2_ASAP7_75t_SL g568 ( 
.A(n_442),
.B(n_343),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_425),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_455),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_442),
.B(n_456),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_435),
.B(n_387),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_437),
.B(n_387),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_465),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_456),
.B(n_361),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_445),
.B(n_338),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_455),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_459),
.B(n_188),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_485),
.Y(n_579)
);

NOR2x1p5_ASAP7_75t_L g580 ( 
.A(n_447),
.B(n_179),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_469),
.Y(n_581)
);

AND2x2_ASAP7_75t_SL g582 ( 
.A(n_456),
.B(n_371),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_456),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_467),
.B(n_281),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_463),
.B(n_400),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_464),
.B(n_169),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_459),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_469),
.B(n_209),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_466),
.B(n_341),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_474),
.B(n_169),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_459),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_459),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_476),
.B(n_288),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_457),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_459),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_459),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_436),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_467),
.B(n_282),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_475),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_462),
.Y(n_600)
);

BUFx4f_ASAP7_75t_L g601 ( 
.A(n_462),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_478),
.B(n_288),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_475),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_438),
.B(n_352),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_487),
.B(n_209),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_462),
.Y(n_606)
);

OAI22xp33_ASAP7_75t_SL g607 ( 
.A1(n_477),
.A2(n_411),
.B1(n_250),
.B2(n_274),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_462),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_462),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_462),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_462),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_458),
.A2(n_374),
.B1(n_199),
.B2(n_212),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_480),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_479),
.B(n_191),
.C(n_190),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_483),
.B(n_379),
.Y(n_615)
);

BUFx10_ASAP7_75t_L g616 ( 
.A(n_457),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_487),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_458),
.A2(n_212),
.B1(n_215),
.B2(n_199),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_416),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_416),
.Y(n_620)
);

NAND2xp33_ASAP7_75t_L g621 ( 
.A(n_480),
.B(n_188),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_419),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_457),
.B(n_193),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_424),
.B(n_434),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_448),
.B(n_230),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_419),
.B(n_363),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_420),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_420),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_480),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_424),
.B(n_205),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_424),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_424),
.B(n_283),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_480),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_430),
.B(n_288),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_434),
.Y(n_635)
);

AND2x6_ASAP7_75t_L g636 ( 
.A(n_434),
.B(n_188),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_SL g637 ( 
.A(n_498),
.B(n_238),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_490),
.B(n_434),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_494),
.B(n_472),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_492),
.B(n_430),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_490),
.B(n_472),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_514),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_507),
.B(n_472),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_525),
.B(n_597),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_504),
.B(n_470),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_494),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_497),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_508),
.B(n_472),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_543),
.A2(n_289),
.B1(n_290),
.B2(n_295),
.Y(n_649)
);

OR2x2_ASAP7_75t_SL g650 ( 
.A(n_625),
.B(n_215),
.Y(n_650)
);

INVxp67_ASAP7_75t_SL g651 ( 
.A(n_493),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_500),
.B(n_484),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_496),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_545),
.A2(n_458),
.B(n_452),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_571),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_497),
.B(n_229),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_630),
.B(n_484),
.Y(n_657)
);

OR2x6_ASAP7_75t_L g658 ( 
.A(n_594),
.B(n_229),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_496),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_499),
.B(n_484),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_543),
.A2(n_330),
.B1(n_308),
.B2(n_234),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_500),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_545),
.A2(n_583),
.B(n_560),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_571),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_506),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_506),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_576),
.B(n_257),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_568),
.B(n_484),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_503),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_501),
.A2(n_274),
.B1(n_303),
.B2(n_234),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_503),
.B(n_427),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_607),
.B(n_488),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_526),
.B(n_266),
.Y(n_673)
);

BUFx6f_ASAP7_75t_SL g674 ( 
.A(n_568),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_582),
.B(n_480),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_522),
.Y(n_676)
);

OAI22xp33_ASAP7_75t_L g677 ( 
.A1(n_604),
.A2(n_248),
.B1(n_271),
.B2(n_291),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_582),
.B(n_480),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_495),
.B(n_301),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_525),
.B(n_310),
.Y(n_680)
);

NOR3xp33_ASAP7_75t_L g681 ( 
.A(n_550),
.B(n_312),
.C(n_259),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_516),
.A2(n_326),
.B1(n_313),
.B2(n_314),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_623),
.B(n_317),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_505),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_516),
.A2(n_319),
.B1(n_321),
.B2(n_248),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_522),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_L g687 ( 
.A(n_618),
.B(n_188),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_505),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_501),
.A2(n_303),
.B1(n_250),
.B2(n_271),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_SL g690 ( 
.A1(n_512),
.A2(n_253),
.B1(n_256),
.B2(n_251),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_501),
.A2(n_321),
.B1(n_319),
.B2(n_308),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_627),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_510),
.B(n_480),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_627),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_616),
.B(n_320),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_628),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_510),
.B(n_291),
.Y(n_697)
);

OR2x6_ASAP7_75t_L g698 ( 
.A(n_594),
.B(n_231),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_628),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_631),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_589),
.B(n_206),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_520),
.B(n_427),
.Y(n_702)
);

O2A1O1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_519),
.A2(n_231),
.B(n_243),
.C(n_287),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_523),
.B(n_452),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_631),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_523),
.B(n_452),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_524),
.B(n_460),
.Y(n_707)
);

AND2x6_ASAP7_75t_SL g708 ( 
.A(n_535),
.B(n_243),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_616),
.B(n_327),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_524),
.B(n_460),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_528),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_554),
.Y(n_712)
);

NOR3xp33_ASAP7_75t_L g713 ( 
.A(n_529),
.B(n_207),
.C(n_217),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_518),
.A2(n_202),
.B1(n_287),
.B2(n_286),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_635),
.Y(n_715)
);

NOR2x1p5_ASAP7_75t_L g716 ( 
.A(n_604),
.B(n_255),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_616),
.B(n_545),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_528),
.B(n_460),
.Y(n_718)
);

INVx4_ASAP7_75t_L g719 ( 
.A(n_493),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_531),
.B(n_202),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_555),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_531),
.B(n_202),
.Y(n_722)
);

INVxp33_ASAP7_75t_L g723 ( 
.A(n_556),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_534),
.B(n_202),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_560),
.A2(n_202),
.B(n_363),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_534),
.B(n_544),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_544),
.B(n_202),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_554),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_558),
.B(n_409),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_558),
.B(n_409),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_560),
.B(n_288),
.Y(n_731)
);

O2A1O1Ixp5_ASAP7_75t_L g732 ( 
.A1(n_518),
.A2(n_413),
.B(n_410),
.C(n_367),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_559),
.B(n_410),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_559),
.B(n_413),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_513),
.A2(n_311),
.B1(n_220),
.B2(n_273),
.Y(n_735)
);

BUFx6f_ASAP7_75t_SL g736 ( 
.A(n_489),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_583),
.B(n_226),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_635),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_564),
.Y(n_739)
);

XOR2xp5_ASAP7_75t_L g740 ( 
.A(n_512),
.B(n_235),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_583),
.A2(n_367),
.B(n_331),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_493),
.B(n_241),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_493),
.B(n_242),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_564),
.B(n_245),
.Y(n_744)
);

O2A1O1Ixp5_ASAP7_75t_L g745 ( 
.A1(n_518),
.A2(n_292),
.B(n_328),
.C(n_325),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_581),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_581),
.B(n_247),
.Y(n_747)
);

NAND2x1p5_ASAP7_75t_L g748 ( 
.A(n_530),
.B(n_255),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_521),
.A2(n_331),
.B1(n_328),
.B2(n_325),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_599),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_599),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_533),
.B(n_249),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_603),
.B(n_617),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_603),
.B(n_262),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_617),
.B(n_263),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_561),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_539),
.B(n_574),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_532),
.B(n_265),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_561),
.B(n_260),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_575),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_575),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_548),
.B(n_268),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_533),
.B(n_323),
.Y(n_763)
);

A2O1A1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_530),
.A2(n_513),
.B(n_612),
.C(n_566),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_563),
.B(n_316),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_619),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_513),
.B(n_315),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_533),
.B(n_293),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_540),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_567),
.B(n_294),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_540),
.B(n_565),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_521),
.A2(n_315),
.B1(n_307),
.B2(n_260),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_540),
.B(n_296),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_521),
.A2(n_307),
.B1(n_286),
.B2(n_292),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_540),
.B(n_304),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_565),
.B(n_632),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_565),
.A2(n_269),
.B1(n_237),
.B2(n_284),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_515),
.B(n_300),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_585),
.B(n_298),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_565),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_620),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_565),
.B(n_584),
.Y(n_782)
);

O2A1O1Ixp5_ASAP7_75t_L g783 ( 
.A1(n_624),
.A2(n_269),
.B(n_276),
.C(n_70),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_614),
.B(n_269),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_622),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_L g786 ( 
.A1(n_516),
.A2(n_269),
.B1(n_16),
.B2(n_17),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_588),
.A2(n_12),
.B1(n_16),
.B2(n_17),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_588),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_592),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_634),
.B(n_23),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_588),
.B(n_82),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_598),
.B(n_76),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_626),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_626),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_527),
.Y(n_795)
);

NOR2x1p5_ASAP7_75t_L g796 ( 
.A(n_597),
.B(n_24),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_605),
.B(n_86),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_605),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_555),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_605),
.B(n_90),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_553),
.B(n_25),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_516),
.B(n_94),
.Y(n_802)
);

OAI221xp5_ASAP7_75t_L g803 ( 
.A1(n_625),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.C(n_30),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_572),
.B(n_26),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_764),
.A2(n_489),
.B1(n_569),
.B2(n_547),
.Y(n_805)
);

OAI21x1_ASAP7_75t_SL g806 ( 
.A1(n_797),
.A2(n_542),
.B(n_633),
.Y(n_806)
);

O2A1O1Ixp5_ASAP7_75t_L g807 ( 
.A1(n_672),
.A2(n_601),
.B(n_590),
.C(n_593),
.Y(n_807)
);

AND2x2_ASAP7_75t_SL g808 ( 
.A(n_687),
.B(n_519),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_652),
.B(n_489),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_771),
.A2(n_601),
.B(n_591),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_782),
.A2(n_601),
.B(n_591),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_652),
.B(n_489),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_799),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_776),
.A2(n_591),
.B(n_592),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_667),
.B(n_538),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_799),
.B(n_569),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_655),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_669),
.B(n_586),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_662),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_669),
.B(n_712),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_647),
.B(n_580),
.Y(n_821)
);

O2A1O1Ixp5_ASAP7_75t_L g822 ( 
.A1(n_745),
.A2(n_602),
.B(n_629),
.C(n_549),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_640),
.B(n_551),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_769),
.A2(n_663),
.B(n_651),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_662),
.B(n_615),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_668),
.B(n_549),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_700),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_721),
.Y(n_828)
);

O2A1O1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_661),
.A2(n_573),
.B(n_578),
.C(n_621),
.Y(n_829)
);

NAND2x1p5_ASAP7_75t_L g830 ( 
.A(n_719),
.B(n_491),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_673),
.A2(n_552),
.B(n_562),
.C(n_613),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_701),
.B(n_546),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_664),
.Y(n_833)
);

A2O1A1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_798),
.A2(n_664),
.B(n_790),
.C(n_784),
.Y(n_834)
);

NAND2x1p5_ASAP7_75t_L g835 ( 
.A(n_719),
.B(n_595),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_712),
.B(n_579),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_719),
.A2(n_587),
.B(n_600),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_728),
.B(n_595),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_642),
.B(n_546),
.Y(n_839)
);

AO21x1_ASAP7_75t_L g840 ( 
.A1(n_637),
.A2(n_621),
.B(n_578),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_717),
.A2(n_657),
.B(n_789),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_645),
.B(n_491),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_798),
.A2(n_606),
.B(n_613),
.C(n_611),
.Y(n_843)
);

O2A1O1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_748),
.A2(n_600),
.B(n_611),
.C(n_610),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_700),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_647),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_791),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_728),
.B(n_570),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_646),
.A2(n_606),
.B(n_610),
.C(n_609),
.Y(n_849)
);

A2O1A1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_646),
.A2(n_608),
.B(n_609),
.C(n_491),
.Y(n_850)
);

O2A1O1Ixp5_ASAP7_75t_L g851 ( 
.A1(n_783),
.A2(n_608),
.B(n_502),
.C(n_596),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_756),
.B(n_793),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_670),
.A2(n_502),
.B1(n_596),
.B2(n_595),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_756),
.B(n_502),
.Y(n_854)
);

O2A1O1Ixp33_ASAP7_75t_SL g855 ( 
.A1(n_800),
.A2(n_570),
.B(n_536),
.C(n_517),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_793),
.B(n_794),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_794),
.B(n_570),
.Y(n_857)
);

A2O1A1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_778),
.A2(n_536),
.B(n_579),
.C(n_509),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_637),
.A2(n_517),
.B1(n_636),
.B2(n_509),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_789),
.A2(n_577),
.B(n_541),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_760),
.B(n_129),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_705),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_723),
.B(n_557),
.Y(n_863)
);

NOR2x1p5_ASAP7_75t_SL g864 ( 
.A(n_795),
.B(n_517),
.Y(n_864)
);

CKINVDCx6p67_ASAP7_75t_R g865 ( 
.A(n_736),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_687),
.A2(n_577),
.B(n_541),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_643),
.A2(n_577),
.B(n_541),
.Y(n_867)
);

A2O1A1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_760),
.A2(n_517),
.B(n_577),
.C(n_541),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_748),
.A2(n_517),
.B(n_636),
.Y(n_869)
);

AND2x2_ASAP7_75t_SL g870 ( 
.A(n_802),
.B(n_791),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_644),
.B(n_541),
.Y(n_871)
);

AO21x1_ASAP7_75t_L g872 ( 
.A1(n_685),
.A2(n_31),
.B(n_37),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_702),
.A2(n_537),
.B(n_511),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_715),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_723),
.B(n_557),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_671),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_648),
.A2(n_537),
.B(n_511),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_639),
.B(n_636),
.Y(n_878)
);

AOI21x1_ASAP7_75t_L g879 ( 
.A1(n_704),
.A2(n_537),
.B(n_511),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_639),
.B(n_636),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_791),
.B(n_780),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_726),
.A2(n_636),
.B(n_113),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_753),
.A2(n_636),
.B(n_107),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_758),
.B(n_31),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_684),
.B(n_39),
.Y(n_885)
);

OAI22x1_ASAP7_75t_L g886 ( 
.A1(n_740),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_761),
.A2(n_779),
.B(n_684),
.C(n_746),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_762),
.B(n_42),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_765),
.B(n_128),
.Y(n_889)
);

O2A1O1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_748),
.A2(n_44),
.B(n_48),
.C(n_49),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_759),
.Y(n_891)
);

AOI21x1_ASAP7_75t_L g892 ( 
.A1(n_706),
.A2(n_138),
.B(n_155),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_638),
.A2(n_135),
.B(n_152),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_761),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_641),
.A2(n_114),
.B(n_151),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_759),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_688),
.A2(n_750),
.B(n_711),
.C(n_746),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_688),
.A2(n_54),
.B(n_55),
.C(n_56),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_660),
.A2(n_75),
.B(n_96),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_711),
.B(n_55),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_698),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_738),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_750),
.B(n_139),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_671),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_773),
.A2(n_140),
.B(n_149),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_689),
.A2(n_162),
.B1(n_691),
.B2(n_714),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_716),
.B(n_735),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_770),
.B(n_649),
.Y(n_908)
);

AOI33xp33_ASAP7_75t_L g909 ( 
.A1(n_677),
.A2(n_735),
.A3(n_777),
.B1(n_787),
.B2(n_788),
.B3(n_749),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_738),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_739),
.A2(n_751),
.B(n_767),
.C(n_766),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_692),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_681),
.B(n_804),
.C(n_801),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_803),
.A2(n_786),
.B(n_697),
.C(n_744),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_SL g915 ( 
.A1(n_792),
.A2(n_731),
.B(n_720),
.C(n_722),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_739),
.B(n_751),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_716),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_650),
.B(n_757),
.Y(n_918)
);

NAND3xp33_ASAP7_75t_L g919 ( 
.A(n_713),
.B(n_679),
.C(n_747),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_754),
.A2(n_755),
.B(n_730),
.C(n_733),
.Y(n_920)
);

NOR2x1_ASAP7_75t_L g921 ( 
.A(n_680),
.B(n_709),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_767),
.B(n_656),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_775),
.A2(n_693),
.B(n_710),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_650),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_692),
.B(n_696),
.Y(n_925)
);

A2O1A1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_766),
.A2(n_781),
.B(n_785),
.C(n_696),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_674),
.A2(n_774),
.B1(n_772),
.B2(n_682),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_656),
.B(n_740),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_694),
.B(n_699),
.Y(n_929)
);

NOR2xp67_ASAP7_75t_L g930 ( 
.A(n_781),
.B(n_785),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_656),
.B(n_690),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_653),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_729),
.B(n_734),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_674),
.B(n_698),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_674),
.B(n_698),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_698),
.B(n_658),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_737),
.A2(n_763),
.B1(n_743),
.B2(n_742),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_752),
.B(n_768),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_703),
.A2(n_718),
.B(n_707),
.C(n_741),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_659),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_658),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_665),
.B(n_666),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_683),
.A2(n_658),
.B1(n_736),
.B2(n_695),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_L g944 ( 
.A(n_787),
.B(n_788),
.C(n_658),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_676),
.A2(n_686),
.B(n_724),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_676),
.A2(n_686),
.B(n_727),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_736),
.A2(n_796),
.B1(n_725),
.B2(n_708),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_796),
.B(n_498),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_655),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_662),
.B(n_514),
.Y(n_950)
);

BUFx4f_ASAP7_75t_L g951 ( 
.A(n_799),
.Y(n_951)
);

AO21x2_ASAP7_75t_L g952 ( 
.A1(n_675),
.A2(n_678),
.B(n_764),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_652),
.B(n_498),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_655),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_764),
.A2(n_668),
.B1(n_678),
.B2(n_675),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_764),
.A2(n_668),
.B1(n_678),
.B2(n_675),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_652),
.B(n_498),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_764),
.A2(n_732),
.B(n_668),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_771),
.A2(n_782),
.B(n_776),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_771),
.A2(n_782),
.B(n_776),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_662),
.A2(n_498),
.B1(n_637),
.B2(n_655),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_771),
.A2(n_782),
.B(n_776),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_764),
.A2(n_732),
.B(n_668),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_764),
.A2(n_732),
.B(n_668),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_662),
.A2(n_498),
.B1(n_637),
.B2(n_655),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_764),
.A2(n_668),
.B1(n_678),
.B2(n_675),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_654),
.A2(n_663),
.B(n_641),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_L g968 ( 
.A(n_667),
.B(n_498),
.C(n_640),
.Y(n_968)
);

NAND2x1p5_ASAP7_75t_L g969 ( 
.A(n_719),
.B(n_791),
.Y(n_969)
);

INVxp67_ASAP7_75t_L g970 ( 
.A(n_662),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_652),
.B(n_498),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_652),
.B(n_498),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_799),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_661),
.A2(n_498),
.B(n_662),
.C(n_672),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_968),
.B(n_953),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_823),
.B(n_891),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_958),
.A2(n_964),
.B(n_963),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_974),
.A2(n_971),
.B(n_957),
.Y(n_978)
);

NOR2xp67_ASAP7_75t_L g979 ( 
.A(n_913),
.B(n_919),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_968),
.B(n_972),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_823),
.B(n_904),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_847),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_813),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_847),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_904),
.B(n_896),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_876),
.B(n_815),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_815),
.B(n_918),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_918),
.B(n_924),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_894),
.B(n_933),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_959),
.A2(n_962),
.B(n_960),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_909),
.A2(n_884),
.B(n_888),
.C(n_944),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_847),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_814),
.A2(n_806),
.B(n_810),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_884),
.A2(n_888),
.B(n_832),
.C(n_914),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_816),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_834),
.A2(n_887),
.B(n_897),
.C(n_948),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_847),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_827),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_894),
.B(n_852),
.Y(n_999)
);

AO31x2_ASAP7_75t_L g1000 ( 
.A1(n_955),
.A2(n_966),
.A3(n_956),
.B(n_840),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_923),
.A2(n_881),
.B(n_824),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_881),
.A2(n_841),
.B(n_811),
.Y(n_1002)
);

AOI21xp33_ASAP7_75t_L g1003 ( 
.A1(n_832),
.A2(n_927),
.B(n_908),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_SL g1004 ( 
.A1(n_872),
.A2(n_890),
.B(n_903),
.Y(n_1004)
);

NAND3xp33_ASAP7_75t_SL g1005 ( 
.A(n_961),
.B(n_965),
.C(n_807),
.Y(n_1005)
);

INVxp67_ASAP7_75t_SL g1006 ( 
.A(n_969),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_951),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_870),
.A2(n_969),
.B1(n_809),
.B2(n_812),
.Y(n_1008)
);

INVx5_ASAP7_75t_L g1009 ( 
.A(n_901),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_870),
.A2(n_856),
.B1(n_808),
.B2(n_930),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_911),
.A2(n_880),
.B(n_878),
.Y(n_1011)
);

INVx5_ASAP7_75t_L g1012 ( 
.A(n_901),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_845),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_922),
.B(n_817),
.Y(n_1014)
);

NOR2xp67_ASAP7_75t_L g1015 ( 
.A(n_917),
.B(n_863),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_822),
.A2(n_826),
.B(n_926),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_833),
.B(n_949),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_954),
.B(n_842),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_808),
.A2(n_938),
.B(n_920),
.C(n_807),
.Y(n_1019)
);

OAI221xp5_ASAP7_75t_L g1020 ( 
.A1(n_928),
.A2(n_839),
.B1(n_907),
.B2(n_819),
.C(n_970),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_973),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_SL g1022 ( 
.A1(n_842),
.A2(n_938),
.B(n_939),
.C(n_829),
.Y(n_1022)
);

BUFx12f_ASAP7_75t_L g1023 ( 
.A(n_828),
.Y(n_1023)
);

NAND2x1p5_ASAP7_75t_L g1024 ( 
.A(n_861),
.B(n_912),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_822),
.A2(n_831),
.B(n_851),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_851),
.A2(n_849),
.B(n_843),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_915),
.A2(n_916),
.B(n_925),
.Y(n_1027)
);

BUFx8_ASAP7_75t_SL g1028 ( 
.A(n_951),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_837),
.A2(n_844),
.B(n_945),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_846),
.B(n_821),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_862),
.Y(n_1031)
);

NOR2x1_ASAP7_75t_SL g1032 ( 
.A(n_889),
.B(n_952),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_819),
.B(n_970),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_929),
.A2(n_835),
.B(n_830),
.Y(n_1034)
);

AOI21xp33_ASAP7_75t_L g1035 ( 
.A1(n_805),
.A2(n_839),
.B(n_818),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_874),
.Y(n_1036)
);

OA21x2_ASAP7_75t_L g1037 ( 
.A1(n_850),
.A2(n_942),
.B(n_900),
.Y(n_1037)
);

AOI21x1_ASAP7_75t_SL g1038 ( 
.A1(n_885),
.A2(n_838),
.B(n_854),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_910),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_SL g1040 ( 
.A(n_863),
.B(n_875),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_857),
.A2(n_906),
.B(n_853),
.Y(n_1041)
);

AOI21xp33_ASAP7_75t_L g1042 ( 
.A1(n_950),
.A2(n_973),
.B(n_825),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_820),
.B(n_912),
.Y(n_1043)
);

NAND3xp33_ASAP7_75t_L g1044 ( 
.A(n_858),
.B(n_875),
.C(n_859),
.Y(n_1044)
);

AOI221xp5_ASAP7_75t_L g1045 ( 
.A1(n_886),
.A2(n_931),
.B1(n_947),
.B2(n_934),
.C(n_935),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_952),
.A2(n_855),
.B(n_869),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_848),
.A2(n_877),
.B(n_867),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_902),
.B(n_861),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_901),
.B(n_821),
.Y(n_1049)
);

OAI21xp33_ASAP7_75t_L g1050 ( 
.A1(n_934),
.A2(n_935),
.B(n_937),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_941),
.B(n_901),
.Y(n_1051)
);

AO31x2_ASAP7_75t_L g1052 ( 
.A1(n_898),
.A2(n_868),
.A3(n_905),
.B(n_882),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_943),
.B(n_921),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_932),
.A2(n_940),
.B(n_866),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_936),
.B(n_871),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_892),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_865),
.A2(n_836),
.B1(n_893),
.B2(n_895),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_864),
.B(n_883),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_899),
.A2(n_823),
.B1(n_870),
.B2(n_953),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_860),
.B(n_514),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_SL g1061 ( 
.A1(n_974),
.A2(n_872),
.B(n_890),
.Y(n_1061)
);

OA21x2_ASAP7_75t_L g1062 ( 
.A1(n_958),
.A2(n_964),
.B(n_963),
.Y(n_1062)
);

O2A1O1Ixp5_ASAP7_75t_L g1063 ( 
.A1(n_840),
.A2(n_851),
.B(n_908),
.C(n_783),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_816),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_847),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_958),
.A2(n_764),
.B(n_668),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_862),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_823),
.B(n_514),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_967),
.A2(n_946),
.B(n_654),
.Y(n_1069)
);

NAND2x1p5_ASAP7_75t_L g1070 ( 
.A(n_847),
.B(n_881),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_968),
.A2(n_815),
.B(n_823),
.C(n_909),
.Y(n_1071)
);

BUFx12f_ASAP7_75t_L g1072 ( 
.A(n_816),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_967),
.A2(n_946),
.B(n_654),
.Y(n_1073)
);

NAND2x1p5_ASAP7_75t_L g1074 ( 
.A(n_847),
.B(n_881),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_968),
.B(n_953),
.Y(n_1075)
);

O2A1O1Ixp5_ASAP7_75t_L g1076 ( 
.A1(n_840),
.A2(n_851),
.B(n_908),
.C(n_783),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_847),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_862),
.Y(n_1078)
);

AOI21xp33_ASAP7_75t_L g1079 ( 
.A1(n_823),
.A2(n_815),
.B(n_667),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_958),
.A2(n_764),
.B(n_668),
.Y(n_1080)
);

OAI21xp33_ASAP7_75t_L g1081 ( 
.A1(n_968),
.A2(n_667),
.B(n_498),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_827),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_862),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_823),
.B(n_514),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_958),
.A2(n_764),
.B(n_668),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_823),
.B(n_514),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_968),
.B(n_953),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_968),
.B(n_953),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_847),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_847),
.Y(n_1090)
);

AOI21x1_ASAP7_75t_L g1091 ( 
.A1(n_826),
.A2(n_879),
.B(n_873),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_968),
.A2(n_815),
.B(n_823),
.C(n_909),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_847),
.B(n_881),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_862),
.Y(n_1094)
);

NOR2x1_ASAP7_75t_L g1095 ( 
.A(n_919),
.B(n_953),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_959),
.A2(n_962),
.B(n_960),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_847),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_958),
.A2(n_764),
.B(n_668),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_959),
.A2(n_962),
.B(n_960),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_968),
.B(n_953),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_865),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_968),
.A2(n_823),
.B1(n_815),
.B2(n_832),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_959),
.A2(n_962),
.B(n_960),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_827),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1079),
.B(n_987),
.Y(n_1105)
);

O2A1O1Ixp5_ASAP7_75t_SL g1106 ( 
.A1(n_1003),
.A2(n_1035),
.B(n_1053),
.C(n_990),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_1009),
.Y(n_1107)
);

INVx3_ASAP7_75t_SL g1108 ( 
.A(n_1101),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_981),
.B(n_989),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_1023),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1068),
.B(n_1084),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_1021),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1017),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_1102),
.B(n_1081),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_1021),
.Y(n_1115)
);

OR2x6_ASAP7_75t_L g1116 ( 
.A(n_1049),
.B(n_1072),
.Y(n_1116)
);

INVx5_ASAP7_75t_L g1117 ( 
.A(n_992),
.Y(n_1117)
);

NAND2x1p5_ASAP7_75t_L g1118 ( 
.A(n_1009),
.B(n_1012),
.Y(n_1118)
);

NOR2xp67_ASAP7_75t_L g1119 ( 
.A(n_1020),
.B(n_1007),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_1028),
.Y(n_1120)
);

OR2x2_ASAP7_75t_L g1121 ( 
.A(n_1086),
.B(n_975),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_983),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_980),
.B(n_1075),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_998),
.Y(n_1124)
);

NOR2xp67_ASAP7_75t_L g1125 ( 
.A(n_1064),
.B(n_979),
.Y(n_1125)
);

AOI21xp33_ASAP7_75t_SL g1126 ( 
.A1(n_1049),
.A2(n_1050),
.B(n_1042),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_1030),
.Y(n_1127)
);

NAND2xp33_ASAP7_75t_L g1128 ( 
.A(n_994),
.B(n_1071),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_SL g1129 ( 
.A1(n_994),
.A2(n_991),
.B(n_1092),
.C(n_1071),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_995),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_976),
.Y(n_1131)
);

AND2x4_ASAP7_75t_SL g1132 ( 
.A(n_1030),
.B(n_1097),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1087),
.B(n_1088),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1100),
.B(n_1092),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_988),
.B(n_986),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1051),
.B(n_1009),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_992),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1013),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1051),
.B(n_1014),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_985),
.B(n_1033),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1009),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_1012),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1045),
.B(n_999),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_991),
.B(n_1018),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1099),
.A2(n_1103),
.B(n_977),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1095),
.B(n_1055),
.Y(n_1146)
);

O2A1O1Ixp5_ASAP7_75t_L g1147 ( 
.A1(n_1063),
.A2(n_1076),
.B(n_1025),
.C(n_1047),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1019),
.A2(n_1080),
.B(n_1098),
.C(n_1085),
.Y(n_1148)
);

BUFx10_ASAP7_75t_L g1149 ( 
.A(n_997),
.Y(n_1149)
);

OR2x6_ASAP7_75t_L g1150 ( 
.A(n_1024),
.B(n_1070),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1039),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1001),
.A2(n_1022),
.B(n_1066),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1022),
.A2(n_1002),
.B(n_1019),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1024),
.A2(n_1006),
.B1(n_1048),
.B2(n_1044),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_1012),
.Y(n_1155)
);

AOI21xp33_ASAP7_75t_L g1156 ( 
.A1(n_1059),
.A2(n_1053),
.B(n_1008),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1061),
.A2(n_996),
.B(n_978),
.C(n_1005),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_996),
.A2(n_1005),
.B(n_1004),
.C(n_1010),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_997),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1043),
.B(n_1062),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_1057),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1062),
.B(n_1060),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_1012),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1015),
.B(n_1040),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_997),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1006),
.B(n_1082),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1104),
.B(n_1036),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1000),
.B(n_984),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1027),
.A2(n_1047),
.B(n_1041),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1031),
.B(n_1083),
.Y(n_1170)
);

CKINVDCx20_ASAP7_75t_R g1171 ( 
.A(n_997),
.Y(n_1171)
);

NOR2x1_ASAP7_75t_L g1172 ( 
.A(n_1097),
.B(n_982),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_982),
.B(n_1077),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_1067),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1078),
.B(n_1094),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1070),
.A2(n_1074),
.B1(n_1093),
.B2(n_1065),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1074),
.A2(n_1093),
.B1(n_1077),
.B2(n_984),
.Y(n_1177)
);

OAI21xp33_ASAP7_75t_L g1178 ( 
.A1(n_1011),
.A2(n_1016),
.B(n_1058),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1063),
.A2(n_1076),
.B(n_1046),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1000),
.B(n_1090),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1065),
.B(n_1089),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1065),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1065),
.A2(n_1089),
.B1(n_1090),
.B2(n_1046),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1032),
.A2(n_1038),
.A3(n_1000),
.B(n_1026),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_1089),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1090),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1090),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1034),
.B(n_1054),
.Y(n_1188)
);

INVx1_ASAP7_75t_SL g1189 ( 
.A(n_1037),
.Y(n_1189)
);

INVxp67_ASAP7_75t_L g1190 ( 
.A(n_1037),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1037),
.B(n_1052),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1091),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_SL g1193 ( 
.A1(n_1038),
.A2(n_1052),
.B(n_993),
.C(n_1056),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_1056),
.B(n_1029),
.Y(n_1194)
);

INVx3_ASAP7_75t_SL g1195 ( 
.A(n_1056),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1069),
.B(n_1073),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1068),
.B(n_1084),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1068),
.B(n_1084),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1009),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1051),
.B(n_1030),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1068),
.B(n_1084),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1068),
.B(n_1084),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1023),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1023),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1079),
.B(n_968),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1068),
.B(n_1084),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1017),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_992),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_992),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1079),
.A2(n_994),
.B(n_968),
.C(n_1071),
.Y(n_1210)
);

NOR2xp67_ASAP7_75t_SL g1211 ( 
.A(n_1023),
.B(n_514),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1079),
.B(n_968),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_990),
.A2(n_1099),
.B(n_1096),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_990),
.A2(n_1099),
.B(n_1096),
.Y(n_1214)
);

NOR2xp67_ASAP7_75t_L g1215 ( 
.A(n_1020),
.B(n_514),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_990),
.A2(n_1099),
.B(n_1096),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1051),
.B(n_1030),
.Y(n_1217)
);

AO32x1_ASAP7_75t_L g1218 ( 
.A1(n_1059),
.A2(n_661),
.A3(n_1010),
.B1(n_685),
.B2(n_956),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1028),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1017),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1023),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1102),
.A2(n_823),
.B1(n_1079),
.B2(n_968),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1102),
.A2(n_823),
.B1(n_1079),
.B2(n_968),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1068),
.B(n_1084),
.Y(n_1224)
);

AO21x2_ASAP7_75t_L g1225 ( 
.A1(n_1025),
.A2(n_1005),
.B(n_977),
.Y(n_1225)
);

INVx6_ASAP7_75t_L g1226 ( 
.A(n_1009),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1068),
.B(n_1084),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1017),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1079),
.B(n_968),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1068),
.B(n_1084),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1021),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1079),
.A2(n_968),
.B1(n_1081),
.B2(n_1003),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1079),
.B(n_968),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1017),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1192),
.Y(n_1235)
);

CKINVDCx6p67_ASAP7_75t_R g1236 ( 
.A(n_1108),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1222),
.A2(n_1223),
.B1(n_1114),
.B2(n_1232),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1171),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1120),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1114),
.A2(n_1232),
.B1(n_1233),
.B2(n_1212),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1124),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1151),
.Y(n_1242)
);

OAI21xp33_ASAP7_75t_L g1243 ( 
.A1(n_1205),
.A2(n_1229),
.B(n_1133),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1142),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_SL g1245 ( 
.A1(n_1161),
.A2(n_1143),
.B1(n_1128),
.B2(n_1164),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1123),
.A2(n_1215),
.B1(n_1119),
.B2(n_1227),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1105),
.B(n_1134),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1156),
.A2(n_1224),
.B1(n_1206),
.B2(n_1230),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1111),
.A2(n_1197),
.B1(n_1198),
.B2(n_1201),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1189),
.Y(n_1250)
);

OAI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1121),
.A2(n_1131),
.B1(n_1135),
.B2(n_1109),
.Y(n_1251)
);

CKINVDCx16_ASAP7_75t_R g1252 ( 
.A(n_1120),
.Y(n_1252)
);

BUFx8_ASAP7_75t_L g1253 ( 
.A(n_1221),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1202),
.A2(n_1146),
.B1(n_1139),
.B2(n_1225),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1167),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1113),
.B(n_1207),
.Y(n_1256)
);

OR2x6_ASAP7_75t_L g1257 ( 
.A(n_1158),
.B(n_1213),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1140),
.B(n_1220),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1225),
.A2(n_1154),
.B1(n_1144),
.B2(n_1178),
.Y(n_1259)
);

OAI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1125),
.A2(n_1234),
.B1(n_1228),
.B2(n_1116),
.Y(n_1260)
);

INVx6_ASAP7_75t_L g1261 ( 
.A(n_1117),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1179),
.A2(n_1147),
.B(n_1169),
.Y(n_1262)
);

BUFx2_ASAP7_75t_R g1263 ( 
.A(n_1219),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1142),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1112),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1200),
.A2(n_1217),
.B1(n_1122),
.B2(n_1130),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1170),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1180),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1200),
.A2(n_1217),
.B1(n_1122),
.B2(n_1152),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1175),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1175),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1112),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1190),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1210),
.B(n_1115),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1190),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1115),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1152),
.A2(n_1211),
.B1(n_1116),
.B2(n_1231),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1127),
.A2(n_1116),
.B1(n_1203),
.B2(n_1110),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1148),
.A2(n_1171),
.B1(n_1210),
.B2(n_1126),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1168),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1142),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1231),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1153),
.A2(n_1150),
.B1(n_1162),
.B2(n_1204),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1166),
.Y(n_1284)
);

BUFx8_ASAP7_75t_L g1285 ( 
.A(n_1159),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1182),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1136),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1108),
.A2(n_1150),
.B1(n_1177),
.B2(n_1174),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1147),
.A2(n_1169),
.B(n_1153),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1142),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1186),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1150),
.A2(n_1176),
.B1(n_1136),
.B2(n_1191),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1187),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1137),
.Y(n_1294)
);

BUFx8_ASAP7_75t_SL g1295 ( 
.A(n_1199),
.Y(n_1295)
);

BUFx2_ASAP7_75t_R g1296 ( 
.A(n_1141),
.Y(n_1296)
);

INVx4_ASAP7_75t_SL g1297 ( 
.A(n_1226),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1160),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1173),
.A2(n_1194),
.B1(n_1188),
.B2(n_1145),
.Y(n_1299)
);

INVx4_ASAP7_75t_R g1300 ( 
.A(n_1141),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1132),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1148),
.B(n_1184),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1173),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1194),
.A2(n_1188),
.B1(n_1145),
.B2(n_1216),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1208),
.Y(n_1305)
);

INVx6_ASAP7_75t_L g1306 ( 
.A(n_1117),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1213),
.A2(n_1214),
.B(n_1193),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1199),
.A2(n_1107),
.B1(n_1155),
.B2(n_1129),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1209),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1106),
.A2(n_1157),
.B(n_1158),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1214),
.A2(n_1165),
.B1(n_1183),
.B2(n_1185),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1196),
.A2(n_1157),
.B(n_1118),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1181),
.B(n_1209),
.Y(n_1313)
);

AOI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1193),
.A2(n_1172),
.B(n_1181),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_1199),
.Y(n_1315)
);

INVx5_ASAP7_75t_L g1316 ( 
.A(n_1117),
.Y(n_1316)
);

AO21x2_ASAP7_75t_L g1317 ( 
.A1(n_1129),
.A2(n_1218),
.B(n_1184),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1195),
.B(n_1118),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1218),
.A2(n_1163),
.B(n_1149),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1123),
.B(n_823),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1213),
.A2(n_1216),
.B(n_1214),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1179),
.A2(n_1147),
.B(n_1169),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1222),
.A2(n_1102),
.B1(n_823),
.B2(n_1079),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1192),
.Y(n_1324)
);

BUFx8_ASAP7_75t_L g1325 ( 
.A(n_1221),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1232),
.A2(n_823),
.B1(n_1102),
.B2(n_1079),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1120),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1138),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1222),
.A2(n_823),
.B1(n_1079),
.B2(n_968),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1162),
.B(n_1123),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1314),
.Y(n_1331)
);

AO21x1_ASAP7_75t_SL g1332 ( 
.A1(n_1237),
.A2(n_1310),
.B(n_1302),
.Y(n_1332)
);

OR2x6_ASAP7_75t_L g1333 ( 
.A(n_1321),
.B(n_1257),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1323),
.A2(n_1329),
.B(n_1326),
.Y(n_1334)
);

AO222x2_ASAP7_75t_L g1335 ( 
.A1(n_1247),
.A2(n_1256),
.B1(n_1240),
.B2(n_1243),
.C1(n_1245),
.C2(n_1249),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1239),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_1296),
.Y(n_1337)
);

INVx2_ASAP7_75t_SL g1338 ( 
.A(n_1265),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1235),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1265),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1324),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1282),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1320),
.A2(n_1246),
.B1(n_1279),
.B2(n_1258),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1291),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1272),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1268),
.B(n_1280),
.Y(n_1346)
);

CKINVDCx6p67_ASAP7_75t_R g1347 ( 
.A(n_1327),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1276),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1251),
.B(n_1256),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_1300),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1273),
.Y(n_1351)
);

BUFx12f_ASAP7_75t_L g1352 ( 
.A(n_1239),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1273),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1299),
.B(n_1275),
.Y(n_1354)
);

INVxp33_ASAP7_75t_L g1355 ( 
.A(n_1238),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1298),
.B(n_1257),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1284),
.B(n_1270),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1250),
.Y(n_1358)
);

AO21x2_ASAP7_75t_L g1359 ( 
.A1(n_1307),
.A2(n_1312),
.B(n_1317),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1259),
.A2(n_1304),
.B(n_1274),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1255),
.Y(n_1361)
);

AOI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1257),
.A2(n_1318),
.B(n_1289),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1248),
.A2(n_1260),
.B1(n_1288),
.B2(n_1269),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1330),
.B(n_1257),
.Y(n_1364)
);

INVx5_ASAP7_75t_L g1365 ( 
.A(n_1316),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1330),
.B(n_1254),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1262),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1313),
.B(n_1262),
.Y(n_1368)
);

BUFx4f_ASAP7_75t_SL g1369 ( 
.A(n_1327),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1322),
.Y(n_1370)
);

OR2x2_ASAP7_75t_SL g1371 ( 
.A(n_1252),
.B(n_1322),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1319),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1307),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1267),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1236),
.A2(n_1278),
.B1(n_1238),
.B2(n_1271),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1241),
.B(n_1242),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1283),
.B(n_1292),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1277),
.B(n_1328),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1311),
.B(n_1287),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1319),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1286),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1266),
.B(n_1303),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1287),
.B(n_1293),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1253),
.A2(n_1325),
.B1(n_1306),
.B2(n_1261),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1368),
.B(n_1294),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1356),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1356),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1371),
.B(n_1318),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1356),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1364),
.B(n_1309),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_SL g1391 ( 
.A(n_1343),
.B(n_1375),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1364),
.B(n_1305),
.Y(n_1392)
);

OAI222xp33_ASAP7_75t_L g1393 ( 
.A1(n_1363),
.A2(n_1308),
.B1(n_1316),
.B2(n_1301),
.C1(n_1315),
.C2(n_1236),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1333),
.B(n_1244),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1346),
.B(n_1244),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1333),
.B(n_1297),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1373),
.B(n_1244),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1373),
.B(n_1290),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1360),
.B(n_1290),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1360),
.B(n_1290),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1345),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1339),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1359),
.B(n_1264),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1348),
.Y(n_1404)
);

AND2x2_ASAP7_75t_SL g1405 ( 
.A(n_1360),
.B(n_1264),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1341),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1338),
.Y(n_1407)
);

INVxp67_ASAP7_75t_SL g1408 ( 
.A(n_1367),
.Y(n_1408)
);

NAND2x1p5_ASAP7_75t_SL g1409 ( 
.A(n_1340),
.B(n_1366),
.Y(n_1409)
);

INVx4_ASAP7_75t_L g1410 ( 
.A(n_1365),
.Y(n_1410)
);

INVxp67_ASAP7_75t_SL g1411 ( 
.A(n_1367),
.Y(n_1411)
);

AOI32xp33_ASAP7_75t_L g1412 ( 
.A1(n_1335),
.A2(n_1301),
.A3(n_1295),
.B1(n_1325),
.B2(n_1253),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1334),
.A2(n_1253),
.B1(n_1325),
.B2(n_1285),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1370),
.B(n_1281),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1380),
.B(n_1281),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1401),
.B(n_1366),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1391),
.B(n_1355),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_SL g1418 ( 
.A(n_1412),
.B(n_1349),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_SL g1419 ( 
.A(n_1393),
.B(n_1365),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1401),
.B(n_1351),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1385),
.B(n_1362),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1385),
.B(n_1362),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1385),
.B(n_1372),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1404),
.B(n_1351),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1413),
.B(n_1347),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1404),
.B(n_1353),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1386),
.B(n_1360),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1393),
.A2(n_1365),
.B(n_1316),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1402),
.B(n_1406),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_SL g1430 ( 
.A(n_1410),
.B(n_1365),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1414),
.B(n_1332),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1390),
.B(n_1342),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1414),
.B(n_1332),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1415),
.Y(n_1434)
);

OAI221xp5_ASAP7_75t_L g1435 ( 
.A1(n_1412),
.A2(n_1363),
.B1(n_1384),
.B2(n_1382),
.C(n_1378),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1413),
.A2(n_1377),
.B1(n_1347),
.B2(n_1357),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_L g1437 ( 
.A(n_1399),
.B(n_1378),
.C(n_1377),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1392),
.B(n_1395),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1392),
.B(n_1369),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1396),
.A2(n_1379),
.B1(n_1354),
.B2(n_1352),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1397),
.B(n_1354),
.Y(n_1441)
);

NAND3xp33_ASAP7_75t_L g1442 ( 
.A(n_1399),
.B(n_1344),
.C(n_1374),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1395),
.B(n_1358),
.Y(n_1443)
);

NAND3xp33_ASAP7_75t_L g1444 ( 
.A(n_1400),
.B(n_1383),
.C(n_1361),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1398),
.B(n_1331),
.Y(n_1445)
);

NAND4xp25_ASAP7_75t_L g1446 ( 
.A(n_1400),
.B(n_1376),
.C(n_1337),
.D(n_1381),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1396),
.A2(n_1379),
.B(n_1350),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1396),
.B(n_1336),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1429),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1429),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1434),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1417),
.B(n_1352),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1416),
.B(n_1408),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1416),
.B(n_1409),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1421),
.B(n_1408),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1421),
.B(n_1411),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1422),
.B(n_1411),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1422),
.B(n_1437),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1420),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1423),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1445),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1437),
.B(n_1409),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1431),
.B(n_1387),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1420),
.Y(n_1464)
);

AND2x4_ASAP7_75t_SL g1465 ( 
.A(n_1431),
.B(n_1396),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1433),
.B(n_1389),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1424),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1433),
.B(n_1389),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1424),
.B(n_1407),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1426),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1442),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1438),
.B(n_1409),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1426),
.B(n_1444),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1427),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1444),
.B(n_1407),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1441),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1442),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1461),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1458),
.B(n_1432),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1455),
.Y(n_1480)
);

NOR2x1_ASAP7_75t_L g1481 ( 
.A(n_1462),
.B(n_1446),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1449),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1449),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1476),
.B(n_1405),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1471),
.B(n_1443),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1450),
.Y(n_1486)
);

INVx3_ASAP7_75t_SL g1487 ( 
.A(n_1462),
.Y(n_1487)
);

NAND2x1p5_ASAP7_75t_L g1488 ( 
.A(n_1454),
.B(n_1410),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1461),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1465),
.B(n_1396),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1450),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1451),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1465),
.B(n_1403),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_SL g1494 ( 
.A(n_1471),
.B(n_1419),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1451),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1465),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1461),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1459),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1476),
.B(n_1405),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_R g1500 ( 
.A(n_1452),
.B(n_1425),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1459),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1463),
.B(n_1394),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1455),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1473),
.B(n_1477),
.Y(n_1504)
);

INVxp67_ASAP7_75t_SL g1505 ( 
.A(n_1475),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1464),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1464),
.Y(n_1507)
);

NAND3xp33_ASAP7_75t_L g1508 ( 
.A(n_1473),
.B(n_1418),
.C(n_1435),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1467),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1467),
.Y(n_1510)
);

NAND2x1p5_ASAP7_75t_L g1511 ( 
.A(n_1454),
.B(n_1410),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1482),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1508),
.B(n_1475),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1482),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1496),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1496),
.B(n_1474),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1496),
.B(n_1466),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1508),
.B(n_1439),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1492),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1487),
.B(n_1493),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1504),
.B(n_1472),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1485),
.B(n_1472),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1505),
.B(n_1458),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1483),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1493),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1487),
.B(n_1468),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1505),
.B(n_1456),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1485),
.B(n_1470),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1483),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1487),
.B(n_1470),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1492),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1495),
.Y(n_1532)
);

OAI21xp33_ASAP7_75t_L g1533 ( 
.A1(n_1481),
.A2(n_1446),
.B(n_1419),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1486),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1481),
.B(n_1469),
.Y(n_1535)
);

AOI21xp33_ASAP7_75t_SL g1536 ( 
.A1(n_1488),
.A2(n_1436),
.B(n_1448),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1478),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1486),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1479),
.B(n_1456),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1478),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1478),
.Y(n_1541)
);

CKINVDCx16_ASAP7_75t_R g1542 ( 
.A(n_1494),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1491),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1495),
.Y(n_1544)
);

AND2x4_ASAP7_75t_SL g1545 ( 
.A(n_1490),
.B(n_1460),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1489),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1491),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1479),
.B(n_1457),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1489),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1498),
.Y(n_1550)
);

AND2x2_ASAP7_75t_SL g1551 ( 
.A(n_1494),
.B(n_1430),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1489),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1498),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1480),
.B(n_1469),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1520),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1518),
.B(n_1263),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_1515),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1542),
.B(n_1488),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1513),
.B(n_1480),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1533),
.A2(n_1436),
.B(n_1488),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1526),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1519),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1512),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1515),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1520),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1551),
.A2(n_1503),
.B1(n_1511),
.B2(n_1440),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1526),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1522),
.B(n_1503),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1512),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1514),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1516),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1525),
.B(n_1490),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1523),
.B(n_1497),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1551),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1514),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1516),
.Y(n_1576)
);

OR2x6_ASAP7_75t_L g1577 ( 
.A(n_1530),
.B(n_1428),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1524),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1545),
.B(n_1511),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1545),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1517),
.B(n_1511),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1535),
.B(n_1502),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1523),
.B(n_1497),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1544),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1521),
.Y(n_1585)
);

NAND3xp33_ASAP7_75t_L g1586 ( 
.A(n_1536),
.B(n_1506),
.C(n_1501),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1524),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1539),
.B(n_1497),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1529),
.Y(n_1589)
);

AND2x4_ASAP7_75t_SL g1590 ( 
.A(n_1517),
.B(n_1490),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1563),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1586),
.A2(n_1528),
.B(n_1554),
.Y(n_1592)
);

OAI21xp33_ASAP7_75t_L g1593 ( 
.A1(n_1574),
.A2(n_1500),
.B(n_1527),
.Y(n_1593)
);

OAI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1585),
.A2(n_1500),
.B1(n_1527),
.B2(n_1388),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1555),
.B(n_1531),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1557),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1565),
.B(n_1532),
.Y(n_1597)
);

AND2x4_ASAP7_75t_SL g1598 ( 
.A(n_1558),
.B(n_1350),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1567),
.B(n_1539),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1563),
.Y(n_1600)
);

AOI332xp33_ASAP7_75t_L g1601 ( 
.A1(n_1562),
.A2(n_1553),
.A3(n_1529),
.B1(n_1550),
.B2(n_1534),
.B3(n_1538),
.C1(n_1547),
.C2(n_1543),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1569),
.Y(n_1602)
);

AOI21xp33_ASAP7_75t_L g1603 ( 
.A1(n_1580),
.A2(n_1558),
.B(n_1559),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1557),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1569),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1584),
.B(n_1548),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1561),
.B(n_1562),
.Y(n_1607)
);

AOI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1560),
.A2(n_1525),
.B(n_1534),
.Y(n_1608)
);

NOR2x2_ASAP7_75t_L g1609 ( 
.A(n_1561),
.B(n_1537),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1570),
.Y(n_1610)
);

INVxp67_ASAP7_75t_SL g1611 ( 
.A(n_1564),
.Y(n_1611)
);

OAI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1577),
.A2(n_1564),
.B1(n_1568),
.B2(n_1571),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1566),
.A2(n_1447),
.B1(n_1516),
.B2(n_1490),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1570),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1582),
.B(n_1548),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_SL g1616 ( 
.A1(n_1577),
.A2(n_1430),
.B1(n_1553),
.B2(n_1550),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1611),
.B(n_1571),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1611),
.B(n_1576),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1593),
.A2(n_1577),
.B1(n_1581),
.B2(n_1590),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1591),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1600),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1596),
.B(n_1576),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1604),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1602),
.Y(n_1624)
);

AO22x2_ASAP7_75t_L g1625 ( 
.A1(n_1605),
.A2(n_1578),
.B1(n_1587),
.B2(n_1575),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1598),
.B(n_1590),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1603),
.B(n_1581),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1607),
.B(n_1568),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1608),
.B(n_1589),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1613),
.B(n_1572),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1594),
.B(n_1579),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1599),
.B(n_1572),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1610),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1609),
.Y(n_1634)
);

AND2x2_ASAP7_75t_SL g1635 ( 
.A(n_1606),
.B(n_1556),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1595),
.Y(n_1636)
);

NAND3xp33_ASAP7_75t_L g1637 ( 
.A(n_1623),
.B(n_1616),
.C(n_1592),
.Y(n_1637)
);

AOI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1617),
.A2(n_1614),
.B(n_1597),
.Y(n_1638)
);

OAI31xp33_ASAP7_75t_SL g1639 ( 
.A1(n_1634),
.A2(n_1594),
.A3(n_1612),
.B(n_1616),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1631),
.A2(n_1629),
.B(n_1635),
.Y(n_1640)
);

AOI221xp5_ASAP7_75t_L g1641 ( 
.A1(n_1636),
.A2(n_1612),
.B1(n_1628),
.B2(n_1627),
.C(n_1618),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1635),
.A2(n_1577),
.B1(n_1615),
.B2(n_1579),
.Y(n_1642)
);

AOI221x1_ASAP7_75t_L g1643 ( 
.A1(n_1625),
.A2(n_1589),
.B1(n_1575),
.B2(n_1587),
.C(n_1578),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1627),
.A2(n_1601),
.B(n_1583),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1625),
.A2(n_1583),
.B(n_1573),
.Y(n_1645)
);

AOI21xp33_ASAP7_75t_SL g1646 ( 
.A1(n_1622),
.A2(n_1632),
.B(n_1630),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1625),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1625),
.A2(n_1573),
.B(n_1572),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1646),
.B(n_1632),
.Y(n_1649)
);

NAND3xp33_ASAP7_75t_L g1650 ( 
.A(n_1639),
.B(n_1619),
.C(n_1630),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1641),
.B(n_1620),
.Y(n_1651)
);

AO22x2_ASAP7_75t_L g1652 ( 
.A1(n_1647),
.A2(n_1633),
.B1(n_1624),
.B2(n_1620),
.Y(n_1652)
);

NOR2x1p5_ASAP7_75t_L g1653 ( 
.A(n_1637),
.B(n_1621),
.Y(n_1653)
);

NOR3x1_ASAP7_75t_L g1654 ( 
.A(n_1640),
.B(n_1624),
.C(n_1621),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1643),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1638),
.B(n_1644),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1648),
.B(n_1633),
.Y(n_1657)
);

NAND3xp33_ASAP7_75t_SL g1658 ( 
.A(n_1642),
.B(n_1626),
.C(n_1588),
.Y(n_1658)
);

AOI211xp5_ASAP7_75t_L g1659 ( 
.A1(n_1656),
.A2(n_1645),
.B(n_1626),
.C(n_1572),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_SL g1660 ( 
.A(n_1650),
.B(n_1588),
.Y(n_1660)
);

NOR3xp33_ASAP7_75t_L g1661 ( 
.A(n_1658),
.B(n_1543),
.C(n_1538),
.Y(n_1661)
);

XNOR2xp5_ASAP7_75t_L g1662 ( 
.A(n_1649),
.B(n_1493),
.Y(n_1662)
);

NOR4xp25_ASAP7_75t_L g1663 ( 
.A(n_1655),
.B(n_1547),
.C(n_1549),
.D(n_1552),
.Y(n_1663)
);

AOI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1660),
.A2(n_1651),
.B1(n_1653),
.B2(n_1652),
.Y(n_1664)
);

NOR2xp67_ASAP7_75t_L g1665 ( 
.A(n_1662),
.B(n_1657),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1661),
.B(n_1654),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1659),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1663),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1662),
.Y(n_1669)
);

NOR2x1_ASAP7_75t_L g1670 ( 
.A(n_1668),
.B(n_1665),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1667),
.B(n_1652),
.Y(n_1671)
);

XNOR2xp5_ASAP7_75t_L g1672 ( 
.A(n_1664),
.B(n_1493),
.Y(n_1672)
);

AOI322xp5_ASAP7_75t_L g1673 ( 
.A1(n_1666),
.A2(n_1669),
.A3(n_1552),
.B1(n_1549),
.B2(n_1546),
.C1(n_1541),
.C2(n_1540),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1667),
.Y(n_1674)
);

INVxp33_ASAP7_75t_L g1675 ( 
.A(n_1672),
.Y(n_1675)
);

NOR3xp33_ASAP7_75t_SL g1676 ( 
.A(n_1674),
.B(n_1447),
.C(n_1453),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1671),
.B(n_1670),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1677),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1678),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1679),
.A2(n_1675),
.B1(n_1673),
.B2(n_1676),
.Y(n_1680)
);

XNOR2xp5_ASAP7_75t_L g1681 ( 
.A(n_1679),
.B(n_1537),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1681),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_SL g1683 ( 
.A1(n_1680),
.A2(n_1546),
.B1(n_1541),
.B2(n_1540),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1683),
.B(n_1501),
.Y(n_1684)
);

AOI211xp5_ASAP7_75t_L g1685 ( 
.A1(n_1682),
.A2(n_1510),
.B(n_1509),
.C(n_1506),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1684),
.A2(n_1510),
.B1(n_1509),
.B2(n_1507),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1686),
.Y(n_1687)
);

OAI221xp5_ASAP7_75t_R g1688 ( 
.A1(n_1687),
.A2(n_1685),
.B1(n_1295),
.B2(n_1507),
.C(n_1285),
.Y(n_1688)
);

AOI211xp5_ASAP7_75t_L g1689 ( 
.A1(n_1688),
.A2(n_1484),
.B(n_1499),
.C(n_1453),
.Y(n_1689)
);


endmodule