module real_jpeg_14921_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_176;
wire n_288;
wire n_221;
wire n_215;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_285;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_3),
.B(n_32),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_3),
.B(n_50),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_3),
.B(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_3),
.B(n_44),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_4),
.B(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_4),
.B(n_53),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_4),
.B(n_50),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_4),
.B(n_61),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_4),
.B(n_30),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_5),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_5),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_5),
.B(n_53),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_5),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_5),
.B(n_32),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_5),
.B(n_61),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_8),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_8),
.B(n_53),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_8),
.B(n_44),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_8),
.B(n_50),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_8),
.B(n_63),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_9),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_9),
.B(n_63),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_13),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_13),
.B(n_44),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_13),
.B(n_30),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_13),
.B(n_50),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_13),
.B(n_61),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_13),
.B(n_53),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_13),
.B(n_32),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_14),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_14),
.B(n_44),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_14),
.B(n_50),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_14),
.B(n_63),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_14),
.B(n_32),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_14),
.B(n_61),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_14),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_15),
.B(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_15),
.B(n_30),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_15),
.B(n_50),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_158),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_157),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_20),
.B(n_122),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_85),
.C(n_100),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_21),
.B(n_85),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_54),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_22),
.B(n_55),
.C(n_72),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.C(n_47),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_23),
.B(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_24),
.B(n_29),
.C(n_36),
.Y(n_99)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_29),
.B(n_154),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_29),
.A2(n_35),
.B1(n_153),
.B2(n_154),
.Y(n_235)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_33),
.B(n_46),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_33),
.B(n_67),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_37),
.A2(n_38),
.B1(n_47),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_38),
.A2(n_39),
.B(n_42),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_40),
.B(n_112),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_40),
.B(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_46),
.B(n_111),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_47),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.C(n_52),
.Y(n_47)
);

FAx1_ASAP7_75t_SL g103 ( 
.A(n_48),
.B(n_49),
.CI(n_52),
.CON(n_103),
.SN(n_103)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_72),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_68),
.C(n_70),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_56),
.B(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.C(n_65),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_57),
.A2(n_58),
.B1(n_83),
.B2(n_84),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_57),
.A2(n_58),
.B1(n_62),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_60),
.B(n_67),
.Y(n_252)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_62),
.Y(n_172)
);

INVx5_ASAP7_75t_SL g111 ( 
.A(n_63),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_65),
.B(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_66),
.B(n_112),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_68),
.A2(n_70),
.B1(n_71),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_78),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_75),
.B(n_76),
.C(n_78),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_76),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_79),
.B(n_82),
.C(n_83),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_81),
.A2(n_82),
.B1(n_105),
.B2(n_106),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_83),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_83),
.A2(n_84),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_83),
.B(n_222),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_93),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_94),
.C(n_99),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_87),
.B(n_90),
.C(n_91),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.C(n_98),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_97),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_100),
.B(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_114),
.C(n_117),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_101),
.B(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.C(n_107),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_102),
.A2(n_103),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_103),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_104),
.B(n_107),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.C(n_113),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_108),
.A2(n_109),
.B1(n_113),
.B2(n_198),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_110),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_113),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_114),
.B(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_156),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_146),
.B2(n_147),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_136),
.B2(n_137),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_144),
.B2(n_145),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_152),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_207),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_183),
.B(n_206),
.Y(n_160)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_161),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_181),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_162),
.B(n_181),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_169),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_166),
.B1(n_169),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.C(n_180),
.Y(n_169)
);

FAx1_ASAP7_75t_SL g189 ( 
.A(n_170),
.B(n_173),
.CI(n_180),
.CON(n_189),
.SN(n_189)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_178),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_174),
.A2(n_175),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_184),
.B(n_187),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_194),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_188),
.A2(n_189),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_189),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_190),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_286)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.C(n_200),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_196),
.B(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_199),
.B(n_200),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.C(n_204),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_288),
.C(n_289),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_282),
.B(n_287),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_267),
.B(n_281),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_237),
.B(n_266),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_224),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_212),
.B(n_224),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.C(n_221),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_227),
.B1(n_228),
.B2(n_230),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_213),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_213),
.B(n_263),
.Y(n_262)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.CI(n_216),
.CON(n_213),
.SN(n_213)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_219),
.B(n_220),
.Y(n_246)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_221),
.Y(n_264)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_231),
.B2(n_236),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_230),
.C(n_236),
.Y(n_268)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_228),
.Y(n_230)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_231),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_232),
.B(n_234),
.C(n_235),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_260),
.B(n_265),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_250),
.B(n_259),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_245),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_240),
.B(n_245),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_248),
.C(n_249),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_254),
.B(n_258),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_252),
.B(n_253),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_268),
.B(n_269),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_273),
.B2(n_274),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_275),
.C(n_280),
.Y(n_283)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_279),
.B2(n_280),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_283),
.B(n_284),
.Y(n_287)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);


endmodule