module real_jpeg_12372_n_16 (n_396, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_397, n_3, n_10, n_9, n_16);

input n_396;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_397;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_0),
.Y(n_104)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_3),
.B(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_3),
.B(n_104),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_3),
.B(n_91),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_3),
.B(n_25),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_3),
.B(n_28),
.Y(n_342)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_5),
.B(n_28),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_5),
.B(n_49),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_5),
.B(n_25),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_5),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_5),
.B(n_37),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_6),
.B(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_6),
.B(n_49),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_6),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_6),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_6),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_6),
.B(n_37),
.Y(n_324)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_8),
.B(n_31),
.Y(n_126)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_8),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_8),
.B(n_104),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_8),
.B(n_28),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_8),
.B(n_37),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_8),
.B(n_42),
.Y(n_303)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_28),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_10),
.B(n_49),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_10),
.B(n_37),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_10),
.B(n_25),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_10),
.B(n_104),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_10),
.B(n_91),
.Y(n_205)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_11),
.B(n_91),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_11),
.B(n_31),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_11),
.B(n_28),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_11),
.B(n_49),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_11),
.B(n_37),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_13),
.B(n_25),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_13),
.B(n_28),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_13),
.B(n_91),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_13),
.B(n_31),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_13),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_13),
.B(n_49),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_13),
.B(n_37),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_13),
.B(n_42),
.Y(n_274)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_14),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_14),
.B(n_91),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_14),
.B(n_31),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_14),
.B(n_25),
.Y(n_322)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_15),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_116),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_115),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_75),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_20),
.B(n_75),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_60),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_44),
.C(n_51),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_22),
.B(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_32),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_23),
.B(n_34),
.C(n_38),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.C(n_30),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_24),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_53),
.C(n_58),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_24),
.A2(n_30),
.B1(n_59),
.B2(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_24),
.A2(n_59),
.B1(n_105),
.B2(n_106),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_24),
.B(n_105),
.C(n_249),
.Y(n_269)
);

INVx5_ASAP7_75t_SL g145 ( 
.A(n_25),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_27),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_27),
.A2(n_79),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_27),
.B(n_287),
.C(n_290),
.Y(n_335)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_29),
.B(n_35),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_30),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_30),
.B(n_89),
.C(n_94),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_30),
.A2(n_82),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_30),
.B(n_197),
.C(n_199),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_30),
.A2(n_82),
.B1(n_89),
.B2(n_90),
.Y(n_369)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_35),
.B(n_133),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_40),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_40),
.B(n_107),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_41),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_41),
.B(n_176),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_41),
.B(n_134),
.Y(n_326)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_44),
.A2(n_51),
.B1(n_52),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.C(n_48),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_45),
.B(n_48),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_46),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_46),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_47),
.B(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_53),
.A2(n_54),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_103),
.C(n_105),
.Y(n_102)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_58),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_57),
.A2(n_58),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_58),
.B(n_94),
.C(n_261),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_74),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_69),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_63),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_85),
.C(n_86),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_63),
.A2(n_67),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_64),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_65),
.A2(n_66),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_66),
.B(n_300),
.C(n_302),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_110),
.C(n_111),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_76),
.B(n_389),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_95),
.C(n_99),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_77),
.B(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_84),
.C(n_88),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_85),
.B(n_86),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_87),
.B(n_131),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_101),
.C(n_108),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_89),
.A2(n_90),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_89),
.A2(n_90),
.B1(n_342),
.B2(n_343),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_89),
.A2(n_90),
.B1(n_108),
.B2(n_357),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_90),
.B(n_157),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_90),
.B(n_340),
.C(n_342),
.Y(n_358)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_92),
.B(n_176),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_94),
.A2(n_258),
.B1(n_259),
.B2(n_262),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_94),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_94),
.A2(n_262),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_95),
.A2(n_99),
.B1(n_100),
.B2(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_95),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_97),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_101),
.A2(n_102),
.B1(n_355),
.B2(n_356),
.Y(n_354)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_103),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_103),
.B(n_136),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_103),
.A2(n_138),
.B1(n_204),
.B2(n_205),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_103),
.A2(n_105),
.B1(n_106),
.B2(n_138),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_103),
.B(n_205),
.C(n_303),
.Y(n_340)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_107),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_108),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_110),
.Y(n_390)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI321xp33_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_379),
.A3(n_387),
.B1(n_391),
.B2(n_392),
.C(n_396),
.Y(n_116)
);

AOI321xp33_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_311),
.A3(n_345),
.B1(n_373),
.B2(n_378),
.C(n_397),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_252),
.C(n_306),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_223),
.B(n_251),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_191),
.B(n_222),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_160),
.B(n_190),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_139),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_123),
.B(n_139),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.C(n_135),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_142),
.B1(n_143),
.B2(n_151),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_124),
.B(n_187),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_126),
.CI(n_127),
.CON(n_124),
.SN(n_124)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_128),
.A2(n_129),
.B1(n_135),
.B2(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_130),
.B(n_132),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_133),
.B(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_134),
.B(n_145),
.Y(n_197)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_152),
.B2(n_159),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_142),
.B(n_151),
.C(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_144),
.B(n_147),
.C(n_150),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_149),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_153),
.B(n_155),
.C(n_156),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_157),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_157),
.A2(n_158),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_157),
.B(n_274),
.C(n_277),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_184),
.B(n_189),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_173),
.B(n_183),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_168),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_163),
.B(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_171),
.C(n_172),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_178),
.B(n_182),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_175),
.B(n_177),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_185),
.B(n_186),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_192),
.B(n_193),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_208),
.B2(n_209),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_210),
.C(n_221),
.Y(n_224)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_202),
.C(n_203),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_206),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_220),
.B2(n_221),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_219),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_216),
.C(n_218),
.Y(n_242)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_214),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_215),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_224),
.B(n_225),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_241),
.B2(n_250),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_240),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_228),
.B(n_240),
.C(n_250),
.Y(n_307)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_236),
.B2(n_237),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_231),
.B(n_238),
.C(n_239),
.Y(n_270)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g394 ( 
.A(n_232),
.Y(n_394)
);

FAx1_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_234),
.CI(n_235),
.CON(n_232),
.SN(n_232)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_233),
.B(n_234),
.C(n_235),
.Y(n_279)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_241),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_243),
.CI(n_247),
.CON(n_241),
.SN(n_241)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_242),
.B(n_243),
.C(n_247),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B(n_246),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_245),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_246),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_246),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI21xp33_ASAP7_75t_L g374 ( 
.A1(n_253),
.A2(n_375),
.B(n_376),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_283),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_254),
.B(n_283),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_271),
.C(n_282),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_255),
.B(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_270),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_263),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_257),
.B(n_263),
.C(n_270),
.Y(n_305)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_260),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_269),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_267),
.C(n_269),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_271),
.A2(n_272),
.B1(n_282),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_278),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_279),
.C(n_281),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_276),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_279),
.Y(n_280)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_305),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_294),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_294),
.C(n_305),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_291),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_292),
.C(n_293),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_297),
.C(n_298),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_302),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_300),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_307),
.B(n_308),
.Y(n_375)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_312),
.A2(n_374),
.B(n_377),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_313),
.B(n_314),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_344),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_316),
.B(n_317),
.C(n_344),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_336),
.B2(n_337),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_318),
.B(n_338),
.C(n_339),
.Y(n_372)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_328),
.B2(n_329),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_320),
.B(n_330),
.C(n_335),
.Y(n_351)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_322),
.B(n_324),
.C(n_326),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_326),
.B2(n_327),
.Y(n_323)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_324),
.Y(n_327)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_330),
.A2(n_331),
.B1(n_334),
.B2(n_335),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_332),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_342),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_346),
.B(n_347),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_372),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_359),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_349),
.B(n_359),
.C(n_372),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_351),
.B1(n_352),
.B2(n_353),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_350),
.B(n_354),
.C(n_358),
.Y(n_386)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_358),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_361),
.B1(n_364),
.B2(n_365),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_360),
.B(n_366),
.C(n_371),
.Y(n_382)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_370),
.B2(n_371),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_371),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_380),
.B(n_381),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_388),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_383),
.CI(n_386),
.CON(n_381),
.SN(n_381)
);


endmodule