module real_aes_8520_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_168;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g115 ( .A(n_0), .Y(n_115) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_1), .A2(n_160), .B(n_163), .C(n_243), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_2), .A2(n_189), .B(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g490 ( .A(n_3), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_4), .B(n_219), .Y(n_218) );
AOI21xp33_ASAP7_75t_L g473 ( .A1(n_5), .A2(n_189), .B(n_474), .Y(n_473) );
AND2x6_ASAP7_75t_L g160 ( .A(n_6), .B(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g256 ( .A(n_7), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_8), .B(n_42), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_9), .A2(n_188), .B(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_10), .B(n_172), .Y(n_245) );
INVx1_ASAP7_75t_L g478 ( .A(n_11), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_12), .B(n_213), .Y(n_513) );
INVx1_ASAP7_75t_L g152 ( .A(n_13), .Y(n_152) );
INVx1_ASAP7_75t_L g525 ( .A(n_14), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_15), .A2(n_79), .B1(n_133), .B2(n_134), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_15), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_16), .A2(n_197), .B(n_278), .C(n_280), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_17), .B(n_219), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_18), .B(n_456), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_19), .B(n_189), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_20), .B(n_203), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_21), .A2(n_213), .B(n_264), .C(n_266), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_22), .B(n_219), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_23), .B(n_172), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_24), .A2(n_199), .B(n_280), .C(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_25), .B(n_172), .Y(n_227) );
CKINVDCx16_ASAP7_75t_R g154 ( .A(n_26), .Y(n_154) );
INVx1_ASAP7_75t_L g226 ( .A(n_27), .Y(n_226) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_28), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_29), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_30), .B(n_172), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_31), .A2(n_104), .B1(n_117), .B2(n_744), .Y(n_103) );
INVx1_ASAP7_75t_L g195 ( .A(n_32), .Y(n_195) );
INVx1_ASAP7_75t_L g468 ( .A(n_33), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_34), .A2(n_130), .B1(n_131), .B2(n_132), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_34), .Y(n_130) );
INVx2_ASAP7_75t_L g158 ( .A(n_35), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_36), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_37), .A2(n_213), .B(n_214), .C(n_216), .Y(n_212) );
INVxp67_ASAP7_75t_L g198 ( .A(n_38), .Y(n_198) );
CKINVDCx14_ASAP7_75t_R g211 ( .A(n_39), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_40), .A2(n_163), .B(n_225), .C(n_229), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_41), .A2(n_160), .B(n_163), .C(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g467 ( .A(n_43), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_44), .A2(n_174), .B(n_254), .C(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_45), .B(n_172), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_46), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_47), .Y(n_191) );
INVx1_ASAP7_75t_L g262 ( .A(n_48), .Y(n_262) );
CKINVDCx16_ASAP7_75t_R g469 ( .A(n_49), .Y(n_469) );
OAI22xp5_ASAP7_75t_SL g738 ( .A1(n_50), .A2(n_59), .B1(n_739), .B2(n_740), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_50), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_51), .B(n_189), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_52), .A2(n_163), .B1(n_266), .B2(n_466), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_53), .Y(n_505) );
CKINVDCx16_ASAP7_75t_R g487 ( .A(n_54), .Y(n_487) );
CKINVDCx14_ASAP7_75t_R g252 ( .A(n_55), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_56), .A2(n_216), .B(n_254), .C(n_477), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_57), .Y(n_537) );
INVx1_ASAP7_75t_L g475 ( .A(n_58), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_59), .Y(n_740) );
INVx1_ASAP7_75t_L g161 ( .A(n_60), .Y(n_161) );
INVx1_ASAP7_75t_L g151 ( .A(n_61), .Y(n_151) );
INVx1_ASAP7_75t_SL g215 ( .A(n_62), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_63), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g737 ( .A1(n_64), .A2(n_738), .B1(n_741), .B2(n_742), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_64), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_65), .B(n_219), .Y(n_268) );
INVx1_ASAP7_75t_L g167 ( .A(n_66), .Y(n_167) );
AOI222xp33_ASAP7_75t_SL g127 ( .A1(n_67), .A2(n_128), .B1(n_129), .B2(n_135), .C1(n_729), .C2(n_731), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_SL g455 ( .A1(n_68), .A2(n_216), .B(n_456), .C(n_457), .Y(n_455) );
INVxp67_ASAP7_75t_L g458 ( .A(n_69), .Y(n_458) );
INVx1_ASAP7_75t_L g110 ( .A(n_70), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_71), .A2(n_189), .B(n_251), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_72), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_73), .A2(n_189), .B(n_275), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_74), .Y(n_471) );
INVx1_ASAP7_75t_L g531 ( .A(n_75), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_76), .A2(n_188), .B(n_190), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g223 ( .A(n_77), .Y(n_223) );
INVx1_ASAP7_75t_L g276 ( .A(n_78), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_79), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_80), .A2(n_160), .B(n_163), .C(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_81), .A2(n_189), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g279 ( .A(n_82), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_83), .B(n_196), .Y(n_502) );
INVx2_ASAP7_75t_L g149 ( .A(n_84), .Y(n_149) );
INVx1_ASAP7_75t_L g244 ( .A(n_85), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_86), .B(n_456), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_87), .A2(n_160), .B(n_163), .C(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g112 ( .A(n_88), .B(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g442 ( .A(n_88), .B(n_114), .Y(n_442) );
INVx2_ASAP7_75t_L g728 ( .A(n_88), .Y(n_728) );
A2O1A1Ixp33_ASAP7_75t_L g162 ( .A1(n_89), .A2(n_163), .B(n_166), .C(n_176), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_90), .B(n_181), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_91), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_92), .A2(n_160), .B(n_163), .C(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_93), .Y(n_517) );
INVx1_ASAP7_75t_L g454 ( .A(n_94), .Y(n_454) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_95), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_96), .B(n_196), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_97), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_98), .B(n_147), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_99), .B(n_147), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_100), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g265 ( .A(n_101), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_102), .A2(n_189), .B(n_453), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx6p67_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g745 ( .A(n_107), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_112), .Y(n_125) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_112), .Y(n_743) );
NOR2x2_ASAP7_75t_L g733 ( .A(n_113), .B(n_728), .Y(n_733) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OR2x2_ASAP7_75t_L g727 ( .A(n_114), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_127), .B1(n_734), .B2(n_735), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_124), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_SL g734 ( .A(n_122), .Y(n_734) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_124), .A2(n_736), .B(n_743), .Y(n_735) );
NOR2xp33_ASAP7_75t_SL g124 ( .A(n_125), .B(n_126), .Y(n_124) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OAI22xp5_ASAP7_75t_SL g135 ( .A1(n_136), .A2(n_442), .B1(n_443), .B2(n_725), .Y(n_135) );
INVx2_ASAP7_75t_L g730 ( .A(n_136), .Y(n_730) );
XOR2xp5_ASAP7_75t_L g736 ( .A(n_136), .B(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_376), .Y(n_136) );
NAND5xp2_ASAP7_75t_L g137 ( .A(n_138), .B(n_305), .C(n_335), .D(n_356), .E(n_362), .Y(n_137) );
AOI221xp5_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_235), .B1(n_269), .B2(n_271), .C(n_282), .Y(n_138) );
INVxp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_232), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_204), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_SL g356 ( .A1(n_143), .A2(n_220), .B(n_357), .C(n_360), .Y(n_356) );
AND2x2_ASAP7_75t_L g426 ( .A(n_143), .B(n_221), .Y(n_426) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_182), .Y(n_143) );
AND2x2_ASAP7_75t_L g284 ( .A(n_144), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g288 ( .A(n_144), .B(n_285), .Y(n_288) );
OR2x2_ASAP7_75t_L g314 ( .A(n_144), .B(n_221), .Y(n_314) );
AND2x2_ASAP7_75t_L g316 ( .A(n_144), .B(n_207), .Y(n_316) );
AND2x2_ASAP7_75t_L g334 ( .A(n_144), .B(n_206), .Y(n_334) );
INVx1_ASAP7_75t_L g367 ( .A(n_144), .Y(n_367) );
INVx2_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
BUFx2_ASAP7_75t_L g234 ( .A(n_145), .Y(n_234) );
AND2x2_ASAP7_75t_L g270 ( .A(n_145), .B(n_207), .Y(n_270) );
AND2x2_ASAP7_75t_L g423 ( .A(n_145), .B(n_221), .Y(n_423) );
AO21x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_153), .B(n_178), .Y(n_145) );
INVx3_ASAP7_75t_L g219 ( .A(n_146), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_146), .B(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_146), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_SL g504 ( .A(n_146), .B(n_505), .Y(n_504) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_147), .Y(n_208) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_147), .A2(n_452), .B(n_459), .Y(n_451) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
AND2x2_ASAP7_75t_SL g181 ( .A(n_149), .B(n_150), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
OAI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_162), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_155), .A2(n_181), .B(n_223), .C(n_224), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_155), .A2(n_241), .B(n_242), .Y(n_240) );
OAI22xp33_ASAP7_75t_L g464 ( .A1(n_155), .A2(n_177), .B1(n_465), .B2(n_469), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_155), .A2(n_487), .B(n_488), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_155), .A2(n_531), .B(n_532), .Y(n_530) );
NAND2x1p5_ASAP7_75t_L g155 ( .A(n_156), .B(n_160), .Y(n_155) );
AND2x4_ASAP7_75t_L g189 ( .A(n_156), .B(n_160), .Y(n_189) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_159), .Y(n_156) );
INVx1_ASAP7_75t_L g200 ( .A(n_157), .Y(n_200) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
INVx1_ASAP7_75t_L g267 ( .A(n_158), .Y(n_267) );
INVx1_ASAP7_75t_L g165 ( .A(n_159), .Y(n_165) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_159), .Y(n_170) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_159), .Y(n_172) );
INVx3_ASAP7_75t_L g197 ( .A(n_159), .Y(n_197) );
INVx1_ASAP7_75t_L g456 ( .A(n_159), .Y(n_456) );
INVx4_ASAP7_75t_SL g177 ( .A(n_160), .Y(n_177) );
BUFx3_ASAP7_75t_L g229 ( .A(n_160), .Y(n_229) );
INVx5_ASAP7_75t_L g192 ( .A(n_163), .Y(n_192) );
AND2x6_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
BUFx3_ASAP7_75t_L g175 ( .A(n_164), .Y(n_175) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_164), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_171), .C(n_173), .Y(n_166) );
O2A1O1Ixp5_ASAP7_75t_L g243 ( .A1(n_168), .A2(n_173), .B(n_244), .C(n_245), .Y(n_243) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OAI22xp5_ASAP7_75t_SL g466 ( .A1(n_169), .A2(n_170), .B1(n_467), .B2(n_468), .Y(n_466) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx4_ASAP7_75t_L g199 ( .A(n_170), .Y(n_199) );
INVx4_ASAP7_75t_L g213 ( .A(n_172), .Y(n_213) );
INVx2_ASAP7_75t_L g254 ( .A(n_172), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_173), .A2(n_502), .B(n_503), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_173), .A2(n_534), .B(n_535), .Y(n_533) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g280 ( .A(n_175), .Y(n_280) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_SL g190 ( .A1(n_177), .A2(n_191), .B(n_192), .C(n_193), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_177), .A2(n_192), .B(n_211), .C(n_212), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_SL g251 ( .A1(n_177), .A2(n_192), .B(n_252), .C(n_253), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_SL g261 ( .A1(n_177), .A2(n_192), .B(n_262), .C(n_263), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_SL g275 ( .A1(n_177), .A2(n_192), .B(n_276), .C(n_277), .Y(n_275) );
O2A1O1Ixp33_ASAP7_75t_L g453 ( .A1(n_177), .A2(n_192), .B(n_454), .C(n_455), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g474 ( .A1(n_177), .A2(n_192), .B(n_475), .C(n_476), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_177), .A2(n_192), .B(n_522), .C(n_523), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
INVx1_ASAP7_75t_L g203 ( .A(n_180), .Y(n_203) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_180), .A2(n_509), .B(n_516), .Y(n_508) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g239 ( .A(n_181), .Y(n_239) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_181), .A2(n_250), .B(n_257), .Y(n_249) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_181), .A2(n_520), .B(n_526), .Y(n_519) );
AND2x2_ASAP7_75t_L g304 ( .A(n_182), .B(n_205), .Y(n_304) );
OR2x2_ASAP7_75t_L g308 ( .A(n_182), .B(n_221), .Y(n_308) );
AND2x2_ASAP7_75t_L g333 ( .A(n_182), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g380 ( .A(n_182), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_182), .B(n_342), .Y(n_428) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_186), .B(n_201), .Y(n_182) );
INVx1_ASAP7_75t_L g286 ( .A(n_183), .Y(n_286) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_183), .A2(n_530), .B(n_536), .Y(n_529) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AOI21xp5_ASAP7_75t_SL g498 ( .A1(n_184), .A2(n_499), .B(n_500), .Y(n_498) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AO21x2_ASAP7_75t_L g463 ( .A1(n_185), .A2(n_464), .B(n_470), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_185), .B(n_471), .Y(n_470) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_185), .A2(n_486), .B(n_493), .Y(n_485) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_187), .A2(n_202), .B(n_286), .Y(n_285) );
BUFx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_194), .B(n_200), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B1(n_198), .B2(n_199), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_196), .A2(n_226), .B(n_227), .C(n_228), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_196), .A2(n_490), .B(n_491), .C(n_492), .Y(n_489) );
INVx5_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_197), .B(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_197), .B(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_197), .B(n_478), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_199), .B(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_199), .B(n_279), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_199), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g228 ( .A(n_200), .Y(n_228) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
OAI322xp33_ASAP7_75t_L g429 ( .A1(n_204), .A2(n_365), .A3(n_388), .B1(n_409), .B2(n_430), .C1(n_432), .C2(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_205), .B(n_285), .Y(n_432) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_220), .Y(n_205) );
AND2x2_ASAP7_75t_L g233 ( .A(n_206), .B(n_234), .Y(n_233) );
AND2x4_ASAP7_75t_L g301 ( .A(n_206), .B(n_221), .Y(n_301) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g342 ( .A(n_207), .B(n_221), .Y(n_342) );
AND2x2_ASAP7_75t_L g386 ( .A(n_207), .B(n_220), .Y(n_386) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_218), .Y(n_207) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_208), .A2(n_260), .B(n_268), .Y(n_259) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_208), .A2(n_274), .B(n_281), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_213), .B(n_215), .Y(n_214) );
INVx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_217), .Y(n_514) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_219), .A2(n_473), .B(n_479), .Y(n_472) );
AND2x2_ASAP7_75t_L g269 ( .A(n_220), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g287 ( .A(n_220), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_220), .B(n_316), .Y(n_440) );
INVx3_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g232 ( .A(n_221), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_221), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g354 ( .A(n_221), .B(n_285), .Y(n_354) );
AND2x2_ASAP7_75t_L g381 ( .A(n_221), .B(n_316), .Y(n_381) );
OR2x2_ASAP7_75t_L g437 ( .A(n_221), .B(n_288), .Y(n_437) );
OR2x6_ASAP7_75t_L g221 ( .A(n_222), .B(n_230), .Y(n_221) );
INVx1_ASAP7_75t_SL g323 ( .A(n_232), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_233), .B(n_354), .Y(n_355) );
AND2x2_ASAP7_75t_L g389 ( .A(n_233), .B(n_379), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_233), .B(n_312), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_233), .B(n_434), .Y(n_433) );
OAI31xp33_ASAP7_75t_L g407 ( .A1(n_235), .A2(n_269), .A3(n_408), .B(n_410), .Y(n_407) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_248), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_236), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g390 ( .A(n_236), .B(n_325), .Y(n_390) );
OR2x2_ASAP7_75t_L g397 ( .A(n_236), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g409 ( .A(n_236), .B(n_298), .Y(n_409) );
CKINVDCx16_ASAP7_75t_R g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g343 ( .A(n_237), .B(n_344), .Y(n_343) );
BUFx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g271 ( .A(n_238), .B(n_272), .Y(n_271) );
INVx4_ASAP7_75t_L g292 ( .A(n_238), .Y(n_292) );
AND2x2_ASAP7_75t_L g329 ( .A(n_238), .B(n_273), .Y(n_329) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_246), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_239), .B(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_239), .B(n_517), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_239), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g328 ( .A(n_248), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g398 ( .A(n_248), .Y(n_398) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_258), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_249), .B(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g298 ( .A(n_249), .B(n_259), .Y(n_298) );
INVx2_ASAP7_75t_L g318 ( .A(n_249), .Y(n_318) );
AND2x2_ASAP7_75t_L g332 ( .A(n_249), .B(n_259), .Y(n_332) );
AND2x2_ASAP7_75t_L g339 ( .A(n_249), .B(n_295), .Y(n_339) );
BUFx3_ASAP7_75t_L g349 ( .A(n_249), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_249), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g294 ( .A(n_258), .Y(n_294) );
AND2x2_ASAP7_75t_L g302 ( .A(n_258), .B(n_292), .Y(n_302) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g272 ( .A(n_259), .B(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_259), .Y(n_326) );
INVx2_ASAP7_75t_L g492 ( .A(n_266), .Y(n_492) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_SL g309 ( .A(n_270), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_270), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_270), .B(n_379), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_271), .B(n_349), .Y(n_402) );
INVx1_ASAP7_75t_SL g436 ( .A(n_271), .Y(n_436) );
INVx1_ASAP7_75t_SL g344 ( .A(n_272), .Y(n_344) );
INVx1_ASAP7_75t_SL g295 ( .A(n_273), .Y(n_295) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_273), .Y(n_306) );
OR2x2_ASAP7_75t_L g317 ( .A(n_273), .B(n_292), .Y(n_317) );
AND2x2_ASAP7_75t_L g331 ( .A(n_273), .B(n_292), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_273), .B(n_321), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_287), .B(n_289), .C(n_300), .Y(n_282) );
AOI31xp33_ASAP7_75t_L g399 ( .A1(n_283), .A2(n_400), .A3(n_401), .B(n_402), .Y(n_399) );
AND2x2_ASAP7_75t_L g372 ( .A(n_284), .B(n_301), .Y(n_372) );
BUFx3_ASAP7_75t_L g312 ( .A(n_285), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_285), .B(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g348 ( .A(n_285), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_285), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g303 ( .A(n_288), .Y(n_303) );
OAI222xp33_ASAP7_75t_L g412 ( .A1(n_288), .A2(n_413), .B1(n_416), .B2(n_417), .C1(n_418), .C2(n_419), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_296), .Y(n_289) );
INVx1_ASAP7_75t_L g418 ( .A(n_290), .Y(n_418) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_292), .B(n_295), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_292), .B(n_318), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_292), .B(n_293), .Y(n_388) );
INVx1_ASAP7_75t_L g439 ( .A(n_292), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_293), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g441 ( .A(n_293), .Y(n_441) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx2_ASAP7_75t_L g321 ( .A(n_294), .Y(n_321) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_295), .Y(n_364) );
AOI32xp33_ASAP7_75t_L g300 ( .A1(n_296), .A2(n_301), .A3(n_302), .B1(n_303), .B2(n_304), .Y(n_300) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_298), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g375 ( .A(n_298), .Y(n_375) );
OR2x2_ASAP7_75t_L g416 ( .A(n_298), .B(n_317), .Y(n_416) );
INVx1_ASAP7_75t_L g352 ( .A(n_299), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_301), .B(n_312), .Y(n_337) );
INVx3_ASAP7_75t_L g346 ( .A(n_301), .Y(n_346) );
AOI322xp5_ASAP7_75t_L g362 ( .A1(n_301), .A2(n_346), .A3(n_363), .B1(n_365), .B2(n_368), .C1(n_372), .C2(n_373), .Y(n_362) );
AND2x2_ASAP7_75t_L g338 ( .A(n_302), .B(n_339), .Y(n_338) );
INVxp67_ASAP7_75t_L g415 ( .A(n_302), .Y(n_415) );
A2O1A1O1Ixp25_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B(n_310), .C(n_318), .D(n_319), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_306), .B(n_349), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
OAI221xp5_ASAP7_75t_L g319 ( .A1(n_308), .A2(n_320), .B1(n_323), .B2(n_324), .C(n_327), .Y(n_319) );
INVx1_ASAP7_75t_SL g434 ( .A(n_308), .Y(n_434) );
AOI21xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_315), .B(n_317), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_312), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI221xp5_ASAP7_75t_SL g404 ( .A1(n_314), .A2(n_398), .B1(n_405), .B2(n_406), .C(n_407), .Y(n_404) );
OAI222xp33_ASAP7_75t_L g435 ( .A1(n_315), .A2(n_436), .B1(n_437), .B2(n_438), .C1(n_440), .C2(n_441), .Y(n_435) );
AND2x2_ASAP7_75t_L g393 ( .A(n_316), .B(n_379), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_316), .A2(n_331), .B(n_378), .Y(n_405) );
INVx1_ASAP7_75t_L g419 ( .A(n_316), .Y(n_419) );
INVx2_ASAP7_75t_SL g322 ( .A(n_317), .Y(n_322) );
AND2x2_ASAP7_75t_L g325 ( .A(n_318), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_SL g359 ( .A(n_321), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_321), .B(n_331), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_322), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_322), .B(n_332), .Y(n_361) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OAI21xp5_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_330), .B(n_333), .Y(n_327) );
INVx1_ASAP7_75t_SL g345 ( .A(n_329), .Y(n_345) );
AND2x2_ASAP7_75t_L g392 ( .A(n_329), .B(n_375), .Y(n_392) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
AND2x2_ASAP7_75t_L g431 ( .A(n_331), .B(n_349), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_332), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g417 ( .A(n_333), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_338), .B1(n_340), .B2(n_347), .C(n_350), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .B1(n_345), .B2(n_346), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OAI22xp33_ASAP7_75t_L g350 ( .A1(n_344), .A2(n_351), .B1(n_353), .B2(n_355), .Y(n_350) );
OR2x2_ASAP7_75t_L g421 ( .A(n_345), .B(n_349), .Y(n_421) );
OR2x2_ASAP7_75t_L g424 ( .A(n_345), .B(n_359), .Y(n_424) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_366), .A2(n_421), .B1(n_422), .B2(n_424), .C(n_425), .Y(n_420) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND3xp33_ASAP7_75t_SL g376 ( .A(n_377), .B(n_391), .C(n_403), .Y(n_376) );
AOI222xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_382), .B1(n_384), .B2(n_387), .C1(n_389), .C2(n_390), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_379), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g401 ( .A(n_381), .Y(n_401) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B1(n_394), .B2(n_396), .C(n_399), .Y(n_391) );
INVx1_ASAP7_75t_L g406 ( .A(n_392), .Y(n_406) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OAI21xp33_ASAP7_75t_L g425 ( .A1(n_396), .A2(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
NOR5xp2_ASAP7_75t_L g403 ( .A(n_404), .B(n_412), .C(n_420), .D(n_429), .E(n_435), .Y(n_403) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVxp67_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_442), .A2(n_444), .B1(n_725), .B2(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_SL g444 ( .A(n_445), .B(n_662), .Y(n_444) );
NOR4xp25_ASAP7_75t_L g445 ( .A(n_446), .B(n_592), .C(n_623), .D(n_642), .Y(n_445) );
NAND4xp25_ASAP7_75t_L g446 ( .A(n_447), .B(n_550), .C(n_565), .D(n_583), .Y(n_446) );
AOI222xp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_495), .B1(n_527), .B2(n_538), .C1(n_543), .C2(n_545), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_480), .Y(n_448) );
INVx1_ASAP7_75t_L g606 ( .A(n_449), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_460), .Y(n_449) );
AND2x2_ASAP7_75t_L g481 ( .A(n_450), .B(n_472), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_450), .B(n_484), .Y(n_635) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g542 ( .A(n_451), .B(n_462), .Y(n_542) );
AND2x2_ASAP7_75t_L g551 ( .A(n_451), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g577 ( .A(n_451), .Y(n_577) );
AND2x2_ASAP7_75t_L g598 ( .A(n_451), .B(n_462), .Y(n_598) );
BUFx2_ASAP7_75t_L g621 ( .A(n_451), .Y(n_621) );
AND2x2_ASAP7_75t_L g645 ( .A(n_451), .B(n_463), .Y(n_645) );
AND2x2_ASAP7_75t_L g709 ( .A(n_451), .B(n_472), .Y(n_709) );
AND2x2_ASAP7_75t_L g610 ( .A(n_460), .B(n_541), .Y(n_610) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_461), .B(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_472), .Y(n_461) );
OR2x2_ASAP7_75t_L g570 ( .A(n_462), .B(n_485), .Y(n_570) );
AND2x2_ASAP7_75t_L g582 ( .A(n_462), .B(n_541), .Y(n_582) );
BUFx2_ASAP7_75t_L g714 ( .A(n_462), .Y(n_714) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g483 ( .A(n_463), .B(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g564 ( .A(n_463), .B(n_485), .Y(n_564) );
AND2x2_ASAP7_75t_L g617 ( .A(n_463), .B(n_472), .Y(n_617) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_463), .Y(n_653) );
AND2x2_ASAP7_75t_L g540 ( .A(n_472), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_SL g552 ( .A(n_472), .Y(n_552) );
INVx2_ASAP7_75t_L g563 ( .A(n_472), .Y(n_563) );
BUFx2_ASAP7_75t_L g587 ( .A(n_472), .Y(n_587) );
AND2x2_ASAP7_75t_SL g644 ( .A(n_472), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
AOI332xp33_ASAP7_75t_L g565 ( .A1(n_481), .A2(n_566), .A3(n_570), .B1(n_571), .B2(n_575), .B3(n_578), .C1(n_579), .C2(n_581), .Y(n_565) );
NAND2x1_ASAP7_75t_L g650 ( .A(n_481), .B(n_541), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_481), .B(n_555), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_SL g583 ( .A1(n_482), .A2(n_584), .B(n_587), .C(n_588), .Y(n_583) );
AND2x2_ASAP7_75t_L g722 ( .A(n_482), .B(n_563), .Y(n_722) );
INVx3_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g619 ( .A(n_483), .B(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g624 ( .A(n_483), .B(n_621), .Y(n_624) );
INVx1_ASAP7_75t_L g555 ( .A(n_484), .Y(n_555) );
AND2x2_ASAP7_75t_L g658 ( .A(n_484), .B(n_617), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_484), .B(n_598), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_484), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_484), .B(n_576), .Y(n_684) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx3_ASAP7_75t_L g541 ( .A(n_485), .Y(n_541) );
OAI31xp33_ASAP7_75t_L g723 ( .A1(n_495), .A2(n_644), .A3(n_651), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_506), .Y(n_495) );
AND2x2_ASAP7_75t_L g527 ( .A(n_496), .B(n_528), .Y(n_527) );
NAND2x1_ASAP7_75t_SL g546 ( .A(n_496), .B(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_496), .Y(n_633) );
AND2x2_ASAP7_75t_L g638 ( .A(n_496), .B(n_549), .Y(n_638) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_497), .A2(n_551), .B(n_553), .C(n_556), .Y(n_550) );
OR2x2_ASAP7_75t_L g567 ( .A(n_497), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g580 ( .A(n_497), .Y(n_580) );
AND2x2_ASAP7_75t_L g586 ( .A(n_497), .B(n_529), .Y(n_586) );
INVx2_ASAP7_75t_L g604 ( .A(n_497), .Y(n_604) );
AND2x2_ASAP7_75t_L g615 ( .A(n_497), .B(n_569), .Y(n_615) );
AND2x2_ASAP7_75t_L g647 ( .A(n_497), .B(n_605), .Y(n_647) );
AND2x2_ASAP7_75t_L g651 ( .A(n_497), .B(n_574), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_497), .B(n_506), .Y(n_656) );
AND2x2_ASAP7_75t_L g690 ( .A(n_497), .B(n_691), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_497), .B(n_593), .Y(n_724) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_504), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_506), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g632 ( .A(n_506), .Y(n_632) );
AND2x2_ASAP7_75t_L g694 ( .A(n_506), .B(n_615), .Y(n_694) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
OR2x2_ASAP7_75t_L g548 ( .A(n_507), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g558 ( .A(n_507), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_507), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g666 ( .A(n_507), .Y(n_666) );
AND2x2_ASAP7_75t_L g683 ( .A(n_507), .B(n_529), .Y(n_683) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g574 ( .A(n_508), .B(n_518), .Y(n_574) );
AND2x2_ASAP7_75t_L g603 ( .A(n_508), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g614 ( .A(n_508), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_508), .B(n_569), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_515), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_514), .Y(n_511) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g528 ( .A(n_519), .B(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g549 ( .A(n_519), .Y(n_549) );
AND2x2_ASAP7_75t_L g605 ( .A(n_519), .B(n_569), .Y(n_605) );
INVx1_ASAP7_75t_L g707 ( .A(n_527), .Y(n_707) );
INVx1_ASAP7_75t_L g711 ( .A(n_528), .Y(n_711) );
INVx2_ASAP7_75t_L g569 ( .A(n_529), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_542), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_540), .B(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_540), .B(n_645), .Y(n_703) );
OR2x2_ASAP7_75t_L g544 ( .A(n_541), .B(n_542), .Y(n_544) );
INVx1_ASAP7_75t_SL g596 ( .A(n_541), .Y(n_596) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_547), .A2(n_600), .B1(n_602), .B2(n_606), .C(n_607), .Y(n_599) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g627 ( .A(n_548), .B(n_591), .Y(n_627) );
INVx2_ASAP7_75t_L g559 ( .A(n_549), .Y(n_559) );
INVx1_ASAP7_75t_L g585 ( .A(n_549), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_549), .B(n_569), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_549), .B(n_572), .Y(n_679) );
INVx1_ASAP7_75t_L g687 ( .A(n_549), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_551), .B(n_555), .Y(n_601) );
AND2x4_ASAP7_75t_L g576 ( .A(n_552), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g689 ( .A(n_555), .B(n_645), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_557), .B(n_560), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_558), .B(n_590), .Y(n_589) );
INVxp67_ASAP7_75t_L g697 ( .A(n_559), .Y(n_697) );
INVxp67_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g597 ( .A(n_563), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g669 ( .A(n_563), .B(n_645), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_563), .B(n_582), .Y(n_675) );
AOI322xp5_ASAP7_75t_L g629 ( .A1(n_564), .A2(n_598), .A3(n_605), .B1(n_630), .B2(n_633), .C1(n_634), .C2(n_636), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_564), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g695 ( .A(n_567), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g641 ( .A(n_568), .Y(n_641) );
INVx2_ASAP7_75t_L g572 ( .A(n_569), .Y(n_572) );
INVx1_ASAP7_75t_L g631 ( .A(n_569), .Y(n_631) );
CKINVDCx16_ASAP7_75t_R g578 ( .A(n_570), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
AND2x2_ASAP7_75t_L g667 ( .A(n_572), .B(n_580), .Y(n_667) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g579 ( .A(n_574), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g622 ( .A(n_574), .B(n_615), .Y(n_622) );
AND2x2_ASAP7_75t_L g626 ( .A(n_574), .B(n_586), .Y(n_626) );
OAI21xp33_ASAP7_75t_SL g636 ( .A1(n_575), .A2(n_637), .B(n_639), .Y(n_636) );
OAI22xp33_ASAP7_75t_L g706 ( .A1(n_575), .A2(n_707), .B1(n_708), .B2(n_710), .Y(n_706) );
INVx3_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g581 ( .A(n_576), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_576), .B(n_596), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_578), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g718 ( .A(n_585), .Y(n_718) );
INVx4_ASAP7_75t_L g591 ( .A(n_586), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_586), .B(n_613), .Y(n_661) );
INVx1_ASAP7_75t_SL g673 ( .A(n_587), .Y(n_673) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp67_ASAP7_75t_L g686 ( .A(n_591), .B(n_687), .Y(n_686) );
OAI211xp5_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_594), .B(n_599), .C(n_616), .Y(n_592) );
OAI221xp5_ASAP7_75t_SL g712 ( .A1(n_594), .A2(n_632), .B1(n_711), .B2(n_713), .C(n_715), .Y(n_712) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_596), .B(n_709), .Y(n_708) );
OAI31xp33_ASAP7_75t_L g688 ( .A1(n_597), .A2(n_674), .A3(n_689), .B(n_690), .Y(n_688) );
INVx1_ASAP7_75t_L g628 ( .A(n_598), .Y(n_628) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g678 ( .A(n_603), .Y(n_678) );
AND2x2_ASAP7_75t_L g691 ( .A(n_605), .B(n_614), .Y(n_691) );
AOI21xp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B(n_611), .Y(n_607) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
INVxp67_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_615), .B(n_718), .Y(n_717) );
OAI21xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B(n_622), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OAI221xp5_ASAP7_75t_SL g623 ( .A1(n_624), .A2(n_625), .B1(n_627), .B2(n_628), .C(n_629), .Y(n_623) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_624), .A2(n_693), .B(n_695), .C(n_698), .Y(n_692) );
CKINVDCx16_ASAP7_75t_R g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_627), .B(n_677), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx1_ASAP7_75t_L g654 ( .A(n_635), .Y(n_654) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g640 ( .A(n_638), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g682 ( .A(n_638), .B(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI211xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B(n_648), .C(n_657), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g719 ( .A1(n_646), .A2(n_656), .B1(n_720), .B2(n_721), .C(n_723), .Y(n_719) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_651), .B1(n_652), .B2(n_655), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI21xp5_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_659), .B(n_660), .Y(n_657) );
INVx1_ASAP7_75t_SL g720 ( .A(n_659), .Y(n_720) );
INVxp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NOR4xp25_ASAP7_75t_L g662 ( .A(n_663), .B(n_692), .C(n_712), .D(n_719), .Y(n_662) );
OAI211xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_668), .B(n_670), .C(n_688), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
O2A1O1Ixp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_674), .B(n_676), .C(n_680), .Y(n_670) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g699 ( .A(n_677), .Y(n_699) );
OR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
OR2x2_ASAP7_75t_L g710 ( .A(n_678), .B(n_711), .Y(n_710) );
OAI21xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_684), .B(n_685), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B1(n_702), .B2(n_704), .C(n_706), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVxp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_709), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_738), .Y(n_742) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
endmodule