module fake_jpeg_30698_n_458 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_458);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_458;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_14),
.B(n_13),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_6),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_49),
.A2(n_45),
.B1(n_48),
.B2(n_38),
.Y(n_123)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_16),
.B(n_6),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_20),
.Y(n_110)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_32),
.B(n_6),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_67),
.B(n_91),
.Y(n_124)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_69),
.Y(n_137)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_33),
.B(n_20),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_90),
.Y(n_100)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_80),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_25),
.Y(n_87)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_89),
.A2(n_94),
.B1(n_45),
.B2(n_34),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_16),
.B(n_8),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

BUFx24_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_92),
.Y(n_149)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_93),
.B(n_27),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_58),
.A2(n_63),
.B1(n_76),
.B2(n_56),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_108),
.A2(n_123),
.B1(n_136),
.B2(n_69),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_110),
.B(n_21),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_53),
.A2(n_47),
.B1(n_48),
.B2(n_44),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_111),
.A2(n_140),
.B1(n_143),
.B2(n_89),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_59),
.A2(n_45),
.B1(n_34),
.B2(n_24),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_114),
.A2(n_27),
.B1(n_21),
.B2(n_37),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_119),
.A2(n_82),
.B1(n_81),
.B2(n_57),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_60),
.B(n_47),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_126),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_44),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_130),
.B(n_37),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_L g136 ( 
.A1(n_62),
.A2(n_42),
.B1(n_46),
.B2(n_26),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_54),
.B(n_43),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_144),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_65),
.A2(n_43),
.B1(n_39),
.B2(n_38),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_87),
.A2(n_24),
.B1(n_34),
.B2(n_42),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_54),
.B(n_39),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_95),
.B(n_26),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_28),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_153),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_154),
.A2(n_176),
.B1(n_181),
.B2(n_192),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_105),
.B(n_64),
.C(n_70),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_155),
.B(n_146),
.C(n_135),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_156),
.A2(n_167),
.B1(n_172),
.B2(n_178),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g216 ( 
.A1(n_157),
.A2(n_196),
.B1(n_101),
.B2(n_104),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_158),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

INVx3_ASAP7_75t_SL g202 ( 
.A(n_159),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_117),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_168),
.Y(n_203)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_161),
.Y(n_233)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_162),
.Y(n_232)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_127),
.A2(n_94),
.B1(n_74),
.B2(n_79),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_165),
.Y(n_236)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

INVx4_ASAP7_75t_SL g168 ( 
.A(n_104),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_173),
.Y(n_204)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_170),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_124),
.A2(n_72),
.B1(n_85),
.B2(n_77),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_179),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_116),
.A2(n_34),
.B1(n_24),
.B2(n_73),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_116),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_182),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_102),
.A2(n_75),
.B1(n_92),
.B2(n_34),
.Y(n_178)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_112),
.A2(n_37),
.B1(n_27),
.B2(n_21),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_199),
.B1(n_114),
.B2(n_119),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_137),
.A2(n_37),
.B1(n_27),
.B2(n_21),
.Y(n_181)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_184),
.Y(n_229)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_186),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_137),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_107),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_187),
.Y(n_230)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_190),
.Y(n_225)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_97),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_189),
.B(n_195),
.Y(n_235)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_125),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_194),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_108),
.A2(n_92),
.B1(n_10),
.B2(n_12),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_197),
.B(n_101),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

AO22x2_ASAP7_75t_SL g196 ( 
.A1(n_136),
.A2(n_37),
.B1(n_27),
.B2(n_21),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_198),
.B(n_4),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_103),
.A2(n_28),
.B1(n_5),
.B2(n_8),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_118),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_220),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_206),
.A2(n_211),
.B1(n_216),
.B2(n_224),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_120),
.B(n_145),
.C(n_143),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_209),
.A2(n_214),
.B(n_193),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_157),
.A2(n_102),
.B1(n_131),
.B2(n_112),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_172),
.A2(n_131),
.B1(n_146),
.B2(n_135),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_213),
.A2(n_163),
.B1(n_191),
.B2(n_188),
.Y(n_264)
);

O2A1O1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_196),
.A2(n_147),
.B(n_149),
.C(n_106),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_110),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_L g270 ( 
.A1(n_221),
.A2(n_234),
.B(n_8),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_156),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_192),
.A2(n_103),
.B1(n_100),
.B2(n_142),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_155),
.A2(n_28),
.B1(n_1),
.B2(n_2),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_226),
.A2(n_208),
.B1(n_206),
.B2(n_200),
.Y(n_250)
);

AOI32xp33_ASAP7_75t_L g227 ( 
.A1(n_174),
.A2(n_28),
.A3(n_5),
.B1(n_8),
.B2(n_15),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_227),
.B(n_15),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_153),
.B(n_0),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_238),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_171),
.B(n_4),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_237),
.Y(n_239)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_239),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_228),
.B(n_166),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_240),
.B(n_254),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_210),
.B(n_195),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_243),
.B(n_247),
.Y(n_283)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_189),
.C(n_184),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_245),
.B(n_255),
.C(n_256),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_262),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_250),
.A2(n_265),
.B1(n_200),
.B2(n_213),
.Y(n_282)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_251),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_216),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_209),
.A2(n_220),
.B(n_205),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_253),
.A2(n_229),
.B(n_226),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_152),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_161),
.C(n_183),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_170),
.Y(n_256)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_238),
.B(n_165),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_260),
.Y(n_284)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_259),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_203),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_201),
.Y(n_261)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_261),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_212),
.B(n_190),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_162),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_263),
.B(n_271),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_264),
.A2(n_266),
.B1(n_202),
.B2(n_224),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_211),
.A2(n_179),
.B1(n_194),
.B2(n_173),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_216),
.A2(n_159),
.B1(n_185),
.B2(n_187),
.Y(n_266)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_217),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_267),
.A2(n_202),
.B1(n_257),
.B2(n_218),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_208),
.A2(n_168),
.B(n_175),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_268),
.A2(n_216),
.B(n_207),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_231),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_269),
.Y(n_297)
);

OAI21xp33_ASAP7_75t_L g300 ( 
.A1(n_270),
.A2(n_272),
.B(n_273),
.Y(n_300)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_229),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_L g273 ( 
.A1(n_234),
.A2(n_9),
.B(n_13),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_254),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_275),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_243),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_276),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_278),
.B(n_292),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_235),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_281),
.B(n_247),
.C(n_246),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_282),
.A2(n_288),
.B1(n_293),
.B2(n_302),
.Y(n_308)
);

AND2x2_ASAP7_75t_SL g285 ( 
.A(n_259),
.B(n_261),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_285),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_287),
.A2(n_268),
.B(n_266),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_248),
.A2(n_216),
.B1(n_209),
.B2(n_214),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_291),
.B(n_250),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_290),
.A2(n_303),
.B1(n_265),
.B2(n_251),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_252),
.A2(n_214),
.B1(n_202),
.B2(n_236),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_258),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_306),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_298),
.A2(n_241),
.B(n_240),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_248),
.A2(n_227),
.B1(n_204),
.B2(n_218),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_256),
.A2(n_204),
.B1(n_225),
.B2(n_218),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_263),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_307),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_309),
.B(n_312),
.C(n_333),
.Y(n_340)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_311),
.A2(n_316),
.B(n_332),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_241),
.C(n_262),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_317),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_276),
.B(n_242),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_326),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_299),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_320),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_289),
.A2(n_271),
.B(n_242),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_322),
.Y(n_352)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_299),
.Y(n_323)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_323),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_324),
.A2(n_330),
.B1(n_282),
.B2(n_275),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_283),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_325),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_279),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_327),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_288),
.A2(n_302),
.B1(n_293),
.B2(n_289),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_328),
.A2(n_329),
.B1(n_303),
.B2(n_306),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_289),
.A2(n_264),
.B1(n_249),
.B2(n_267),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_290),
.A2(n_244),
.B1(n_239),
.B2(n_267),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_283),
.A2(n_236),
.B(n_222),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_331),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_284),
.A2(n_222),
.B(n_233),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_274),
.B(n_230),
.C(n_233),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_298),
.A2(n_215),
.B(n_230),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g344 ( 
.A(n_334),
.B(n_280),
.CI(n_305),
.CON(n_344),
.SN(n_344)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_274),
.B(n_232),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_286),
.C(n_297),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_307),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_336),
.B(n_344),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_338),
.A2(n_348),
.B1(n_349),
.B2(n_354),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_341),
.A2(n_345),
.B1(n_310),
.B2(n_326),
.Y(n_384)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_342),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_324),
.A2(n_311),
.B1(n_330),
.B2(n_325),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_346),
.B(n_357),
.C(n_318),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_286),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_322),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_308),
.A2(n_304),
.B1(n_301),
.B2(n_305),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_308),
.A2(n_304),
.B1(n_301),
.B2(n_285),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_328),
.A2(n_285),
.B1(n_291),
.B2(n_297),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_309),
.B(n_285),
.C(n_280),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_329),
.A2(n_284),
.B1(n_295),
.B2(n_300),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_358),
.A2(n_354),
.B1(n_349),
.B2(n_338),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_319),
.B(n_295),
.Y(n_360)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_360),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_360),
.Y(n_364)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_364),
.Y(n_392)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_337),
.Y(n_365)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_365),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_340),
.B(n_335),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_370),
.Y(n_391)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_367),
.Y(n_399)
);

XOR2x2_ASAP7_75t_L g368 ( 
.A(n_347),
.B(n_316),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_368),
.B(n_382),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_357),
.B(n_333),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_369),
.B(n_373),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_346),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_348),
.A2(n_313),
.B1(n_314),
.B2(n_321),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_377),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_358),
.B(n_313),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_375),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_376),
.B(n_378),
.C(n_380),
.Y(n_389)
);

AO21x1_ASAP7_75t_L g377 ( 
.A1(n_339),
.A2(n_334),
.B(n_315),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_342),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_350),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_352),
.B(n_344),
.C(n_339),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_350),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_381),
.B(n_383),
.Y(n_390)
);

OAI21xp33_ASAP7_75t_L g382 ( 
.A1(n_352),
.A2(n_315),
.B(n_314),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_SL g383 ( 
.A(n_356),
.B(n_331),
.Y(n_383)
);

XNOR2x1_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_345),
.Y(n_398)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_363),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_385),
.B(n_394),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_359),
.C(n_353),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_393),
.B(n_402),
.C(n_368),
.Y(n_408)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_362),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_395),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_398),
.B(n_373),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_372),
.B(n_359),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_400),
.Y(n_414)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_380),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_401),
.B(n_369),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_353),
.C(n_344),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_408),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_396),
.A2(n_371),
.B1(n_341),
.B2(n_374),
.Y(n_404)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_404),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_387),
.A2(n_371),
.B1(n_336),
.B2(n_355),
.Y(n_405)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_405),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_407),
.B(n_323),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_391),
.B(n_378),
.C(n_376),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_412),
.C(n_413),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_389),
.B(n_377),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_398),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_332),
.C(n_361),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_389),
.B(n_401),
.C(n_388),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_388),
.B(n_393),
.C(n_402),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_386),
.C(n_351),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_392),
.A2(n_382),
.B1(n_361),
.B2(n_355),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_416),
.A2(n_387),
.B1(n_385),
.B2(n_399),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_423),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_420),
.B(n_424),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_414),
.A2(n_397),
.B1(n_390),
.B2(n_400),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_421),
.A2(n_426),
.B1(n_425),
.B2(n_406),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_413),
.A2(n_395),
.B(n_386),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_422),
.B(n_277),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_343),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_403),
.A2(n_343),
.B1(n_327),
.B2(n_320),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_426),
.B(n_416),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_427),
.B(n_429),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_408),
.B(n_317),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_430),
.B(n_420),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_428),
.A2(n_411),
.B(n_415),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_431),
.A2(n_433),
.B(n_424),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_419),
.A2(n_409),
.B(n_412),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_434),
.B(n_435),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_421),
.A2(n_277),
.B1(n_215),
.B2(n_232),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_438),
.B(n_9),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_9),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_439),
.B(n_423),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_431),
.B(n_417),
.C(n_429),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_440),
.A2(n_444),
.B(n_430),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_442),
.B(n_445),
.Y(n_449)
);

NOR2x1_ASAP7_75t_SL g443 ( 
.A(n_432),
.B(n_417),
.Y(n_443)
);

O2A1O1Ixp33_ASAP7_75t_SL g447 ( 
.A1(n_443),
.A2(n_436),
.B(n_437),
.C(n_434),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_446),
.B(n_15),
.C(n_1),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_447),
.A2(n_450),
.B(n_441),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g453 ( 
.A(n_448),
.Y(n_453)
);

AO21x1_ASAP7_75t_L g451 ( 
.A1(n_449),
.A2(n_441),
.B(n_15),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_451),
.A2(n_452),
.B(n_0),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_454),
.A2(n_453),
.B(n_2),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_455),
.A2(n_2),
.B(n_3),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_456),
.A2(n_3),
.B(n_360),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_457),
.B(n_3),
.Y(n_458)
);


endmodule