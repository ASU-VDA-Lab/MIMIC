module fake_jpeg_13795_n_36 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_36);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_15;

INVx8_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_1),
.Y(n_24)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

AO22x1_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_20),
.B1(n_12),
.B2(n_16),
.Y(n_25)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_24),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_16),
.B(n_2),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_2),
.B(n_3),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_25),
.B(n_16),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_29),
.B(n_21),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_12),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_31),
.B(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_3),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_4),
.Y(n_35)
);

OAI321xp33_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_4),
.A3(n_34),
.B1(n_7),
.B2(n_10),
.C(n_11),
.Y(n_36)
);


endmodule