module fake_ariane_2906_n_1743 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1743);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1743;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_45),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_104),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_118),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_1),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_70),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_32),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_80),
.Y(n_164)
);

BUFx10_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_93),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_41),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_61),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_29),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_1),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_0),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_78),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_153),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_13),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_33),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_154),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_101),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_60),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_65),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_47),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_71),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_63),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_46),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_132),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_19),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_119),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_15),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_143),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_46),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_149),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_98),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_39),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_145),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_112),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_82),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_140),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_95),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_107),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_117),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_30),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_3),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_113),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_56),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_66),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_16),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_124),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_67),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_131),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_69),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_0),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_57),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_111),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_18),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_47),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_6),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_23),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_94),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_36),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_33),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_52),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_136),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_5),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_36),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_125),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_97),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_21),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_83),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_8),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_73),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_28),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_144),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_152),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_27),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_12),
.Y(n_240)
);

HB1xp67_ASAP7_75t_SL g241 ( 
.A(n_9),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_59),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_29),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_100),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_103),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_2),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_72),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_4),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_32),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_115),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_15),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_128),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_114),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_39),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_19),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_88),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_30),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_34),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_109),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_3),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_7),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_133),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_22),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_50),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_38),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_51),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_42),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_146),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_123),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_81),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_77),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_9),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_55),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_10),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_99),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_35),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_21),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_17),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_17),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_54),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_2),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_148),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_85),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_89),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_91),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_41),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_38),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_129),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_74),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_4),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_96),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_64),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_34),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_68),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_11),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_137),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_108),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_35),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_23),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_130),
.Y(n_300)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_150),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_43),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_87),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_24),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_37),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_142),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_40),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_11),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_139),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_160),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_168),
.Y(n_311)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_170),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_194),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_203),
.Y(n_314)
);

INVxp33_ASAP7_75t_SL g315 ( 
.A(n_170),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_228),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_215),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_241),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_218),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_220),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_175),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_164),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_180),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_168),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_219),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_219),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_201),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_198),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_210),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_223),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_223),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_244),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_292),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_250),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_224),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_296),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_181),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_229),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_165),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_234),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_156),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_240),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_163),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_239),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_165),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_165),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_251),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_157),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_261),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_157),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_265),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_287),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_176),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_290),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_172),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_239),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_302),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_298),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_176),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_298),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_158),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_158),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_199),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_159),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_307),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_274),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_274),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_189),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_286),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_159),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_161),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_286),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_295),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_295),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_226),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_226),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_191),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_295),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_161),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_230),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_162),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_162),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_318),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_193),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_365),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_365),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_341),
.A2(n_305),
.B1(n_249),
.B2(n_175),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_365),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_337),
.A2(n_187),
.B1(n_185),
.B2(n_304),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_377),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_377),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_378),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_339),
.B(n_166),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_321),
.Y(n_396)
);

CKINVDCx8_ASAP7_75t_R g397 ( 
.A(n_323),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_378),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_322),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_L g400 ( 
.A(n_348),
.B(n_202),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_337),
.A2(n_278),
.B1(n_236),
.B2(n_304),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_360),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_365),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_365),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_382),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_328),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_177),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_312),
.A2(n_171),
.B1(n_182),
.B2(n_293),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_382),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_343),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_311),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_311),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_353),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_324),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_324),
.Y(n_415)
);

AND2x6_ASAP7_75t_L g416 ( 
.A(n_360),
.B(n_230),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_325),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_R g418 ( 
.A(n_380),
.B(n_190),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_325),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_339),
.B(n_166),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_315),
.A2(n_316),
.B1(n_327),
.B2(n_333),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_355),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_326),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_326),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_375),
.B(n_231),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_330),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_327),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_330),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_331),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_331),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_344),
.B(n_356),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_359),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_329),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_361),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_363),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_370),
.B(n_177),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_376),
.B(n_231),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_367),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_348),
.B(n_238),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_310),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_313),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_314),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_332),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_350),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_333),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_368),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_317),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_371),
.B(n_374),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_319),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_320),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_335),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_350),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_338),
.Y(n_453)
);

CKINVDCx11_ASAP7_75t_R g454 ( 
.A(n_410),
.Y(n_454)
);

NAND2xp33_ASAP7_75t_SL g455 ( 
.A(n_418),
.B(n_362),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_424),
.Y(n_456)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_404),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_392),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_345),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_385),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_424),
.Y(n_461)
);

AND2x6_ASAP7_75t_L g462 ( 
.A(n_407),
.B(n_242),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_424),
.Y(n_463)
);

AND2x6_ASAP7_75t_L g464 ( 
.A(n_407),
.B(n_242),
.Y(n_464)
);

AND2x6_ASAP7_75t_L g465 ( 
.A(n_393),
.B(n_280),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_444),
.B(n_362),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_444),
.B(n_364),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_408),
.A2(n_281),
.B1(n_187),
.B2(n_185),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_424),
.Y(n_469)
);

NAND3xp33_ASAP7_75t_L g470 ( 
.A(n_453),
.B(n_366),
.C(n_364),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_393),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_366),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_424),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_395),
.B(n_372),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_420),
.B(n_372),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_416),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_402),
.B(n_373),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_427),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_427),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_402),
.B(n_345),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_394),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_416),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_424),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_396),
.B(n_373),
.Y(n_484)
);

AND3x2_ASAP7_75t_L g485 ( 
.A(n_445),
.B(n_276),
.C(n_340),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_442),
.B(n_447),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_414),
.Y(n_487)
);

NOR2x1p5_ASAP7_75t_L g488 ( 
.A(n_440),
.B(n_346),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_402),
.B(n_346),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_414),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_425),
.A2(n_351),
.B1(n_342),
.B2(n_347),
.Y(n_491)
);

AO22x2_ASAP7_75t_L g492 ( 
.A1(n_391),
.A2(n_280),
.B1(n_291),
.B2(n_358),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_404),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_453),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_431),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_414),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_431),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_413),
.B(n_446),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_453),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_SL g501 ( 
.A1(n_389),
.A2(n_334),
.B1(n_336),
.B2(n_379),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_415),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_415),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_396),
.B(n_381),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_453),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_445),
.B(n_381),
.Y(n_506)
);

NAND3xp33_ASAP7_75t_L g507 ( 
.A(n_453),
.B(n_384),
.C(n_383),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_425),
.A2(n_352),
.B1(n_349),
.B2(n_357),
.Y(n_508)
);

INVx8_ASAP7_75t_L g509 ( 
.A(n_416),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_415),
.Y(n_510)
);

AND3x2_ASAP7_75t_L g511 ( 
.A(n_397),
.B(n_354),
.C(n_291),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_419),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_419),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_398),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_399),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_416),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_398),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_425),
.A2(n_384),
.B1(n_383),
.B2(n_285),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_404),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_419),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_453),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_426),
.Y(n_522)
);

AOI21x1_ASAP7_75t_L g523 ( 
.A1(n_386),
.A2(n_309),
.B(n_205),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_426),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_425),
.B(n_167),
.Y(n_525)
);

AOI21x1_ASAP7_75t_L g526 ( 
.A1(n_386),
.A2(n_222),
.B(n_303),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_404),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_422),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_405),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_405),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_413),
.B(n_167),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_426),
.Y(n_532)
);

AO22x2_ASAP7_75t_L g533 ( 
.A1(n_391),
.A2(n_297),
.B1(n_209),
.B2(n_213),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_442),
.B(n_236),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_428),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_413),
.B(n_446),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_409),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_413),
.B(n_169),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_404),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_437),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_446),
.B(n_169),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_428),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_437),
.B(n_277),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_409),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_406),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_428),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_404),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_437),
.A2(n_255),
.B1(n_232),
.B2(n_243),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_411),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_416),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_387),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_437),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_411),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_412),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_416),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_387),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_440),
.B(n_277),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_412),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_387),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_388),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_442),
.B(n_278),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_388),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_388),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_447),
.B(n_279),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_417),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_441),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_408),
.B(n_421),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_417),
.Y(n_568)
);

NOR3xp33_ASAP7_75t_L g569 ( 
.A(n_401),
.B(n_279),
.C(n_281),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_441),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_423),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_390),
.Y(n_572)
);

OR2x6_ASAP7_75t_L g573 ( 
.A(n_389),
.B(n_214),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_401),
.A2(n_254),
.B1(n_246),
.B2(n_248),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_450),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_390),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_450),
.B(n_173),
.Y(n_577)
);

INVx5_ASAP7_75t_L g578 ( 
.A(n_416),
.Y(n_578)
);

INVxp33_ASAP7_75t_L g579 ( 
.A(n_436),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_390),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_447),
.B(n_299),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_423),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_403),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_403),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_429),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_416),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_403),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_432),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_429),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_435),
.Y(n_590)
);

INVxp67_ASAP7_75t_SL g591 ( 
.A(n_451),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_400),
.B(n_225),
.Y(n_592)
);

OAI22xp33_ASAP7_75t_L g593 ( 
.A1(n_421),
.A2(n_299),
.B1(n_272),
.B2(n_267),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_432),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_433),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_430),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_451),
.B(n_235),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_430),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_448),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_449),
.B(n_256),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_432),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_435),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_478),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_566),
.A2(n_397),
.B1(n_208),
.B2(n_221),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_566),
.A2(n_397),
.B1(n_263),
.B2(n_260),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_478),
.B(n_443),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_496),
.B(n_449),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_459),
.B(n_449),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_590),
.B(n_173),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_496),
.B(n_435),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_498),
.B(n_435),
.Y(n_611)
);

NOR2xp67_ASAP7_75t_L g612 ( 
.A(n_479),
.B(n_434),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_460),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_590),
.B(n_174),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_498),
.B(n_434),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_575),
.B(n_438),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_575),
.B(n_438),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_591),
.B(n_448),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_590),
.B(n_174),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_474),
.B(n_257),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_588),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_484),
.B(n_436),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_458),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_590),
.B(n_178),
.Y(n_624)
);

INVx8_ASAP7_75t_L g625 ( 
.A(n_462),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_528),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_592),
.B(n_178),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_570),
.B(n_179),
.Y(n_628)
);

A2O1A1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_468),
.A2(n_282),
.B(n_300),
.C(n_289),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_460),
.B(n_258),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_590),
.B(n_179),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_588),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_475),
.B(n_183),
.Y(n_633)
);

AO221x1_ASAP7_75t_L g634 ( 
.A1(n_593),
.A2(n_199),
.B1(n_288),
.B2(n_7),
.C(n_8),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_462),
.A2(n_306),
.B1(n_184),
.B2(n_294),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_454),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_484),
.B(n_183),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_466),
.B(n_184),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_471),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_588),
.Y(n_640)
);

NOR2xp67_ASAP7_75t_L g641 ( 
.A(n_470),
.B(n_306),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_588),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_570),
.B(n_186),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_588),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_534),
.B(n_186),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_511),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_590),
.B(n_188),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_470),
.B(n_188),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_570),
.B(n_233),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_507),
.B(n_233),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_528),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_540),
.B(n_283),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_471),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_507),
.A2(n_283),
.B1(n_284),
.B2(n_294),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_481),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_543),
.B(n_284),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_476),
.B(n_301),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_467),
.B(n_477),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_480),
.B(n_5),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g660 ( 
.A(n_545),
.Y(n_660)
);

NOR2xp67_ASAP7_75t_L g661 ( 
.A(n_515),
.B(n_192),
.Y(n_661)
);

NAND2x1_ASAP7_75t_L g662 ( 
.A(n_476),
.B(n_199),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_481),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_495),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_540),
.B(n_195),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_489),
.B(n_6),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_487),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_552),
.B(n_196),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_552),
.B(n_197),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_L g670 ( 
.A(n_462),
.B(n_301),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_599),
.A2(n_273),
.B1(n_211),
.B2(n_207),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_495),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_534),
.B(n_252),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_462),
.A2(n_247),
.B1(n_275),
.B2(n_271),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_487),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_545),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_490),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_476),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_490),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_595),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_561),
.B(n_245),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_497),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_599),
.B(n_10),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_561),
.B(n_564),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_564),
.B(n_253),
.Y(n_685)
);

INVxp67_ASAP7_75t_SL g686 ( 
.A(n_500),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_504),
.B(n_12),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_506),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_514),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_514),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_476),
.B(n_301),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_509),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_581),
.B(n_237),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_509),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_497),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_581),
.B(n_259),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_462),
.B(n_227),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_517),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_499),
.A2(n_217),
.B(n_270),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_482),
.B(n_301),
.Y(n_700)
);

NOR2x1_ASAP7_75t_L g701 ( 
.A(n_488),
.B(n_199),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_472),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_462),
.B(n_262),
.Y(n_703)
);

BUFx2_ASAP7_75t_R g704 ( 
.A(n_567),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_557),
.B(n_13),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_502),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_502),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_462),
.B(n_216),
.Y(n_708)
);

BUFx12f_ASAP7_75t_L g709 ( 
.A(n_573),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_455),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_464),
.A2(n_212),
.B1(n_269),
.B2(n_268),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_464),
.B(n_266),
.Y(n_712)
);

NOR2xp67_ASAP7_75t_L g713 ( 
.A(n_468),
.B(n_200),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_503),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_464),
.B(n_264),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_557),
.B(n_14),
.Y(n_716)
);

OAI22xp33_ASAP7_75t_L g717 ( 
.A1(n_573),
.A2(n_204),
.B1(n_206),
.B2(n_199),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_517),
.Y(n_718)
);

INVx4_ASAP7_75t_L g719 ( 
.A(n_509),
.Y(n_719)
);

OAI22xp33_ASAP7_75t_L g720 ( 
.A1(n_573),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_482),
.B(n_516),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_529),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_488),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_557),
.B(n_20),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_464),
.B(n_301),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_574),
.B(n_20),
.C(n_22),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_557),
.B(n_24),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_482),
.B(n_301),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_464),
.B(n_301),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_525),
.B(n_25),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_509),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_503),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_482),
.B(n_516),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_464),
.B(n_301),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_516),
.B(n_25),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_509),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_464),
.B(n_26),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_529),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_485),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_510),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_602),
.B(n_26),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_500),
.Y(n_742)
);

BUFx8_ASAP7_75t_L g743 ( 
.A(n_543),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_516),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_541),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_530),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_510),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_550),
.B(n_27),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_550),
.B(n_28),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_512),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_486),
.B(n_31),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_602),
.B(n_31),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_543),
.B(n_37),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_530),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_537),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_537),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_544),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_550),
.B(n_40),
.Y(n_758)
);

OAI21xp5_ASAP7_75t_L g759 ( 
.A1(n_544),
.A2(n_84),
.B(n_127),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_512),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_543),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_486),
.B(n_42),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_501),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_569),
.B(n_43),
.C(n_44),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_602),
.B(n_44),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_602),
.B(n_45),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_549),
.B(n_48),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_518),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_513),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_549),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_553),
.B(n_49),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_553),
.B(n_135),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_623),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_603),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_620),
.A2(n_573),
.B1(n_533),
.B2(n_492),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_620),
.B(n_492),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_667),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_761),
.B(n_550),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_745),
.B(n_688),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_606),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_678),
.B(n_494),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_627),
.A2(n_573),
.B1(n_533),
.B2(n_492),
.Y(n_782)
);

INVxp67_ASAP7_75t_SL g783 ( 
.A(n_692),
.Y(n_783)
);

NOR3xp33_ASAP7_75t_SL g784 ( 
.A(n_720),
.B(n_577),
.C(n_582),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_678),
.B(n_494),
.Y(n_785)
);

A2O1A1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_687),
.A2(n_597),
.B(n_585),
.C(n_598),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_639),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_687),
.A2(n_558),
.B(n_554),
.C(n_598),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_634),
.A2(n_533),
.B1(n_684),
.B2(n_492),
.Y(n_789)
);

NAND2x1p5_ASAP7_75t_L g790 ( 
.A(n_692),
.B(n_694),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_SL g791 ( 
.A1(n_763),
.A2(n_533),
.B1(n_465),
.B2(n_579),
.Y(n_791)
);

NOR3xp33_ASAP7_75t_SL g792 ( 
.A(n_720),
.B(n_565),
.C(n_568),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_667),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_717),
.A2(n_465),
.B1(n_532),
.B2(n_542),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_646),
.B(n_491),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_744),
.B(n_494),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_608),
.B(n_508),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_653),
.Y(n_798)
);

INVx5_ASAP7_75t_L g799 ( 
.A(n_625),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_655),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_663),
.Y(n_801)
);

AND3x1_ASAP7_75t_SL g802 ( 
.A(n_664),
.B(n_558),
.C(n_554),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_744),
.B(n_494),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_626),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_672),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_717),
.A2(n_465),
.B1(n_522),
.B2(n_535),
.Y(n_806)
);

NAND2x1p5_ASAP7_75t_L g807 ( 
.A(n_692),
.B(n_578),
.Y(n_807)
);

CKINVDCx11_ASAP7_75t_R g808 ( 
.A(n_636),
.Y(n_808)
);

NAND2xp33_ASAP7_75t_L g809 ( 
.A(n_625),
.B(n_565),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_695),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_608),
.B(n_568),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_645),
.B(n_618),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_626),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_695),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_651),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_676),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_692),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_SL g818 ( 
.A1(n_622),
.A2(n_548),
.B1(n_582),
.B2(n_596),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_689),
.Y(n_819)
);

A2O1A1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_705),
.A2(n_585),
.B(n_596),
.C(n_571),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_611),
.B(n_571),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_743),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_702),
.B(n_494),
.Y(n_823)
);

BUFx12f_ASAP7_75t_L g824 ( 
.A(n_743),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_740),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_613),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_611),
.B(n_589),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_694),
.B(n_731),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_615),
.B(n_589),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_690),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_698),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_694),
.B(n_521),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_637),
.B(n_536),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_718),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_630),
.B(n_600),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_722),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_738),
.Y(n_837)
);

NOR2x2_ASAP7_75t_L g838 ( 
.A(n_704),
.B(n_456),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_710),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_709),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_694),
.Y(n_841)
);

NOR2x2_ASAP7_75t_L g842 ( 
.A(n_660),
.B(n_456),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_731),
.B(n_737),
.Y(n_843)
);

NOR2x1p5_ASAP7_75t_L g844 ( 
.A(n_656),
.B(n_538),
.Y(n_844)
);

INVx1_ASAP7_75t_SL g845 ( 
.A(n_753),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_746),
.Y(n_846)
);

CKINVDCx11_ASAP7_75t_R g847 ( 
.A(n_753),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_740),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_723),
.Y(n_849)
);

NOR2x2_ASAP7_75t_L g850 ( 
.A(n_656),
.B(n_638),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_754),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_755),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_680),
.B(n_601),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_731),
.Y(n_854)
);

INVx5_ASAP7_75t_L g855 ( 
.A(n_625),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_604),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_739),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_731),
.B(n_521),
.Y(n_858)
);

NOR2x2_ASAP7_75t_L g859 ( 
.A(n_638),
.B(n_461),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_756),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_607),
.B(n_601),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_757),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_R g863 ( 
.A(n_670),
.B(n_523),
.Y(n_863)
);

NAND3xp33_ASAP7_75t_SL g864 ( 
.A(n_633),
.B(n_531),
.C(n_463),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_675),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_683),
.B(n_594),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_770),
.A2(n_521),
.B1(n_500),
.B2(n_505),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_677),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_719),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_719),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_616),
.A2(n_505),
.B1(n_463),
.B2(n_469),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_605),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_640),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_683),
.B(n_594),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_701),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_679),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_736),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_617),
.B(n_522),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_682),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_673),
.B(n_513),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_767),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_658),
.B(n_505),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_658),
.B(n_483),
.Y(n_883)
);

BUFx12f_ASAP7_75t_L g884 ( 
.A(n_736),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_771),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_751),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_R g887 ( 
.A(n_640),
.B(n_526),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_621),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_681),
.B(n_685),
.Y(n_889)
);

AND3x1_ASAP7_75t_L g890 ( 
.A(n_629),
.B(n_519),
.C(n_493),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_705),
.A2(n_524),
.B(n_520),
.C(n_532),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_693),
.B(n_483),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_762),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_696),
.B(n_524),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_610),
.B(n_546),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_612),
.B(n_716),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_659),
.B(n_473),
.Y(n_897)
);

NOR2x1p5_ASAP7_75t_L g898 ( 
.A(n_726),
.B(n_764),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_713),
.B(n_520),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_628),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_716),
.B(n_535),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_706),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_659),
.B(n_461),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_724),
.B(n_546),
.Y(n_904)
);

INVxp67_ASAP7_75t_SL g905 ( 
.A(n_686),
.Y(n_905)
);

O2A1O1Ixp5_ASAP7_75t_L g906 ( 
.A1(n_648),
.A2(n_519),
.B(n_493),
.C(n_539),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_633),
.B(n_542),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_724),
.B(n_465),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_727),
.B(n_465),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_707),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_730),
.A2(n_465),
.B1(n_469),
.B2(n_473),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_666),
.B(n_539),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_714),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_732),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_747),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_654),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_750),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_632),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_727),
.B(n_465),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_760),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_661),
.B(n_578),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_666),
.B(n_560),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_768),
.A2(n_555),
.B1(n_578),
.B2(n_586),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_772),
.B(n_539),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_730),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_643),
.B(n_649),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_SL g927 ( 
.A(n_741),
.B(n_526),
.C(n_523),
.Y(n_927)
);

BUFx8_ASAP7_75t_L g928 ( 
.A(n_642),
.Y(n_928)
);

INVx4_ASAP7_75t_L g929 ( 
.A(n_644),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_769),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_765),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_629),
.B(n_572),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_652),
.B(n_560),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_735),
.A2(n_555),
.B1(n_586),
.B2(n_578),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_665),
.B(n_560),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_741),
.A2(n_560),
.B(n_576),
.C(n_572),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_671),
.Y(n_937)
);

NAND3xp33_ASAP7_75t_SL g938 ( 
.A(n_635),
.B(n_587),
.C(n_584),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_752),
.B(n_556),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_752),
.B(n_556),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_759),
.B(n_493),
.Y(n_941)
);

NAND2xp33_ASAP7_75t_L g942 ( 
.A(n_766),
.B(n_609),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_668),
.B(n_669),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_648),
.B(n_556),
.Y(n_944)
);

BUFx5_ASAP7_75t_L g945 ( 
.A(n_721),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_641),
.B(n_556),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_735),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_748),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_742),
.B(n_576),
.Y(n_949)
);

NOR2x2_ASAP7_75t_L g950 ( 
.A(n_650),
.B(n_587),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_725),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_729),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_748),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_749),
.A2(n_555),
.B1(n_586),
.B2(n_578),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_650),
.B(n_563),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_749),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_734),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_758),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_758),
.B(n_519),
.Y(n_959)
);

OR2x6_ASAP7_75t_L g960 ( 
.A(n_721),
.B(n_562),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_773),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_784),
.A2(n_674),
.B(n_711),
.C(n_715),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_804),
.B(n_563),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_813),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_784),
.A2(n_697),
.B(n_712),
.C(n_708),
.Y(n_965)
);

AO31x2_ASAP7_75t_L g966 ( 
.A1(n_891),
.A2(n_703),
.A3(n_551),
.B(n_562),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_884),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_811),
.A2(n_733),
.B(n_728),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_856),
.B(n_609),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_889),
.A2(n_614),
.B(n_624),
.C(n_631),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_791),
.A2(n_647),
.B1(n_619),
.B2(n_624),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_SL g972 ( 
.A1(n_786),
.A2(n_647),
.B(n_619),
.C(n_631),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_804),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_777),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_821),
.A2(n_733),
.B(n_728),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_824),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_793),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_780),
.B(n_779),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_810),
.Y(n_979)
);

NOR3xp33_ASAP7_75t_L g980 ( 
.A(n_818),
.B(n_614),
.C(n_699),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_928),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_779),
.B(n_563),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_872),
.A2(n_916),
.B1(n_937),
.B2(n_775),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_816),
.B(n_555),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_845),
.B(n_572),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_827),
.A2(n_700),
.B(n_691),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_774),
.B(n_586),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_941),
.A2(n_700),
.B(n_691),
.Y(n_988)
);

OAI33xp33_ASAP7_75t_L g989 ( 
.A1(n_812),
.A2(n_657),
.A3(n_580),
.B1(n_584),
.B2(n_583),
.B3(n_559),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_835),
.B(n_563),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_787),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_815),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_792),
.A2(n_657),
.B1(n_662),
.B2(n_576),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_815),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_817),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_941),
.A2(n_493),
.B(n_519),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_795),
.A2(n_782),
.B1(n_789),
.B2(n_797),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_943),
.A2(n_576),
.B(n_572),
.C(n_580),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_900),
.B(n_527),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_SL g1000 ( 
.A1(n_943),
.A2(n_931),
.B(n_942),
.C(n_935),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_939),
.A2(n_539),
.B(n_527),
.Y(n_1001)
);

BUFx12f_ASAP7_75t_L g1002 ( 
.A(n_808),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_792),
.A2(n_551),
.B(n_583),
.C(n_559),
.Y(n_1003)
);

OR2x6_ASAP7_75t_L g1004 ( 
.A(n_822),
.B(n_527),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_925),
.B(n_547),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_798),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_786),
.A2(n_788),
.B(n_882),
.C(n_956),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_940),
.A2(n_547),
.B(n_457),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_795),
.B(n_547),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_826),
.B(n_833),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_829),
.A2(n_547),
.B1(n_578),
.B2(n_586),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_788),
.A2(n_457),
.B(n_547),
.C(n_586),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_926),
.A2(n_457),
.B(n_62),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_928),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_820),
.A2(n_457),
.B1(n_75),
.B2(n_76),
.Y(n_1015)
);

OAI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_881),
.A2(n_457),
.B(n_79),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_924),
.A2(n_457),
.B(n_86),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_853),
.B(n_58),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_826),
.B(n_90),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_924),
.A2(n_922),
.B(n_904),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_857),
.Y(n_1021)
);

NAND2xp33_ASAP7_75t_SL g1022 ( 
.A(n_844),
.B(n_92),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_800),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_849),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_820),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_901),
.A2(n_116),
.B(n_122),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_882),
.B(n_126),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_896),
.B(n_778),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_799),
.B(n_855),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_886),
.A2(n_893),
.B(n_885),
.C(n_776),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_817),
.Y(n_1031)
);

NAND3xp33_ASAP7_75t_L g1032 ( 
.A(n_890),
.B(n_892),
.C(n_789),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_847),
.B(n_839),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_866),
.A2(n_874),
.B(n_809),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_898),
.A2(n_778),
.B1(n_948),
.B2(n_958),
.Y(n_1035)
);

OR2x6_ASAP7_75t_L g1036 ( 
.A(n_840),
.B(n_899),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_L g1037 ( 
.A(n_864),
.B(n_919),
.C(n_908),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_799),
.B(n_855),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_781),
.A2(n_796),
.B(n_785),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_873),
.Y(n_1040)
);

BUFx8_ASAP7_75t_SL g1041 ( 
.A(n_817),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_892),
.A2(n_953),
.B(n_947),
.C(n_944),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_R g1043 ( 
.A(n_799),
.B(n_855),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_801),
.B(n_805),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_781),
.A2(n_796),
.B(n_785),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_842),
.Y(n_1046)
);

AOI21x1_ASAP7_75t_L g1047 ( 
.A1(n_897),
.A2(n_903),
.B(n_912),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_819),
.B(n_830),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_803),
.A2(n_903),
.B(n_897),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_803),
.A2(n_909),
.B(n_912),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_950),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_959),
.A2(n_936),
.B(n_878),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_814),
.Y(n_1053)
);

AOI21x1_ASAP7_75t_L g1054 ( 
.A1(n_843),
.A2(n_823),
.B(n_959),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_873),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_831),
.B(n_834),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_932),
.Y(n_1057)
);

NAND2x1p5_ASAP7_75t_L g1058 ( 
.A(n_799),
.B(n_855),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_836),
.B(n_837),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_846),
.B(n_851),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_907),
.B(n_870),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_852),
.A2(n_860),
.B1(n_862),
.B2(n_794),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_905),
.B(n_948),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_936),
.A2(n_933),
.B(n_895),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_902),
.Y(n_1065)
);

OAI21xp33_ASAP7_75t_L g1066 ( 
.A1(n_935),
.A2(n_880),
.B(n_894),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_870),
.B(n_817),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_891),
.A2(n_927),
.B(n_906),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_949),
.A2(n_858),
.B(n_832),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_888),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_794),
.A2(n_806),
.B1(n_923),
.B2(n_877),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_SL g1072 ( 
.A(n_870),
.B(n_929),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_861),
.B(n_910),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_913),
.B(n_920),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_832),
.A2(n_858),
.B(n_843),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_806),
.A2(n_923),
.B1(n_911),
.B2(n_927),
.Y(n_1076)
);

AOI21x1_ASAP7_75t_L g1077 ( 
.A1(n_823),
.A2(n_883),
.B(n_955),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_825),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_802),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_870),
.B(n_945),
.Y(n_1080)
);

AOI22x1_ASAP7_75t_L g1081 ( 
.A1(n_946),
.A2(n_929),
.B1(n_869),
.B2(n_877),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_790),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_865),
.A2(n_879),
.B1(n_930),
.B2(n_868),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_883),
.B(n_888),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_915),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_850),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_867),
.A2(n_944),
.B(n_871),
.C(n_875),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_918),
.B(n_917),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_848),
.B(n_914),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_876),
.Y(n_1090)
);

NOR2x1_ASAP7_75t_L g1091 ( 
.A(n_921),
.B(n_918),
.Y(n_1091)
);

AOI221xp5_ASAP7_75t_L g1092 ( 
.A1(n_938),
.A2(n_863),
.B1(n_934),
.B2(n_954),
.C(n_887),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_828),
.A2(n_869),
.B(n_783),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_960),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_802),
.A2(n_945),
.B1(n_960),
.B2(n_921),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_828),
.A2(n_960),
.B(n_957),
.C(n_951),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_934),
.A2(n_954),
.B(n_854),
.C(n_841),
.Y(n_1097)
);

INVx8_ASAP7_75t_L g1098 ( 
.A(n_841),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_952),
.B(n_945),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_945),
.A2(n_854),
.B1(n_790),
.B2(n_859),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_945),
.A2(n_863),
.B(n_887),
.C(n_838),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_SL g1102 ( 
.A1(n_807),
.A2(n_872),
.B1(n_856),
.B2(n_501),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_807),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_945),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_799),
.B(n_855),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_792),
.A2(n_784),
.B1(n_811),
.B2(n_775),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_813),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_773),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_811),
.A2(n_827),
.B(n_821),
.Y(n_1109)
);

O2A1O1Ixp5_ASAP7_75t_L g1110 ( 
.A1(n_1106),
.A2(n_1015),
.B(n_1076),
.C(n_1068),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_983),
.B(n_969),
.Y(n_1111)
);

NAND2x1p5_ASAP7_75t_L g1112 ( 
.A(n_981),
.B(n_967),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1106),
.A2(n_1032),
.B(n_1007),
.C(n_970),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1000),
.A2(n_1015),
.B(n_1010),
.C(n_962),
.Y(n_1114)
);

AO21x2_ASAP7_75t_L g1115 ( 
.A1(n_1068),
.A2(n_1064),
.B(n_1052),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_961),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_967),
.Y(n_1117)
);

AO31x2_ASAP7_75t_L g1118 ( 
.A1(n_1076),
.A2(n_965),
.A3(n_1042),
.B(n_1020),
.Y(n_1118)
);

AO31x2_ASAP7_75t_L g1119 ( 
.A1(n_1049),
.A2(n_1109),
.A3(n_1025),
.B(n_1071),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1102),
.A2(n_997),
.B1(n_1057),
.B2(n_1051),
.Y(n_1120)
);

AO22x2_ASAP7_75t_L g1121 ( 
.A1(n_1062),
.A2(n_1025),
.B1(n_1046),
.B2(n_1094),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_SL g1122 ( 
.A1(n_1079),
.A2(n_1086),
.B1(n_1046),
.B2(n_1027),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1107),
.B(n_992),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1047),
.A2(n_1050),
.B(n_1077),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_SL g1125 ( 
.A1(n_1095),
.A2(n_1062),
.B(n_1035),
.Y(n_1125)
);

AOI221x1_ASAP7_75t_L g1126 ( 
.A1(n_980),
.A2(n_1037),
.B1(n_1016),
.B2(n_1066),
.C(n_1075),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_SL g1127 ( 
.A1(n_1019),
.A2(n_1080),
.B(n_1030),
.C(n_1101),
.Y(n_1127)
);

AO21x1_ASAP7_75t_L g1128 ( 
.A1(n_1022),
.A2(n_1096),
.B(n_1012),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_974),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1034),
.A2(n_988),
.A3(n_1084),
.B(n_1045),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_SL g1131 ( 
.A1(n_1029),
.A2(n_1105),
.B(n_1092),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1054),
.A2(n_996),
.B(n_1039),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_968),
.A2(n_975),
.B(n_986),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1017),
.A2(n_1069),
.B(n_1001),
.Y(n_1134)
);

AO32x2_ASAP7_75t_L g1135 ( 
.A1(n_1055),
.A2(n_966),
.A3(n_1014),
.B1(n_1011),
.B2(n_989),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1008),
.A2(n_1099),
.B(n_1061),
.Y(n_1136)
);

AO31x2_ASAP7_75t_L g1137 ( 
.A1(n_1104),
.A2(n_1003),
.A3(n_1097),
.B(n_1011),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_972),
.A2(n_1013),
.B(n_1087),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_1036),
.B(n_1040),
.Y(n_1139)
);

INVxp67_ASAP7_75t_L g1140 ( 
.A(n_964),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1107),
.B(n_994),
.Y(n_1141)
);

AO31x2_ASAP7_75t_L g1142 ( 
.A1(n_1073),
.A2(n_998),
.A3(n_1053),
.B(n_1078),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1044),
.B(n_1060),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1056),
.B(n_982),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1081),
.A2(n_1093),
.B(n_1026),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1048),
.B(n_1059),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1072),
.A2(n_1005),
.B(n_1028),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1058),
.A2(n_1100),
.B(n_1038),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1072),
.A2(n_990),
.B(n_1063),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_963),
.B(n_1108),
.Y(n_1150)
);

AOI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_971),
.A2(n_1018),
.B(n_1088),
.Y(n_1151)
);

CKINVDCx20_ASAP7_75t_R g1152 ( 
.A(n_1002),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1058),
.A2(n_1067),
.B(n_1091),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_1041),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_1033),
.B(n_1023),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_993),
.A2(n_984),
.B(n_991),
.Y(n_1156)
);

AO31x2_ASAP7_75t_L g1157 ( 
.A1(n_977),
.A2(n_979),
.A3(n_1089),
.B(n_1065),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1074),
.A2(n_987),
.B(n_1006),
.Y(n_1158)
);

INVx5_ASAP7_75t_L g1159 ( 
.A(n_967),
.Y(n_1159)
);

O2A1O1Ixp5_ASAP7_75t_SL g1160 ( 
.A1(n_1085),
.A2(n_1090),
.B(n_1021),
.C(n_999),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1009),
.A2(n_1083),
.B(n_985),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1029),
.A2(n_1105),
.B(n_1098),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1004),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1098),
.A2(n_1031),
.B(n_995),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1070),
.B(n_1036),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1004),
.A2(n_1024),
.B1(n_1036),
.B2(n_1098),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_966),
.A2(n_1043),
.B(n_1103),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_976),
.Y(n_1168)
);

INVxp67_ASAP7_75t_L g1169 ( 
.A(n_1082),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_966),
.A2(n_1031),
.B(n_1103),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_SL g1171 ( 
.A(n_1103),
.B(n_1082),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1082),
.A2(n_620),
.B(n_592),
.C(n_925),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1020),
.A2(n_1064),
.B(n_1047),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1010),
.B(n_978),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_961),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_974),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1010),
.B(n_978),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1109),
.A2(n_1034),
.B(n_811),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1010),
.B(n_978),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_981),
.Y(n_1180)
);

AOI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1020),
.A2(n_1064),
.B(n_1047),
.Y(n_1181)
);

BUFx10_ASAP7_75t_L g1182 ( 
.A(n_967),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_SL g1183 ( 
.A1(n_1101),
.A2(n_811),
.B(n_1071),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1041),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_983),
.B(n_622),
.Y(n_1185)
);

NOR4xp25_ASAP7_75t_L g1186 ( 
.A(n_1106),
.B(n_720),
.C(n_1007),
.D(n_629),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1109),
.A2(n_1034),
.B(n_811),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1007),
.A2(n_1106),
.B(n_1052),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_961),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_983),
.B(n_622),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1010),
.B(n_978),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1002),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1049),
.A2(n_1047),
.B(n_1020),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1106),
.A2(n_916),
.B1(n_620),
.B2(n_937),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_978),
.B(n_973),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_983),
.B(n_622),
.Y(n_1196)
);

AOI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1020),
.A2(n_1064),
.B(n_1047),
.Y(n_1197)
);

AOI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1020),
.A2(n_1064),
.B(n_1047),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_981),
.B(n_799),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_1107),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1109),
.A2(n_620),
.B(n_627),
.Y(n_1201)
);

AOI211x1_ASAP7_75t_L g1202 ( 
.A1(n_1106),
.A2(n_720),
.B(n_726),
.C(n_764),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1109),
.A2(n_1034),
.B(n_811),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_964),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1029),
.Y(n_1205)
);

AOI211x1_ASAP7_75t_L g1206 ( 
.A1(n_1106),
.A2(n_720),
.B(n_726),
.C(n_764),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_964),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1076),
.A2(n_891),
.A3(n_965),
.B(n_1064),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1010),
.B(n_978),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1010),
.B(n_978),
.Y(n_1210)
);

NAND3x1_ASAP7_75t_L g1211 ( 
.A(n_983),
.B(n_775),
.C(n_969),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_961),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1109),
.A2(n_1034),
.B(n_811),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1049),
.A2(n_1047),
.B(n_1020),
.Y(n_1214)
);

NAND3xp33_ASAP7_75t_SL g1215 ( 
.A(n_983),
.B(n_872),
.C(n_856),
.Y(n_1215)
);

INVx4_ASAP7_75t_L g1216 ( 
.A(n_1041),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1107),
.Y(n_1217)
);

CKINVDCx8_ASAP7_75t_R g1218 ( 
.A(n_967),
.Y(n_1218)
);

NOR4xp25_ASAP7_75t_L g1219 ( 
.A(n_1106),
.B(n_720),
.C(n_1007),
.D(n_629),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1010),
.B(n_978),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1049),
.A2(n_1047),
.B(n_1020),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_964),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1007),
.A2(n_1106),
.B(n_1052),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1076),
.A2(n_891),
.A3(n_965),
.B(n_1064),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1010),
.B(n_978),
.Y(n_1225)
);

AO32x2_ASAP7_75t_L g1226 ( 
.A1(n_1106),
.A2(n_1076),
.A3(n_1062),
.B1(n_818),
.B2(n_1015),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1010),
.B(n_978),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_SL g1228 ( 
.A1(n_1000),
.A2(n_786),
.B(n_1007),
.C(n_788),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1029),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1076),
.A2(n_891),
.A3(n_965),
.B(n_1064),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_SL g1231 ( 
.A1(n_1106),
.A2(n_1095),
.B(n_1062),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1010),
.B(n_978),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1049),
.A2(n_1047),
.B(n_1020),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1106),
.A2(n_916),
.B1(n_620),
.B2(n_937),
.Y(n_1234)
);

NOR2xp67_ASAP7_75t_L g1235 ( 
.A(n_1029),
.B(n_1105),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1107),
.B(n_804),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1109),
.A2(n_1034),
.B(n_811),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_964),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_SL g1239 ( 
.A1(n_1106),
.A2(n_1095),
.B(n_1062),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1010),
.B(n_978),
.Y(n_1240)
);

OA21x2_ASAP7_75t_L g1241 ( 
.A1(n_1068),
.A2(n_1020),
.B(n_1064),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1010),
.B(n_978),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1010),
.B(n_978),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1106),
.A2(n_916),
.B1(n_620),
.B2(n_937),
.Y(n_1244)
);

CKINVDCx14_ASAP7_75t_R g1245 ( 
.A(n_1002),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1106),
.A2(n_916),
.B1(n_620),
.B2(n_937),
.Y(n_1246)
);

OA21x2_ASAP7_75t_L g1247 ( 
.A1(n_1068),
.A2(n_1020),
.B(n_1064),
.Y(n_1247)
);

INVxp67_ASAP7_75t_SL g1248 ( 
.A(n_964),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_974),
.Y(n_1249)
);

NAND3xp33_ASAP7_75t_SL g1250 ( 
.A(n_1194),
.B(n_1244),
.C(n_1234),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1185),
.A2(n_1196),
.B1(n_1190),
.B2(n_1111),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1235),
.B(n_1205),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1143),
.B(n_1174),
.Y(n_1253)
);

OA21x2_ASAP7_75t_L g1254 ( 
.A1(n_1133),
.A2(n_1126),
.B(n_1110),
.Y(n_1254)
);

OA21x2_ASAP7_75t_L g1255 ( 
.A1(n_1193),
.A2(n_1221),
.B(n_1214),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1246),
.A2(n_1215),
.B1(n_1121),
.B2(n_1120),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1257)
);

AO21x2_ASAP7_75t_L g1258 ( 
.A1(n_1170),
.A2(n_1138),
.B(n_1203),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1181),
.A2(n_1197),
.B(n_1198),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1226),
.B(n_1188),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1233),
.A2(n_1223),
.B(n_1188),
.Y(n_1261)
);

INVx4_ASAP7_75t_L g1262 ( 
.A(n_1139),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1128),
.A2(n_1113),
.A3(n_1187),
.B(n_1213),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1236),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1237),
.A2(n_1132),
.B(n_1124),
.Y(n_1265)
);

BUFx12f_ASAP7_75t_L g1266 ( 
.A(n_1184),
.Y(n_1266)
);

AO21x2_ASAP7_75t_L g1267 ( 
.A1(n_1170),
.A2(n_1151),
.B(n_1125),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1114),
.A2(n_1228),
.B(n_1172),
.C(n_1223),
.Y(n_1268)
);

OA21x2_ASAP7_75t_L g1269 ( 
.A1(n_1167),
.A2(n_1239),
.B(n_1231),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1136),
.A2(n_1241),
.B(n_1247),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1177),
.B(n_1179),
.Y(n_1271)
);

O2A1O1Ixp5_ASAP7_75t_L g1272 ( 
.A1(n_1156),
.A2(n_1149),
.B(n_1147),
.C(n_1141),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1241),
.A2(n_1247),
.B(n_1148),
.Y(n_1273)
);

NAND2x1p5_ASAP7_75t_L g1274 ( 
.A(n_1235),
.B(n_1205),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1158),
.A2(n_1153),
.B(n_1160),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1183),
.A2(n_1164),
.B(n_1161),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1229),
.B(n_1162),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1161),
.A2(n_1163),
.B(n_1131),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1211),
.A2(n_1202),
.B1(n_1206),
.B2(n_1144),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1229),
.B(n_1139),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1157),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1226),
.B(n_1186),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1157),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1115),
.A2(n_1127),
.B(n_1146),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1175),
.A2(n_1189),
.B(n_1212),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1226),
.A2(n_1122),
.B(n_1186),
.C(n_1219),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1150),
.A2(n_1249),
.B(n_1129),
.Y(n_1287)
);

O2A1O1Ixp33_ASAP7_75t_L g1288 ( 
.A1(n_1219),
.A2(n_1227),
.B(n_1243),
.C(n_1242),
.Y(n_1288)
);

BUFx2_ASAP7_75t_SL g1289 ( 
.A(n_1218),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1207),
.Y(n_1290)
);

AO21x2_ASAP7_75t_L g1291 ( 
.A1(n_1115),
.A2(n_1176),
.B(n_1225),
.Y(n_1291)
);

AO32x2_ASAP7_75t_L g1292 ( 
.A1(n_1166),
.A2(n_1121),
.A3(n_1135),
.B1(n_1118),
.B2(n_1224),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1191),
.B(n_1232),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1119),
.A2(n_1118),
.B(n_1224),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1119),
.A2(n_1210),
.B(n_1209),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_SL g1296 ( 
.A1(n_1122),
.A2(n_1155),
.B1(n_1240),
.B2(n_1220),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1202),
.A2(n_1206),
.B(n_1119),
.C(n_1217),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1248),
.A2(n_1140),
.B(n_1238),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1130),
.A2(n_1199),
.B(n_1165),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1142),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1130),
.A2(n_1208),
.B(n_1230),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1204),
.A2(n_1222),
.B1(n_1123),
.B2(n_1200),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1169),
.B(n_1195),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1171),
.A2(n_1118),
.B(n_1230),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1184),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1159),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1168),
.A2(n_1112),
.B(n_1171),
.Y(n_1307)
);

NAND2x1p5_ASAP7_75t_L g1308 ( 
.A(n_1159),
.B(n_1117),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1130),
.A2(n_1208),
.B(n_1230),
.Y(n_1309)
);

AO21x1_ASAP7_75t_L g1310 ( 
.A1(n_1135),
.A2(n_1224),
.B(n_1208),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1154),
.A2(n_1159),
.B1(n_1216),
.B2(n_1184),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1216),
.B(n_1137),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1137),
.A2(n_1182),
.B(n_1180),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1245),
.A2(n_1152),
.B(n_1182),
.C(n_1137),
.Y(n_1314)
);

AO21x2_ASAP7_75t_L g1315 ( 
.A1(n_1192),
.A2(n_1170),
.B(n_1068),
.Y(n_1315)
);

OA21x2_ASAP7_75t_L g1316 ( 
.A1(n_1133),
.A2(n_1126),
.B(n_1110),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_SL g1317 ( 
.A1(n_1113),
.A2(n_1007),
.B(n_1000),
.C(n_1201),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1194),
.B(n_1234),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1226),
.B(n_1188),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1139),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1236),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1136),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_SL g1326 ( 
.A1(n_1111),
.A2(n_1185),
.B1(n_1196),
.B2(n_1190),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1226),
.B(n_1188),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1235),
.B(n_1205),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1111),
.A2(n_1246),
.B1(n_1244),
.B2(n_1234),
.Y(n_1331)
);

NAND2x1p5_ASAP7_75t_L g1332 ( 
.A(n_1235),
.B(n_1205),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1245),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1139),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1194),
.A2(n_620),
.B(n_1234),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1116),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1194),
.A2(n_620),
.B(n_1234),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1185),
.A2(n_1196),
.B1(n_1190),
.B2(n_501),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1226),
.B(n_1188),
.Y(n_1342)
);

AOI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1138),
.A2(n_1181),
.B(n_1173),
.Y(n_1343)
);

O2A1O1Ixp33_ASAP7_75t_SL g1344 ( 
.A1(n_1113),
.A2(n_1007),
.B(n_1000),
.C(n_1201),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1226),
.B(n_1188),
.Y(n_1345)
);

NAND2x1p5_ASAP7_75t_L g1346 ( 
.A(n_1235),
.B(n_1205),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_SL g1347 ( 
.A(n_1218),
.B(n_1002),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1143),
.B(n_1174),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1139),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1226),
.B(n_1188),
.Y(n_1351)
);

OR2x6_ASAP7_75t_L g1352 ( 
.A(n_1131),
.B(n_1183),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1194),
.A2(n_1234),
.B1(n_1246),
.B2(n_1244),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1355)
);

AOI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1138),
.A2(n_1181),
.B(n_1173),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1201),
.A2(n_1109),
.B(n_1178),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1116),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1194),
.A2(n_1244),
.B(n_1246),
.C(n_1234),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1143),
.B(n_1174),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1157),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1194),
.A2(n_620),
.B(n_1234),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1157),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1226),
.B(n_1188),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1133),
.A2(n_1126),
.B(n_1110),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1205),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1194),
.B(n_1234),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1134),
.A2(n_1145),
.B(n_1173),
.Y(n_1372)
);

AO21x2_ASAP7_75t_L g1373 ( 
.A1(n_1170),
.A2(n_1068),
.B(n_1138),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1116),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1185),
.A2(n_1196),
.B1(n_1190),
.B2(n_501),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1111),
.A2(n_1246),
.B1(n_1244),
.B2(n_1234),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1257),
.A2(n_1323),
.B(n_1322),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_1308),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1285),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1337),
.A2(n_1364),
.B(n_1339),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1261),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_SL g1382 ( 
.A1(n_1352),
.A2(n_1359),
.B(n_1354),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1264),
.B(n_1321),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1331),
.A2(n_1376),
.B1(n_1251),
.B2(n_1318),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1290),
.B(n_1271),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1312),
.B(n_1260),
.Y(n_1386)
);

INVxp67_ASAP7_75t_L g1387 ( 
.A(n_1290),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1318),
.A2(n_1371),
.B1(n_1326),
.B2(n_1340),
.Y(n_1388)
);

O2A1O1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1250),
.A2(n_1371),
.B(n_1317),
.C(n_1344),
.Y(n_1389)
);

O2A1O1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1317),
.A2(n_1344),
.B(n_1375),
.C(n_1268),
.Y(n_1390)
);

OA22x2_ASAP7_75t_L g1391 ( 
.A1(n_1352),
.A2(n_1319),
.B1(n_1367),
.B2(n_1328),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1349),
.B(n_1361),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1303),
.B(n_1350),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1256),
.A2(n_1286),
.B1(n_1352),
.B2(n_1282),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1350),
.B(n_1320),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1261),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1357),
.A2(n_1352),
.B(n_1284),
.Y(n_1397)
);

NOR2xp67_ASAP7_75t_L g1398 ( 
.A(n_1311),
.B(n_1306),
.Y(n_1398)
);

O2A1O1Ixp5_ASAP7_75t_L g1399 ( 
.A1(n_1286),
.A2(n_1272),
.B(n_1297),
.C(n_1279),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_SL g1400 ( 
.A1(n_1314),
.A2(n_1288),
.B(n_1295),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1293),
.B(n_1302),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1260),
.A2(n_1328),
.B1(n_1319),
.B2(n_1345),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1297),
.A2(n_1298),
.B(n_1342),
.C(n_1351),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1342),
.B(n_1345),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1320),
.B(n_1335),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1296),
.A2(n_1367),
.B1(n_1351),
.B2(n_1347),
.Y(n_1406)
);

INVx2_ASAP7_75t_SL g1407 ( 
.A(n_1305),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1335),
.B(n_1280),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1333),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1312),
.B(n_1277),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1289),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1333),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1280),
.B(n_1315),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_1266),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1338),
.B(n_1358),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1374),
.B(n_1280),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1261),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1287),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1266),
.Y(n_1419)
);

OA21x2_ASAP7_75t_L g1420 ( 
.A1(n_1325),
.A2(n_1341),
.B(n_1334),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1291),
.B(n_1262),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1291),
.B(n_1262),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1262),
.A2(n_1316),
.B1(n_1254),
.B2(n_1369),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1281),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1301),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1369),
.A2(n_1305),
.B1(n_1269),
.B2(n_1277),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1308),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1315),
.Y(n_1428)
);

O2A1O1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1307),
.A2(n_1304),
.B(n_1306),
.C(n_1324),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_SL g1430 ( 
.A1(n_1252),
.A2(n_1329),
.B(n_1274),
.Y(n_1430)
);

O2A1O1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1324),
.A2(n_1373),
.B(n_1310),
.C(n_1267),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1283),
.Y(n_1432)
);

AOI211xp5_ASAP7_75t_L g1433 ( 
.A1(n_1276),
.A2(n_1313),
.B(n_1299),
.C(n_1309),
.Y(n_1433)
);

AOI21x1_ASAP7_75t_SL g1434 ( 
.A1(n_1252),
.A2(n_1263),
.B(n_1356),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_SL g1435 ( 
.A1(n_1274),
.A2(n_1346),
.B(n_1332),
.Y(n_1435)
);

OA21x2_ASAP7_75t_L g1436 ( 
.A1(n_1325),
.A2(n_1372),
.B(n_1368),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1327),
.A2(n_1372),
.B(n_1368),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1283),
.Y(n_1438)
);

O2A1O1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1267),
.A2(n_1258),
.B(n_1269),
.C(n_1294),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1327),
.A2(n_1330),
.B(n_1363),
.Y(n_1440)
);

OAI211xp5_ASAP7_75t_L g1441 ( 
.A1(n_1294),
.A2(n_1343),
.B(n_1269),
.C(n_1299),
.Y(n_1441)
);

AND2x4_ASAP7_75t_SL g1442 ( 
.A(n_1370),
.B(n_1300),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1278),
.B(n_1276),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1278),
.B(n_1273),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1292),
.B(n_1332),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1329),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1346),
.A2(n_1294),
.B1(n_1255),
.B2(n_1263),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1273),
.B(n_1270),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1292),
.B(n_1263),
.Y(n_1449)
);

AOI21x1_ASAP7_75t_SL g1450 ( 
.A1(n_1275),
.A2(n_1259),
.B(n_1255),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1255),
.A2(n_1292),
.B1(n_1362),
.B2(n_1366),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1292),
.A2(n_1275),
.B(n_1259),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1265),
.A2(n_1330),
.B(n_1334),
.C(n_1336),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1265),
.B(n_1336),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_SL g1455 ( 
.A1(n_1348),
.A2(n_1353),
.B(n_1355),
.Y(n_1455)
);

CKINVDCx14_ASAP7_75t_R g1456 ( 
.A(n_1353),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1355),
.B(n_1365),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1365),
.A2(n_1360),
.B(n_1363),
.Y(n_1458)
);

OA22x2_ASAP7_75t_L g1459 ( 
.A1(n_1360),
.A2(n_1326),
.B1(n_1339),
.B2(n_1337),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1333),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1264),
.B(n_1253),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1379),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1404),
.B(n_1402),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1456),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1456),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1448),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1450),
.A2(n_1458),
.B(n_1397),
.Y(n_1467)
);

OA21x2_ASAP7_75t_L g1468 ( 
.A1(n_1380),
.A2(n_1399),
.B(n_1441),
.Y(n_1468)
);

OR2x6_ASAP7_75t_L g1469 ( 
.A(n_1391),
.B(n_1443),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1410),
.B(n_1443),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1418),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1401),
.B(n_1449),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1384),
.A2(n_1389),
.B(n_1388),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1386),
.B(n_1381),
.Y(n_1474)
);

AND2x4_ASAP7_75t_SL g1475 ( 
.A(n_1410),
.B(n_1386),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1385),
.Y(n_1476)
);

OR2x6_ASAP7_75t_L g1477 ( 
.A(n_1391),
.B(n_1443),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1439),
.A2(n_1434),
.B(n_1453),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1396),
.B(n_1417),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1415),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1444),
.B(n_1448),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1421),
.B(n_1422),
.Y(n_1482)
);

AO21x2_ASAP7_75t_L g1483 ( 
.A1(n_1452),
.A2(n_1451),
.B(n_1400),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1423),
.A2(n_1431),
.B(n_1447),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1445),
.B(n_1425),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1428),
.B(n_1426),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1382),
.B(n_1459),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1413),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_SL g1489 ( 
.A1(n_1390),
.A2(n_1394),
.B(n_1403),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1461),
.B(n_1383),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1459),
.A2(n_1406),
.B1(n_1392),
.B2(n_1387),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1457),
.B(n_1454),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1416),
.B(n_1429),
.Y(n_1493)
);

OR2x6_ASAP7_75t_L g1494 ( 
.A(n_1430),
.B(n_1435),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1411),
.B(n_1407),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1414),
.A2(n_1446),
.B1(n_1409),
.B2(n_1398),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1377),
.B(n_1437),
.Y(n_1497)
);

AO21x2_ASAP7_75t_L g1498 ( 
.A1(n_1455),
.A2(n_1432),
.B(n_1424),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1471),
.Y(n_1499)
);

AO21x2_ASAP7_75t_L g1500 ( 
.A1(n_1484),
.A2(n_1438),
.B(n_1433),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1492),
.B(n_1377),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1492),
.B(n_1481),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1497),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1469),
.Y(n_1504)
);

AOI21xp5_ASAP7_75t_SL g1505 ( 
.A1(n_1487),
.A2(n_1378),
.B(n_1427),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1497),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1479),
.B(n_1393),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1473),
.A2(n_1408),
.B1(n_1405),
.B2(n_1414),
.Y(n_1508)
);

NOR2x1_ASAP7_75t_L g1509 ( 
.A(n_1483),
.B(n_1436),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1471),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1463),
.B(n_1436),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1481),
.Y(n_1512)
);

AND2x4_ASAP7_75t_SL g1513 ( 
.A(n_1470),
.B(n_1395),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1466),
.B(n_1442),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1498),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1498),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1479),
.B(n_1420),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1463),
.B(n_1472),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1462),
.Y(n_1519)
);

NOR2x1_ASAP7_75t_L g1520 ( 
.A(n_1483),
.B(n_1420),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1474),
.B(n_1440),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1518),
.B(n_1472),
.Y(n_1522)
);

AND2x2_ASAP7_75t_SL g1523 ( 
.A(n_1513),
.B(n_1475),
.Y(n_1523)
);

AO21x2_ASAP7_75t_L g1524 ( 
.A1(n_1515),
.A2(n_1484),
.B(n_1483),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1499),
.Y(n_1525)
);

OAI33xp33_ASAP7_75t_L g1526 ( 
.A1(n_1511),
.A2(n_1491),
.A3(n_1493),
.B1(n_1482),
.B2(n_1490),
.B3(n_1480),
.Y(n_1526)
);

NAND3xp33_ASAP7_75t_L g1527 ( 
.A(n_1509),
.B(n_1473),
.C(n_1487),
.Y(n_1527)
);

OAI21xp5_ASAP7_75t_SL g1528 ( 
.A1(n_1508),
.A2(n_1491),
.B(n_1496),
.Y(n_1528)
);

AOI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1517),
.A2(n_1489),
.B1(n_1493),
.B2(n_1483),
.C(n_1484),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1499),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1518),
.B(n_1476),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1500),
.A2(n_1489),
.B1(n_1469),
.B2(n_1477),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_SL g1533 ( 
.A1(n_1504),
.A2(n_1484),
.B1(n_1465),
.B2(n_1464),
.Y(n_1533)
);

OAI221xp5_ASAP7_75t_L g1534 ( 
.A1(n_1508),
.A2(n_1486),
.B1(n_1496),
.B2(n_1464),
.C(n_1465),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1509),
.A2(n_1478),
.B(n_1467),
.Y(n_1535)
);

AND2x2_ASAP7_75t_SL g1536 ( 
.A(n_1513),
.B(n_1475),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1503),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1500),
.A2(n_1477),
.B1(n_1469),
.B2(n_1488),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1510),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1508),
.A2(n_1463),
.B1(n_1468),
.B2(n_1477),
.Y(n_1540)
);

INVx4_ASAP7_75t_L g1541 ( 
.A(n_1514),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1502),
.B(n_1485),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1519),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1519),
.Y(n_1544)
);

NAND3xp33_ASAP7_75t_L g1545 ( 
.A(n_1509),
.B(n_1468),
.C(n_1486),
.Y(n_1545)
);

INVxp67_ASAP7_75t_L g1546 ( 
.A(n_1507),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1502),
.B(n_1485),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1510),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1518),
.B(n_1490),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1527),
.A2(n_1529),
.B(n_1528),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1524),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1525),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1524),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1524),
.Y(n_1554)
);

OA21x2_ASAP7_75t_L g1555 ( 
.A1(n_1545),
.A2(n_1515),
.B(n_1516),
.Y(n_1555)
);

AND4x1_ASAP7_75t_L g1556 ( 
.A(n_1527),
.B(n_1520),
.C(n_1505),
.D(n_1495),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1530),
.Y(n_1557)
);

INVxp67_ASAP7_75t_SL g1558 ( 
.A(n_1545),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1537),
.B(n_1511),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1540),
.A2(n_1468),
.B(n_1494),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1535),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1535),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1541),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1543),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1539),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1522),
.B(n_1518),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1548),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1523),
.B(n_1520),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1542),
.B(n_1506),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1541),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1541),
.B(n_1512),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_SL g1572 ( 
.A(n_1558),
.B(n_1523),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1566),
.B(n_1549),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1550),
.B(n_1549),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1566),
.B(n_1531),
.Y(n_1575)
);

AOI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1550),
.A2(n_1526),
.B1(n_1532),
.B2(n_1533),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1555),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1555),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1565),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1555),
.Y(n_1580)
);

NAND2x1p5_ASAP7_75t_L g1581 ( 
.A(n_1556),
.B(n_1523),
.Y(n_1581)
);

NOR2x1_ASAP7_75t_L g1582 ( 
.A(n_1550),
.B(n_1409),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1564),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1565),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1565),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1555),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1558),
.B(n_1536),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1567),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1563),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1558),
.B(n_1536),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1567),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1563),
.B(n_1536),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1564),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1567),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1564),
.B(n_1412),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1552),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1569),
.B(n_1546),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1563),
.B(n_1541),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1563),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1552),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1570),
.B(n_1542),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1559),
.B(n_1544),
.Y(n_1602)
);

NAND2xp33_ASAP7_75t_R g1603 ( 
.A(n_1570),
.B(n_1412),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1552),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1557),
.Y(n_1605)
);

OR2x6_ASAP7_75t_L g1606 ( 
.A(n_1560),
.B(n_1494),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1555),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1570),
.B(n_1547),
.Y(n_1608)
);

OAI31xp33_ASAP7_75t_L g1609 ( 
.A1(n_1561),
.A2(n_1534),
.A3(n_1538),
.B(n_1486),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1559),
.B(n_1517),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1559),
.B(n_1517),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1604),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1582),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1574),
.B(n_1569),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1577),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1593),
.Y(n_1616)
);

INVxp67_ASAP7_75t_L g1617 ( 
.A(n_1595),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1581),
.B(n_1570),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1596),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1583),
.B(n_1569),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1581),
.B(n_1587),
.Y(n_1621)
);

OAI21xp33_ASAP7_75t_SL g1622 ( 
.A1(n_1587),
.A2(n_1568),
.B(n_1560),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1575),
.B(n_1557),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1576),
.B(n_1569),
.Y(n_1624)
);

OR2x6_ASAP7_75t_L g1625 ( 
.A(n_1606),
.B(n_1494),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1577),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1600),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1573),
.B(n_1521),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1575),
.B(n_1557),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1581),
.B(n_1590),
.Y(n_1630)
);

CKINVDCx16_ASAP7_75t_R g1631 ( 
.A(n_1603),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1605),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1585),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1573),
.B(n_1521),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1590),
.B(n_1521),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1578),
.Y(n_1636)
);

OAI21xp33_ASAP7_75t_L g1637 ( 
.A1(n_1572),
.A2(n_1562),
.B(n_1561),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1578),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1580),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1592),
.B(n_1571),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1585),
.Y(n_1641)
);

NOR2x1p5_ASAP7_75t_SL g1642 ( 
.A(n_1580),
.B(n_1551),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1599),
.B(n_1521),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1609),
.A2(n_1556),
.B(n_1520),
.Y(n_1644)
);

OAI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1606),
.A2(n_1556),
.B1(n_1561),
.B2(n_1562),
.C(n_1555),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1597),
.B(n_1501),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1619),
.Y(n_1647)
);

INVx1_ASAP7_75t_SL g1648 ( 
.A(n_1631),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1615),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1631),
.B(n_1460),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1615),
.Y(n_1651)
);

AOI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1624),
.A2(n_1622),
.B1(n_1645),
.B2(n_1630),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1616),
.B(n_1601),
.Y(n_1653)
);

CKINVDCx16_ASAP7_75t_R g1654 ( 
.A(n_1613),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1617),
.B(n_1601),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1621),
.B(n_1592),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1619),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1621),
.B(n_1608),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1627),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1626),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1612),
.B(n_1608),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1630),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1612),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1613),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1618),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1623),
.B(n_1602),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1627),
.Y(n_1667)
);

OR2x6_ASAP7_75t_L g1668 ( 
.A(n_1625),
.B(n_1606),
.Y(n_1668)
);

CKINVDCx16_ASAP7_75t_R g1669 ( 
.A(n_1644),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1622),
.A2(n_1606),
.B1(n_1586),
.B2(n_1607),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1618),
.Y(n_1671)
);

O2A1O1Ixp33_ASAP7_75t_SL g1672 ( 
.A1(n_1648),
.A2(n_1637),
.B(n_1589),
.C(n_1614),
.Y(n_1672)
);

AOI21xp33_ASAP7_75t_L g1673 ( 
.A1(n_1664),
.A2(n_1641),
.B(n_1633),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1647),
.Y(n_1674)
);

NOR4xp75_ASAP7_75t_L g1675 ( 
.A(n_1655),
.B(n_1620),
.C(n_1640),
.D(n_1635),
.Y(n_1675)
);

OAI22xp33_ASAP7_75t_SL g1676 ( 
.A1(n_1669),
.A2(n_1607),
.B1(n_1586),
.B2(n_1625),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1654),
.B(n_1623),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1658),
.B(n_1656),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1669),
.A2(n_1652),
.B1(n_1654),
.B2(n_1656),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1658),
.Y(n_1680)
);

INVx1_ASAP7_75t_SL g1681 ( 
.A(n_1662),
.Y(n_1681)
);

AOI21xp33_ASAP7_75t_SL g1682 ( 
.A1(n_1650),
.A2(n_1589),
.B(n_1568),
.Y(n_1682)
);

A2O1A1Ixp33_ASAP7_75t_L g1683 ( 
.A1(n_1670),
.A2(n_1642),
.B(n_1562),
.C(n_1561),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1647),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1671),
.B(n_1640),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1665),
.B(n_1629),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1657),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1671),
.Y(n_1688)
);

AOI322xp5_ASAP7_75t_L g1689 ( 
.A1(n_1649),
.A2(n_1634),
.A3(n_1628),
.B1(n_1626),
.B2(n_1636),
.C1(n_1638),
.C2(n_1639),
.Y(n_1689)
);

OAI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1668),
.A2(n_1625),
.B1(n_1562),
.B2(n_1561),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1678),
.B(n_1653),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1680),
.B(n_1663),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1680),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1681),
.B(n_1666),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1674),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1677),
.B(n_1666),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1688),
.B(n_1685),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1684),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1686),
.B(n_1661),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_SL g1700 ( 
.A1(n_1679),
.A2(n_1419),
.B1(n_1667),
.B2(n_1659),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1687),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1700),
.A2(n_1683),
.B1(n_1676),
.B2(n_1690),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1696),
.A2(n_1683),
.B1(n_1690),
.B2(n_1649),
.Y(n_1703)
);

NAND4xp25_ASAP7_75t_L g1704 ( 
.A(n_1694),
.B(n_1673),
.C(n_1672),
.D(n_1682),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1692),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1691),
.A2(n_1672),
.B(n_1660),
.Y(n_1706)
);

NAND3xp33_ASAP7_75t_SL g1707 ( 
.A(n_1693),
.B(n_1675),
.C(n_1689),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1697),
.B(n_1657),
.Y(n_1708)
);

OAI31xp33_ASAP7_75t_L g1709 ( 
.A1(n_1701),
.A2(n_1660),
.A3(n_1651),
.B(n_1562),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_SL g1710 ( 
.A(n_1697),
.B(n_1651),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1708),
.Y(n_1711)
);

NAND4xp25_ASAP7_75t_L g1712 ( 
.A(n_1706),
.B(n_1699),
.C(n_1698),
.D(n_1695),
.Y(n_1712)
);

OAI211xp5_ASAP7_75t_SL g1713 ( 
.A1(n_1702),
.A2(n_1667),
.B(n_1659),
.C(n_1633),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1703),
.A2(n_1629),
.B1(n_1643),
.B2(n_1668),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1710),
.B(n_1632),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1711),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1715),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1712),
.B(n_1705),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1714),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1713),
.B(n_1598),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1715),
.Y(n_1721)
);

A2O1A1Ixp33_ASAP7_75t_L g1722 ( 
.A1(n_1718),
.A2(n_1707),
.B(n_1709),
.C(n_1704),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1716),
.Y(n_1723)
);

NOR2x1_ASAP7_75t_L g1724 ( 
.A(n_1718),
.B(n_1641),
.Y(n_1724)
);

AOI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1717),
.A2(n_1639),
.B1(n_1638),
.B2(n_1636),
.C(n_1632),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_L g1726 ( 
.A(n_1716),
.B(n_1668),
.C(n_1584),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1723),
.Y(n_1727)
);

XNOR2x1_ASAP7_75t_L g1728 ( 
.A(n_1724),
.B(n_1719),
.Y(n_1728)
);

OAI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1726),
.A2(n_1721),
.B(n_1720),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1728),
.Y(n_1730)
);

AOI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1730),
.A2(n_1722),
.B1(n_1729),
.B2(n_1725),
.Y(n_1731)
);

BUFx6f_ASAP7_75t_L g1732 ( 
.A(n_1731),
.Y(n_1732)
);

NOR3xp33_ASAP7_75t_L g1733 ( 
.A(n_1731),
.B(n_1727),
.C(n_1716),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1733),
.B(n_1579),
.Y(n_1734)
);

BUFx2_ASAP7_75t_L g1735 ( 
.A(n_1732),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1734),
.A2(n_1594),
.B1(n_1588),
.B2(n_1591),
.Y(n_1736)
);

CKINVDCx20_ASAP7_75t_R g1737 ( 
.A(n_1735),
.Y(n_1737)
);

NAND2xp33_ASAP7_75t_SL g1738 ( 
.A(n_1737),
.B(n_1734),
.Y(n_1738)
);

NAND2x1p5_ASAP7_75t_L g1739 ( 
.A(n_1738),
.B(n_1736),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1739),
.A2(n_1668),
.B(n_1642),
.Y(n_1740)
);

OAI211xp5_ASAP7_75t_L g1741 ( 
.A1(n_1740),
.A2(n_1602),
.B(n_1551),
.C(n_1554),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1741),
.A2(n_1646),
.B1(n_1611),
.B2(n_1610),
.Y(n_1742)
);

AOI211xp5_ASAP7_75t_L g1743 ( 
.A1(n_1742),
.A2(n_1551),
.B(n_1554),
.C(n_1553),
.Y(n_1743)
);


endmodule