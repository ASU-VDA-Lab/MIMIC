module fake_netlist_1_5540_n_471 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_471);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_471;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g67 ( .A(n_35), .Y(n_67) );
INVxp33_ASAP7_75t_L g68 ( .A(n_7), .Y(n_68) );
CKINVDCx5p33_ASAP7_75t_R g69 ( .A(n_33), .Y(n_69) );
CKINVDCx5p33_ASAP7_75t_R g70 ( .A(n_0), .Y(n_70) );
INVxp33_ASAP7_75t_L g71 ( .A(n_54), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_46), .Y(n_72) );
INVxp33_ASAP7_75t_L g73 ( .A(n_31), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_42), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_58), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_34), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_28), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_40), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_53), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_27), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_16), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_48), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_3), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_51), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_65), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_7), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_43), .Y(n_87) );
INVxp33_ASAP7_75t_SL g88 ( .A(n_47), .Y(n_88) );
INVxp33_ASAP7_75t_L g89 ( .A(n_14), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_19), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_20), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_49), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_41), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_14), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_10), .Y(n_95) );
CKINVDCx16_ASAP7_75t_R g96 ( .A(n_50), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_13), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_30), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_38), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_9), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_57), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_36), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_64), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_29), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_17), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_67), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_67), .Y(n_107) );
BUFx2_ASAP7_75t_L g108 ( .A(n_96), .Y(n_108) );
AND2x4_ASAP7_75t_L g109 ( .A(n_97), .B(n_0), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_82), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_82), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_72), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_70), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_74), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_100), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_74), .Y(n_117) );
BUFx8_ASAP7_75t_L g118 ( .A(n_75), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_88), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_75), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_76), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_86), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_122) );
NOR2xp33_ASAP7_75t_R g123 ( .A(n_69), .B(n_32), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_97), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_76), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_98), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_77), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_80), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_108), .B(n_71), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_111), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_108), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_127), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_118), .B(n_73), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_109), .B(n_83), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_127), .Y(n_136) );
INVx5_ASAP7_75t_L g137 ( .A(n_127), .Y(n_137) );
NAND3xp33_ASAP7_75t_L g138 ( .A(n_118), .B(n_105), .C(n_83), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_118), .B(n_129), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_127), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_111), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_127), .Y(n_142) );
INVxp67_ASAP7_75t_L g143 ( .A(n_116), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_127), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_106), .B(n_68), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_111), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_111), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_111), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_111), .Y(n_149) );
AO22x2_ASAP7_75t_L g150 ( .A1(n_109), .A2(n_113), .B1(n_125), .B2(n_106), .Y(n_150) );
INVx2_ASAP7_75t_SL g151 ( .A(n_118), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_119), .B(n_87), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_107), .B(n_89), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_128), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_109), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_128), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_154), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_145), .A2(n_126), .B1(n_109), .B2(n_114), .Y(n_159) );
NOR3xp33_ASAP7_75t_SL g160 ( .A(n_152), .B(n_81), .C(n_94), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_154), .Y(n_161) );
NOR2x1p5_ASAP7_75t_L g162 ( .A(n_130), .B(n_145), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_154), .Y(n_163) );
BUFx2_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_148), .Y(n_165) );
NOR3xp33_ASAP7_75t_SL g166 ( .A(n_134), .B(n_94), .C(n_95), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_156), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_153), .B(n_107), .Y(n_168) );
NOR3xp33_ASAP7_75t_SL g169 ( .A(n_139), .B(n_95), .C(n_101), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_135), .B(n_122), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_156), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_155), .Y(n_173) );
NAND2x1p5_ASAP7_75t_L g174 ( .A(n_155), .B(n_128), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_132), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_155), .A2(n_128), .B(n_125), .C(n_121), .Y(n_177) );
OAI22xp5_ASAP7_75t_L g178 ( .A1(n_150), .A2(n_117), .B1(n_113), .B2(n_121), .Y(n_178) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_150), .Y(n_180) );
OR2x6_ASAP7_75t_L g181 ( .A(n_150), .B(n_115), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_135), .B(n_115), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_156), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_135), .B(n_117), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_135), .B(n_112), .Y(n_185) );
NOR2xp67_ASAP7_75t_L g186 ( .A(n_143), .B(n_112), .Y(n_186) );
NOR3xp33_ASAP7_75t_SL g187 ( .A(n_138), .B(n_85), .C(n_79), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_155), .Y(n_188) );
BUFx12f_ASAP7_75t_SL g189 ( .A(n_148), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_137), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_181), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_178), .B(n_120), .Y(n_192) );
BUFx4f_ASAP7_75t_L g193 ( .A(n_181), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_182), .B(n_120), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_158), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_184), .B(n_110), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_177), .A2(n_110), .B(n_79), .C(n_84), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_157), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_179), .B(n_124), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_159), .B(n_124), .Y(n_200) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_172), .A2(n_133), .B(n_136), .Y(n_201) );
OR2x2_ASAP7_75t_L g202 ( .A(n_176), .B(n_124), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_168), .B(n_124), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_158), .Y(n_204) );
INVx3_ASAP7_75t_SL g205 ( .A(n_181), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_161), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_167), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_181), .B(n_78), .Y(n_208) );
INVxp67_ASAP7_75t_SL g209 ( .A(n_175), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_180), .B(n_78), .Y(n_210) );
INVx2_ASAP7_75t_SL g211 ( .A(n_157), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_161), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_157), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_163), .Y(n_214) );
NOR2x1_ASAP7_75t_SL g215 ( .A(n_157), .B(n_84), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_167), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_163), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_162), .B(n_92), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_170), .B(n_92), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_171), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_189), .Y(n_221) );
BUFx12f_ASAP7_75t_L g222 ( .A(n_176), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_173), .Y(n_223) );
BUFx2_ASAP7_75t_L g224 ( .A(n_164), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_157), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_203), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_193), .B(n_170), .Y(n_227) );
INVx2_ASAP7_75t_SL g228 ( .A(n_193), .Y(n_228) );
INVxp67_ASAP7_75t_L g229 ( .A(n_202), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_222), .Y(n_230) );
NOR2xp33_ASAP7_75t_SL g231 ( .A(n_193), .B(n_189), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_202), .B(n_170), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_193), .B(n_174), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_205), .Y(n_234) );
INVx4_ASAP7_75t_SL g235 ( .A(n_205), .Y(n_235) );
NAND2xp33_ASAP7_75t_SL g236 ( .A(n_205), .B(n_164), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_222), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_195), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_219), .A2(n_188), .B1(n_173), .B2(n_186), .Y(n_239) );
AND2x2_ASAP7_75t_SL g240 ( .A(n_208), .B(n_185), .Y(n_240) );
AO31x2_ASAP7_75t_L g241 ( .A1(n_192), .A2(n_147), .A3(n_149), .B(n_146), .Y(n_241) );
NOR2xp67_ASAP7_75t_L g242 ( .A(n_222), .B(n_1), .Y(n_242) );
AND2x4_ASAP7_75t_SL g243 ( .A(n_221), .B(n_166), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_224), .A2(n_188), .B1(n_160), .B2(n_169), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_195), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_191), .B(n_173), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_208), .A2(n_174), .B1(n_183), .B2(n_171), .Y(n_247) );
AOI221xp5_ASAP7_75t_L g248 ( .A1(n_200), .A2(n_187), .B1(n_183), .B2(n_174), .C(n_104), .Y(n_248) );
NAND2x1p5_ASAP7_75t_L g249 ( .A(n_191), .B(n_93), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_203), .Y(n_250) );
INVx2_ASAP7_75t_SL g251 ( .A(n_221), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_207), .B(n_190), .Y(n_252) );
CKINVDCx11_ASAP7_75t_R g253 ( .A(n_219), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_219), .A2(n_190), .B1(n_93), .B2(n_99), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_226), .B(n_207), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_246), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_253), .A2(n_219), .B1(n_218), .B2(n_224), .Y(n_257) );
INVx1_ASAP7_75t_SL g258 ( .A(n_230), .Y(n_258) );
OR2x2_ASAP7_75t_L g259 ( .A(n_232), .B(n_216), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_232), .B(n_218), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_227), .B(n_199), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_238), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_248), .A2(n_210), .B1(n_191), .B2(n_216), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_238), .Y(n_264) );
AOI211xp5_ASAP7_75t_L g265 ( .A1(n_242), .A2(n_197), .B(n_194), .C(n_196), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_233), .B(n_223), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_240), .A2(n_192), .B1(n_209), .B2(n_194), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_245), .Y(n_268) );
AOI21xp33_ASAP7_75t_L g269 ( .A1(n_244), .A2(n_196), .B(n_209), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_245), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_250), .A2(n_210), .B1(n_223), .B2(n_220), .Y(n_271) );
AOI22xp33_ASAP7_75t_SL g272 ( .A1(n_227), .A2(n_215), .B1(n_210), .B2(n_220), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_229), .A2(n_210), .B1(n_223), .B2(n_220), .C(n_217), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_252), .A2(n_223), .B1(n_206), .B2(n_217), .Y(n_274) );
OR2x2_ASAP7_75t_SL g275 ( .A(n_235), .B(n_99), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_240), .A2(n_206), .B1(n_217), .B2(n_195), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_241), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_252), .A2(n_206), .B1(n_214), .B2(n_204), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_277), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_266), .Y(n_280) );
OAI211xp5_ASAP7_75t_L g281 ( .A1(n_257), .A2(n_254), .B(n_239), .C(n_236), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_262), .Y(n_282) );
OAI222xp33_ASAP7_75t_L g283 ( .A1(n_257), .A2(n_249), .B1(n_228), .B2(n_230), .C1(n_247), .C2(n_251), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_264), .Y(n_284) );
AO22x1_ASAP7_75t_L g285 ( .A1(n_277), .A2(n_237), .B1(n_228), .B2(n_234), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_264), .Y(n_286) );
OAI21xp5_ASAP7_75t_L g287 ( .A1(n_267), .A2(n_249), .B(n_204), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_270), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_262), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g290 ( .A1(n_260), .A2(n_243), .B1(n_236), .B2(n_237), .C(n_251), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_268), .B(n_241), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_268), .B(n_241), .Y(n_292) );
OA21x2_ASAP7_75t_L g293 ( .A1(n_276), .A2(n_102), .B(n_103), .Y(n_293) );
AOI33xp33_ASAP7_75t_L g294 ( .A1(n_258), .A2(n_243), .A3(n_102), .B1(n_103), .B2(n_104), .B3(n_91), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_270), .Y(n_295) );
AND4x1_ASAP7_75t_L g296 ( .A(n_265), .B(n_231), .C(n_235), .D(n_233), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_255), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_255), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_266), .B(n_241), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_259), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_266), .B(n_241), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_291), .B(n_256), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_279), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_279), .Y(n_304) );
OAI221xp5_ASAP7_75t_L g305 ( .A1(n_290), .A2(n_263), .B1(n_272), .B2(n_261), .C(n_265), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_289), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_291), .B(n_292), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_291), .B(n_256), .Y(n_308) );
NOR3xp33_ASAP7_75t_L g309 ( .A(n_281), .B(n_269), .C(n_273), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_282), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_284), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_292), .B(n_256), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_288), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_290), .B(n_235), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_298), .B(n_275), .Y(n_315) );
OAI321xp33_ASAP7_75t_L g316 ( .A1(n_281), .A2(n_249), .A3(n_274), .B1(n_271), .B2(n_259), .C(n_278), .Y(n_316) );
NAND2x1_ASAP7_75t_SL g317 ( .A(n_292), .B(n_275), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_283), .A2(n_90), .B1(n_234), .B2(n_246), .C(n_214), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_299), .B(n_204), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_297), .B(n_246), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_299), .B(n_212), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_288), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_289), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_297), .B(n_212), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_299), .B(n_212), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_285), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_284), .Y(n_327) );
AOI33xp33_ASAP7_75t_L g328 ( .A1(n_300), .A2(n_149), .A3(n_147), .B1(n_146), .B2(n_140), .B3(n_142), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_284), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_301), .B(n_214), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_296), .B(n_235), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_301), .A2(n_225), .B1(n_211), .B2(n_198), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_310), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_306), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_306), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_307), .B(n_301), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_307), .B(n_286), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_308), .B(n_312), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_310), .B(n_300), .Y(n_339) );
AOI21xp33_ASAP7_75t_L g340 ( .A1(n_305), .A2(n_293), .B(n_280), .Y(n_340) );
NOR2xp67_ASAP7_75t_SL g341 ( .A(n_331), .B(n_293), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_326), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_323), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_323), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_308), .B(n_286), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_303), .B(n_286), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_327), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_327), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_311), .Y(n_349) );
NAND4xp25_ASAP7_75t_SL g350 ( .A(n_318), .B(n_294), .C(n_287), .D(n_296), .Y(n_350) );
OAI21x1_ASAP7_75t_SL g351 ( .A1(n_318), .A2(n_293), .B(n_295), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_305), .B(n_280), .Y(n_352) );
NOR2x1_ASAP7_75t_SL g353 ( .A(n_314), .B(n_280), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_329), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_312), .B(n_295), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_302), .B(n_288), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_329), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_320), .B(n_285), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_311), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_302), .B(n_288), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_311), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_302), .B(n_288), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_304), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_302), .B(n_288), .Y(n_364) );
CKINVDCx16_ASAP7_75t_R g365 ( .A(n_315), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_319), .B(n_288), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_319), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_321), .B(n_293), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_321), .B(n_293), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_313), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_313), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_325), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_350), .A2(n_316), .B(n_326), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_333), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_337), .Y(n_375) );
INVxp33_ASAP7_75t_L g376 ( .A(n_353), .Y(n_376) );
OAI211xp5_ASAP7_75t_SL g377 ( .A1(n_340), .A2(n_309), .B(n_328), .C(n_332), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_365), .B(n_330), .Y(n_378) );
NOR2xp33_ASAP7_75t_SL g379 ( .A(n_341), .B(n_365), .Y(n_379) );
AOI32xp33_ASAP7_75t_L g380 ( .A1(n_352), .A2(n_316), .A3(n_317), .B1(n_324), .B2(n_313), .Y(n_380) );
INVxp67_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_336), .B(n_322), .Y(n_382) );
AOI32xp33_ASAP7_75t_L g383 ( .A1(n_342), .A2(n_324), .A3(n_313), .B1(n_322), .B2(n_6), .Y(n_383) );
AOI222xp33_ASAP7_75t_L g384 ( .A1(n_353), .A2(n_215), .B1(n_4), .B2(n_5), .C1(n_6), .C2(n_8), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_338), .B(n_2), .Y(n_385) );
OAI322xp33_ASAP7_75t_L g386 ( .A1(n_363), .A2(n_4), .A3(n_5), .B1(n_8), .B2(n_9), .C1(n_10), .C2(n_11), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_338), .B(n_11), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_334), .B(n_12), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_345), .B(n_12), .Y(n_389) );
AOI211xp5_ASAP7_75t_L g390 ( .A1(n_341), .A2(n_358), .B(n_342), .C(n_368), .Y(n_390) );
OAI221xp5_ASAP7_75t_SL g391 ( .A1(n_367), .A2(n_13), .B1(n_15), .B2(n_16), .C(n_17), .Y(n_391) );
OAI21xp33_ASAP7_75t_L g392 ( .A1(n_355), .A2(n_141), .B(n_131), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_349), .Y(n_393) );
AOI211xp5_ASAP7_75t_L g394 ( .A1(n_368), .A2(n_18), .B(n_123), .C(n_148), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g395 ( .A1(n_335), .A2(n_141), .B1(n_131), .B2(n_140), .C(n_144), .Y(n_395) );
NAND3xp33_ASAP7_75t_SL g396 ( .A(n_369), .B(n_18), .C(n_141), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_349), .Y(n_397) );
AO22x1_ASAP7_75t_L g398 ( .A1(n_372), .A2(n_213), .B1(n_198), .B2(n_23), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_372), .A2(n_201), .B1(n_148), .B2(n_213), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_346), .B(n_148), .Y(n_400) );
OAI211xp5_ASAP7_75t_L g401 ( .A1(n_343), .A2(n_142), .B(n_133), .C(n_137), .Y(n_401) );
XNOR2xp5_ASAP7_75t_L g402 ( .A(n_356), .B(n_21), .Y(n_402) );
OAI22xp33_ASAP7_75t_SL g403 ( .A1(n_346), .A2(n_22), .B1(n_24), .B2(n_25), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_344), .B(n_26), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_381), .B(n_347), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_394), .A2(n_366), .B1(n_348), .B2(n_357), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_393), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_375), .B(n_348), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_374), .B(n_357), .Y(n_409) );
AOI21xp33_ASAP7_75t_L g410 ( .A1(n_384), .A2(n_354), .B(n_371), .Y(n_410) );
BUFx4f_ASAP7_75t_SL g411 ( .A(n_389), .Y(n_411) );
XNOR2xp5_ASAP7_75t_L g412 ( .A(n_402), .B(n_364), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_379), .B(n_351), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_387), .B(n_354), .Y(n_414) );
AOI21xp33_ASAP7_75t_L g415 ( .A1(n_385), .A2(n_371), .B(n_370), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_386), .A2(n_351), .B1(n_364), .B2(n_362), .C(n_360), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_386), .A2(n_370), .B1(n_361), .B2(n_359), .C(n_366), .Y(n_417) );
NAND4xp25_ASAP7_75t_SL g418 ( .A(n_383), .B(n_37), .C(n_39), .D(n_44), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_373), .A2(n_213), .B1(n_198), .B2(n_137), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_397), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_390), .B(n_213), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_382), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_378), .B(n_45), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_390), .B(n_198), .Y(n_424) );
INVx2_ASAP7_75t_SL g425 ( .A(n_400), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_388), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_404), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_376), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_426), .B(n_380), .Y(n_429) );
O2A1O1Ixp33_ASAP7_75t_L g430 ( .A1(n_424), .A2(n_403), .B(n_391), .C(n_377), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_410), .A2(n_396), .B1(n_403), .B2(n_392), .C(n_398), .Y(n_431) );
AND3x4_ASAP7_75t_L g432 ( .A(n_411), .B(n_401), .C(n_399), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_409), .Y(n_433) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_406), .A2(n_395), .B(n_137), .Y(n_434) );
OAI31xp33_ASAP7_75t_SL g435 ( .A1(n_424), .A2(n_52), .A3(n_55), .B(n_56), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_418), .A2(n_198), .B1(n_137), .B2(n_165), .Y(n_436) );
AOI32xp33_ASAP7_75t_L g437 ( .A1(n_421), .A2(n_59), .A3(n_60), .B1(n_61), .B2(n_62), .Y(n_437) );
INVxp67_ASAP7_75t_L g438 ( .A(n_405), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_411), .Y(n_439) );
INVxp67_ASAP7_75t_L g440 ( .A(n_414), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_425), .Y(n_441) );
NOR2xp33_ASAP7_75t_R g442 ( .A(n_428), .B(n_63), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_421), .A2(n_137), .B1(n_66), .B2(n_165), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_413), .A2(n_416), .B1(n_422), .B2(n_427), .Y(n_444) );
OA21x2_ASAP7_75t_L g445 ( .A1(n_415), .A2(n_165), .B(n_408), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_441), .Y(n_446) );
XNOR2xp5_ASAP7_75t_L g447 ( .A(n_439), .B(n_412), .Y(n_447) );
NAND4xp25_ASAP7_75t_L g448 ( .A(n_430), .B(n_419), .C(n_417), .D(n_423), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_440), .B(n_407), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_442), .Y(n_450) );
OR2x6_ASAP7_75t_L g451 ( .A(n_443), .B(n_420), .Y(n_451) );
XOR2x1_ASAP7_75t_L g452 ( .A(n_443), .B(n_435), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_432), .A2(n_438), .B1(n_431), .B2(n_433), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_434), .A2(n_436), .B1(n_437), .B2(n_445), .Y(n_454) );
AOI321xp33_ASAP7_75t_L g455 ( .A1(n_444), .A2(n_430), .A3(n_429), .B1(n_385), .B2(n_413), .C(n_373), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_444), .B(n_429), .Y(n_456) );
AOI22xp5_ASAP7_75t_SL g457 ( .A1(n_439), .A2(n_440), .B1(n_441), .B2(n_429), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_444), .A2(n_429), .B1(n_432), .B2(n_440), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_450), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_457), .B(n_446), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_449), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_452), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_456), .A2(n_454), .B1(n_448), .B2(n_451), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_461), .Y(n_464) );
NAND3xp33_ASAP7_75t_SL g465 ( .A(n_463), .B(n_455), .C(n_458), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_464), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_465), .B(n_462), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_466), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_467), .Y(n_469) );
OAI221xp5_ASAP7_75t_R g470 ( .A1(n_469), .A2(n_447), .B1(n_453), .B2(n_459), .C(n_460), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_470), .A2(n_460), .B(n_468), .Y(n_471) );
endmodule