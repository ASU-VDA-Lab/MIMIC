module real_aes_6906_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_1066;
wire n_684;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_1106;
wire n_778;
wire n_618;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_979;
wire n_759;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_1034;
wire n_491;
wire n_923;
wire n_894;
wire n_694;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_1137;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_932;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_638;
wire n_564;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_1160;
wire n_550;
wire n_966;
wire n_1108;
wire n_990;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_1072;
wire n_994;
wire n_1078;
wire n_384;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_931;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_1148;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_1152;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_504;
wire n_960;
wire n_455;
wire n_725;
wire n_671;
wire n_1084;
wire n_973;
wire n_1081;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1017;
wire n_1013;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_867;
wire n_722;
wire n_398;
wire n_1100;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_432;
wire n_1103;
wire n_1031;
wire n_1037;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_1041;
wire n_501;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_756;
wire n_404;
wire n_1073;
wire n_728;
wire n_598;
wire n_713;
wire n_735;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1157;
wire n_1158;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_727;
wire n_1014;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_1155;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_1136;
wire n_720;
wire n_1127;
wire n_968;
wire n_435;
wire n_972;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_928;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1052;
wire n_787;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_1090;
wire n_456;
wire n_717;
wire n_982;
wire n_1133;
wire n_1164;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_1162;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_929;
wire n_1143;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_1045;
wire n_566;
wire n_719;
wire n_837;
wire n_1114;
wire n_871;
wire n_967;
wire n_474;
wire n_1156;
wire n_1159;
wire n_829;
wire n_1030;
wire n_988;
wire n_1088;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1151;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_1040;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_1097;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1101;
wire n_447;
wire n_1102;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_1039;
wire n_1119;
wire n_802;
wire n_868;
wire n_877;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_0), .A2(n_286), .B1(n_528), .B2(n_529), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_1), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g1072 ( .A(n_2), .Y(n_1072) );
CKINVDCx20_ASAP7_75t_R g888 ( .A(n_3), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_4), .A2(n_51), .B1(n_726), .B2(n_728), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g1018 ( .A(n_5), .Y(n_1018) );
AOI221xp5_ASAP7_75t_L g753 ( .A1(n_6), .A2(n_14), .B1(n_511), .B2(n_754), .C(n_756), .Y(n_753) );
AOI221xp5_ASAP7_75t_L g735 ( .A1(n_7), .A2(n_270), .B1(n_692), .B2(n_736), .C(n_738), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_8), .A2(n_140), .B1(n_688), .B2(n_844), .Y(n_843) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_9), .Y(n_416) );
AO22x2_ASAP7_75t_L g405 ( .A1(n_10), .A2(n_220), .B1(n_406), .B2(n_407), .Y(n_405) );
INVx1_ASAP7_75t_L g1104 ( .A(n_10), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_11), .A2(n_160), .B1(n_531), .B2(n_634), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_12), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g924 ( .A(n_13), .Y(n_924) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_15), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_16), .A2(n_288), .B1(n_608), .B2(n_609), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_17), .A2(n_106), .B1(n_634), .B2(n_911), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_18), .A2(n_54), .B1(n_549), .B2(n_550), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g1030 ( .A(n_19), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_20), .A2(n_244), .B1(n_638), .B2(n_639), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_21), .B(n_653), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g896 ( .A(n_22), .Y(n_896) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_23), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_24), .A2(n_358), .B1(n_489), .B2(n_591), .Y(n_590) );
CKINVDCx20_ASAP7_75t_R g1006 ( .A(n_25), .Y(n_1006) );
AOI222xp33_ASAP7_75t_L g623 ( .A1(n_26), .A2(n_56), .B1(n_340), .B2(n_504), .C1(n_575), .C2(n_624), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g1038 ( .A(n_27), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_28), .A2(n_124), .B1(n_461), .B2(n_465), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_29), .A2(n_55), .B1(n_488), .B2(n_913), .Y(n_983) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_30), .Y(n_870) );
AO22x2_ASAP7_75t_L g409 ( .A1(n_31), .A2(n_112), .B1(n_406), .B2(n_410), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_32), .A2(n_734), .B1(n_760), .B2(n_761), .Y(n_733) );
INVx1_ASAP7_75t_L g760 ( .A(n_32), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_33), .A2(n_372), .B1(n_479), .B2(n_482), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g1009 ( .A1(n_34), .A2(n_1010), .B1(n_1040), .B2(n_1041), .Y(n_1009) );
CKINVDCx20_ASAP7_75t_R g1040 ( .A(n_34), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_35), .A2(n_245), .B1(n_465), .B2(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g1118 ( .A(n_36), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_37), .A2(n_116), .B1(n_524), .B2(n_525), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_38), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_39), .A2(n_63), .B1(n_844), .B2(n_916), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_40), .A2(n_163), .B1(n_706), .B2(n_707), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g994 ( .A1(n_41), .A2(n_275), .B1(n_470), .B2(n_844), .Y(n_994) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_42), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_43), .B(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_44), .B(n_418), .Y(n_976) );
CKINVDCx20_ASAP7_75t_R g979 ( .A(n_45), .Y(n_979) );
CKINVDCx20_ASAP7_75t_R g978 ( .A(n_46), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_47), .A2(n_190), .B1(n_619), .B2(n_634), .Y(n_1013) );
AOI22xp5_ASAP7_75t_L g1007 ( .A1(n_48), .A2(n_214), .B1(n_450), .B2(n_625), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_49), .A2(n_331), .B1(n_589), .B2(n_772), .Y(n_1125) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_50), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g975 ( .A(n_52), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_53), .A2(n_125), .B1(n_916), .B2(n_917), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_57), .A2(n_147), .B1(n_540), .B2(n_642), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_58), .A2(n_243), .B1(n_638), .B2(n_639), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_59), .A2(n_285), .B1(n_594), .B2(n_597), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_60), .B(n_653), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_61), .A2(n_312), .B1(n_540), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_62), .A2(n_109), .B1(n_689), .B2(n_769), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_64), .A2(n_827), .B1(n_850), .B2(n_851), .Y(n_826) );
INVx1_ASAP7_75t_L g850 ( .A(n_64), .Y(n_850) );
AOI22xp33_ASAP7_75t_SL g1059 ( .A1(n_65), .A2(n_273), .B1(n_541), .B2(n_543), .Y(n_1059) );
CKINVDCx20_ASAP7_75t_R g1075 ( .A(n_66), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_67), .A2(n_342), .B1(n_638), .B2(n_639), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_68), .A2(n_295), .B1(n_594), .B2(n_1127), .Y(n_1126) );
CKINVDCx20_ASAP7_75t_R g1112 ( .A(n_69), .Y(n_1112) );
INVx1_ASAP7_75t_L g946 ( .A(n_70), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_71), .A2(n_356), .B1(n_539), .B2(n_540), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g1023 ( .A(n_72), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_73), .A2(n_104), .B1(n_402), .B2(n_465), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_74), .A2(n_339), .B1(n_540), .B2(n_846), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_75), .A2(n_100), .B1(n_591), .B2(n_876), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_76), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_77), .B(n_728), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_78), .A2(n_289), .B1(n_621), .B2(n_622), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g930 ( .A(n_79), .Y(n_930) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_80), .A2(n_210), .B1(n_503), .B2(n_504), .Y(n_502) );
INVx1_ASAP7_75t_L g991 ( .A(n_81), .Y(n_991) );
CKINVDCx20_ASAP7_75t_R g1032 ( .A(n_82), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_83), .A2(n_186), .B1(n_709), .B2(n_1160), .Y(n_1159) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_84), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_85), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_86), .A2(n_208), .B1(n_554), .B2(n_688), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_87), .A2(n_133), .B1(n_546), .B2(n_547), .Y(n_731) );
AO22x2_ASAP7_75t_L g415 ( .A1(n_88), .A2(n_250), .B1(n_406), .B2(n_407), .Y(n_415) );
INVx1_ASAP7_75t_L g1101 ( .A(n_88), .Y(n_1101) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_89), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_90), .A2(n_91), .B1(n_608), .B2(n_622), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_92), .A2(n_230), .B1(n_531), .B2(n_634), .Y(n_1158) );
AOI22xp5_ASAP7_75t_L g997 ( .A1(n_93), .A2(n_110), .B1(n_640), .B2(n_880), .Y(n_997) );
AOI22xp5_ASAP7_75t_L g892 ( .A1(n_94), .A2(n_225), .B1(n_419), .B2(n_800), .Y(n_892) );
AOI22x1_ASAP7_75t_L g965 ( .A1(n_95), .A2(n_966), .B1(n_987), .B2(n_988), .Y(n_965) );
INVx1_ASAP7_75t_L g987 ( .A(n_95), .Y(n_987) );
CKINVDCx20_ASAP7_75t_R g1145 ( .A(n_96), .Y(n_1145) );
AOI222xp33_ASAP7_75t_L g759 ( .A1(n_97), .A2(n_107), .B1(n_138), .B2(n_549), .C1(n_575), .C2(n_624), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_98), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_99), .A2(n_254), .B1(n_525), .B2(n_772), .Y(n_1155) );
INVx1_ASAP7_75t_L g657 ( .A(n_101), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g1076 ( .A(n_102), .Y(n_1076) );
CKINVDCx20_ASAP7_75t_R g1070 ( .A(n_103), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_105), .A2(n_183), .B1(n_615), .B2(n_616), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_108), .A2(n_363), .B1(n_473), .B2(n_556), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g969 ( .A(n_111), .Y(n_969) );
INVx1_ASAP7_75t_L g1105 ( .A(n_112), .Y(n_1105) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_113), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g1001 ( .A(n_114), .Y(n_1001) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_115), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_117), .A2(n_215), .B1(n_482), .B2(n_543), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g891 ( .A(n_118), .Y(n_891) );
CKINVDCx20_ASAP7_75t_R g1029 ( .A(n_119), .Y(n_1029) );
CKINVDCx20_ASAP7_75t_R g1048 ( .A(n_120), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_121), .B(n_653), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_122), .A2(n_290), .B1(n_461), .B2(n_634), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_123), .A2(n_135), .B1(n_554), .B2(n_692), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g899 ( .A1(n_126), .A2(n_301), .B1(n_463), .B2(n_465), .Y(n_899) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_127), .Y(n_423) );
AOI22xp33_ASAP7_75t_SL g807 ( .A1(n_128), .A2(n_178), .B1(n_677), .B2(n_808), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_129), .A2(n_209), .B1(n_846), .B2(n_920), .Y(n_919) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_130), .A2(n_296), .B1(n_489), .B2(n_608), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g1152 ( .A(n_131), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_132), .A2(n_330), .B1(n_419), .B2(n_808), .Y(n_1073) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_134), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_136), .A2(n_303), .B1(n_450), .B2(n_579), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g1055 ( .A1(n_137), .A2(n_321), .B1(n_616), .B2(n_800), .Y(n_1055) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_139), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_141), .A2(n_326), .B1(n_539), .B2(n_605), .Y(n_604) );
AOI222xp33_ASAP7_75t_L g557 ( .A1(n_142), .A2(n_222), .B1(n_306), .B2(n_403), .C1(n_427), .C2(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_143), .A2(n_196), .B1(n_522), .B2(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_144), .A2(n_201), .B1(n_531), .B2(n_533), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g1000 ( .A(n_145), .Y(n_1000) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_146), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g1144 ( .A(n_148), .Y(n_1144) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_149), .B(n_1052), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_150), .A2(n_200), .B1(n_470), .B2(n_473), .Y(n_469) );
AND2x6_ASAP7_75t_L g385 ( .A(n_151), .B(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g1098 ( .A(n_151), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_152), .A2(n_237), .B1(n_688), .B2(n_689), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_153), .A2(n_276), .B1(n_425), .B2(n_550), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_154), .A2(n_176), .B1(n_483), .B2(n_621), .Y(n_1082) );
INVx1_ASAP7_75t_L g684 ( .A(n_155), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_156), .A2(n_263), .B1(n_650), .B2(n_880), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_157), .A2(n_278), .B1(n_482), .B2(n_642), .Y(n_986) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_158), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_159), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_161), .A2(n_185), .B1(n_520), .B2(n_522), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g1107 ( .A1(n_162), .A2(n_1108), .B1(n_1128), .B2(n_1129), .Y(n_1107) );
CKINVDCx20_ASAP7_75t_R g1128 ( .A(n_162), .Y(n_1128) );
AOI22xp5_ASAP7_75t_SL g938 ( .A1(n_164), .A2(n_939), .B1(n_959), .B2(n_960), .Y(n_938) );
INVx1_ASAP7_75t_L g960 ( .A(n_164), .Y(n_960) );
AOI22xp33_ASAP7_75t_SL g1049 ( .A1(n_165), .A2(n_280), .B1(n_514), .B2(n_625), .Y(n_1049) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_166), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g995 ( .A1(n_167), .A2(n_300), .B1(n_483), .B2(n_533), .Y(n_995) );
NAND2xp5_ASAP7_75t_SL g804 ( .A(n_168), .B(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g942 ( .A(n_169), .Y(n_942) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_170), .Y(n_786) );
AO22x2_ASAP7_75t_L g413 ( .A1(n_171), .A2(n_241), .B1(n_406), .B2(n_410), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g1102 ( .A(n_171), .B(n_1103), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_172), .A2(n_181), .B1(n_605), .B2(n_642), .Y(n_1123) );
AOI22xp33_ASAP7_75t_SL g814 ( .A1(n_173), .A2(n_258), .B1(n_707), .B2(n_815), .Y(n_814) );
XNOR2x2_ASAP7_75t_L g535 ( .A(n_174), .B(n_536), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_175), .A2(n_357), .B1(n_594), .B2(n_597), .Y(n_593) );
AOI22xp33_ASAP7_75t_SL g799 ( .A1(n_177), .A2(n_268), .B1(n_503), .B2(n_800), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g973 ( .A(n_179), .Y(n_973) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_180), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_182), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_184), .A2(n_316), .B1(n_531), .B2(n_543), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_187), .Y(n_886) );
AOI22xp33_ASAP7_75t_SL g813 ( .A1(n_188), .A2(n_199), .B1(n_554), .B2(n_640), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g998 ( .A1(n_189), .A2(n_228), .B1(n_608), .B2(n_901), .Y(n_998) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_191), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_192), .A2(n_310), .B1(n_482), .B2(n_642), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_193), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_194), .B(n_1036), .Y(n_1035) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_195), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_197), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_198), .A2(n_366), .B1(n_608), .B2(n_609), .Y(n_607) );
AOI22xp33_ASAP7_75t_SL g810 ( .A1(n_202), .A2(n_355), .B1(n_479), .B2(n_605), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_203), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_204), .B(n_653), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_205), .Y(n_432) );
AOI22xp33_ASAP7_75t_SL g1058 ( .A1(n_206), .A2(n_255), .B1(n_465), .B2(n_621), .Y(n_1058) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_207), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_211), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_212), .A2(n_219), .B1(n_503), .B2(n_867), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_213), .A2(n_327), .B1(n_463), .B2(n_556), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_216), .A2(n_253), .B1(n_554), .B2(n_622), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_217), .A2(n_223), .B1(n_528), .B2(n_772), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_218), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_221), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_224), .A2(n_347), .B1(n_690), .B2(n_957), .Y(n_956) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_226), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_227), .A2(n_272), .B1(n_916), .B2(n_917), .Y(n_958) );
OA22x2_ASAP7_75t_L g1064 ( .A1(n_229), .A2(n_1065), .B1(n_1066), .B2(n_1084), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_229), .Y(n_1065) );
CKINVDCx20_ASAP7_75t_R g1148 ( .A(n_231), .Y(n_1148) );
CKINVDCx20_ASAP7_75t_R g926 ( .A(n_232), .Y(n_926) );
CKINVDCx20_ASAP7_75t_R g970 ( .A(n_233), .Y(n_970) );
CKINVDCx20_ASAP7_75t_R g1039 ( .A(n_234), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_235), .B(n_803), .Y(n_802) );
XNOR2x2_ASAP7_75t_L g701 ( .A(n_236), .B(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g390 ( .A(n_238), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_239), .A2(n_630), .B1(n_660), .B2(n_661), .Y(n_629) );
INVx1_ASAP7_75t_L g660 ( .A(n_239), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g931 ( .A(n_240), .Y(n_931) );
AOI22xp5_ASAP7_75t_L g878 ( .A1(n_242), .A2(n_252), .B1(n_461), .B2(n_594), .Y(n_878) );
AOI22xp33_ASAP7_75t_SL g1062 ( .A1(n_246), .A2(n_375), .B1(n_488), .B2(n_901), .Y(n_1062) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_247), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g1061 ( .A1(n_248), .A2(n_369), .B1(n_589), .B2(n_844), .Y(n_1061) );
CKINVDCx20_ASAP7_75t_R g1147 ( .A(n_249), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_251), .A2(n_348), .B1(n_514), .B2(n_515), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g1020 ( .A(n_256), .Y(n_1020) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_257), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g1034 ( .A(n_259), .Y(n_1034) );
CKINVDCx20_ASAP7_75t_R g1139 ( .A(n_260), .Y(n_1139) );
AOI22xp5_ASAP7_75t_L g1140 ( .A1(n_260), .A2(n_1139), .B1(n_1141), .B2(n_1161), .Y(n_1140) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_261), .A2(n_764), .B1(n_790), .B2(n_791), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_261), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_262), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_264), .A2(n_298), .B1(n_481), .B2(n_639), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_265), .A2(n_364), .B1(n_605), .B2(n_846), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_266), .B(n_507), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_267), .A2(n_371), .B1(n_473), .B2(n_815), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_269), .A2(n_352), .B1(n_709), .B2(n_1015), .Y(n_1014) );
CKINVDCx20_ASAP7_75t_R g1069 ( .A(n_271), .Y(n_1069) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_274), .A2(n_383), .B(n_391), .C(n_1106), .Y(n_382) );
INVx1_ASAP7_75t_L g945 ( .A(n_277), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_279), .A2(n_297), .B1(n_487), .B2(n_489), .Y(n_486) );
INVx1_ASAP7_75t_L g949 ( .A(n_281), .Y(n_949) );
INVx1_ASAP7_75t_L g406 ( .A(n_282), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_282), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_283), .A2(n_368), .B1(n_465), .B2(n_880), .Y(n_879) );
CKINVDCx20_ASAP7_75t_R g927 ( .A(n_284), .Y(n_927) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_287), .Y(n_894) );
AOI221xp5_ASAP7_75t_L g744 ( .A1(n_291), .A2(n_305), .B1(n_594), .B2(n_745), .C(n_748), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_292), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_293), .Y(n_493) );
INVx1_ASAP7_75t_L g645 ( .A(n_294), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_299), .B(n_507), .Y(n_613) );
AOI22xp33_ASAP7_75t_SL g527 ( .A1(n_302), .A2(n_361), .B1(n_528), .B2(n_529), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_304), .A2(n_325), .B1(n_463), .B2(n_634), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_307), .A2(n_354), .B1(n_621), .B2(n_901), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_308), .A2(n_338), .B1(n_427), .B2(n_515), .Y(n_1002) );
CKINVDCx20_ASAP7_75t_R g1115 ( .A(n_309), .Y(n_1115) );
INVx1_ASAP7_75t_L g389 ( .A(n_311), .Y(n_389) );
INVx1_ASAP7_75t_L g1119 ( .A(n_313), .Y(n_1119) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_314), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_315), .B(n_728), .Y(n_1149) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_317), .Y(n_816) );
INVx1_ASAP7_75t_L g386 ( .A(n_318), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_319), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_320), .Y(n_749) );
OA22x2_ASAP7_75t_L g1043 ( .A1(n_322), .A2(n_1044), .B1(n_1045), .B2(n_1063), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_322), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_323), .A2(n_360), .B1(n_622), .B2(n_688), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_324), .B(n_806), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_328), .A2(n_341), .B1(n_522), .B2(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_329), .A2(n_332), .B1(n_546), .B2(n_547), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_333), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_334), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g1025 ( .A(n_335), .Y(n_1025) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_336), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_337), .B(n_728), .Y(n_947) );
CKINVDCx20_ASAP7_75t_R g1151 ( .A(n_343), .Y(n_1151) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_344), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g678 ( .A(n_345), .Y(n_678) );
INVx1_ASAP7_75t_L g881 ( .A(n_346), .Y(n_881) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_349), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_350), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g943 ( .A(n_351), .Y(n_943) );
CKINVDCx20_ASAP7_75t_R g869 ( .A(n_353), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_359), .Y(n_782) );
INVx1_ASAP7_75t_L g905 ( .A(n_362), .Y(n_905) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_365), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_367), .B(n_503), .Y(n_1116) );
CKINVDCx20_ASAP7_75t_R g923 ( .A(n_370), .Y(n_923) );
OA22x2_ASAP7_75t_SL g665 ( .A1(n_373), .A2(n_666), .B1(n_667), .B2(n_696), .Y(n_665) );
INVx1_ASAP7_75t_L g696 ( .A(n_373), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g906 ( .A1(n_374), .A2(n_907), .B1(n_932), .B2(n_933), .Y(n_906) );
INVx1_ASAP7_75t_L g932 ( .A(n_374), .Y(n_932) );
CKINVDCx20_ASAP7_75t_R g1111 ( .A(n_376), .Y(n_1111) );
CKINVDCx20_ASAP7_75t_R g839 ( .A(n_377), .Y(n_839) );
INVx1_ASAP7_75t_L g950 ( .A(n_378), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_379), .A2(n_381), .B1(n_531), .B2(n_913), .Y(n_912) );
CKINVDCx20_ASAP7_75t_R g1114 ( .A(n_380), .Y(n_1114) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_385), .B(n_387), .Y(n_384) );
HB1xp67_ASAP7_75t_L g1097 ( .A(n_386), .Y(n_1097) );
OA21x2_ASAP7_75t_L g1137 ( .A1(n_387), .A2(n_1096), .B(n_1138), .Y(n_1137) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_823), .B1(n_1091), .B2(n_1092), .C(n_1093), .Y(n_391) );
INVxp67_ASAP7_75t_L g1091 ( .A(n_392), .Y(n_1091) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_699), .B1(n_700), .B2(n_822), .Y(n_392) );
INVx1_ASAP7_75t_L g822 ( .A(n_393), .Y(n_822) );
XOR2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_561), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_494), .B2(n_495), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
XOR2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_493), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_458), .Y(n_398) );
NOR3xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_431), .C(n_447), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_416), .B1(n_417), .B2(n_423), .C(n_424), .Y(n_400) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_401), .A2(n_501), .B(n_502), .Y(n_500) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_SL g972 ( .A(n_402), .Y(n_972) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx4_ASAP7_75t_L g576 ( .A(n_403), .Y(n_576) );
INVx2_ASAP7_75t_L g723 ( .A(n_403), .Y(n_723) );
INVx2_ASAP7_75t_L g781 ( .A(n_403), .Y(n_781) );
BUFx3_ASAP7_75t_L g1005 ( .A(n_403), .Y(n_1005) );
AND2x6_ASAP7_75t_L g403 ( .A(n_404), .B(n_411), .Y(n_403) );
AND2x4_ASAP7_75t_L g428 ( .A(n_404), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g584 ( .A(n_404), .Y(n_584) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_409), .Y(n_404) );
AND2x2_ASAP7_75t_L g422 ( .A(n_405), .B(n_413), .Y(n_422) );
INVx2_ASAP7_75t_L g438 ( .A(n_405), .Y(n_438) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_408), .Y(n_410) );
OR2x2_ASAP7_75t_L g437 ( .A(n_409), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g446 ( .A(n_409), .B(n_438), .Y(n_446) );
INVx2_ASAP7_75t_L g453 ( .A(n_409), .Y(n_453) );
INVx1_ASAP7_75t_L g492 ( .A(n_409), .Y(n_492) );
AND2x6_ASAP7_75t_L g463 ( .A(n_411), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g472 ( .A(n_411), .B(n_468), .Y(n_472) );
AND2x4_ASAP7_75t_L g481 ( .A(n_411), .B(n_446), .Y(n_481) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_414), .Y(n_411) );
AND2x2_ASAP7_75t_L g440 ( .A(n_412), .B(n_415), .Y(n_440) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g467 ( .A(n_413), .B(n_430), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_413), .B(n_415), .Y(n_476) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g421 ( .A(n_415), .Y(n_421) );
INVx1_ASAP7_75t_L g430 ( .A(n_415), .Y(n_430) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx4f_ASAP7_75t_L g728 ( .A(n_418), .Y(n_728) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_419), .Y(n_503) );
BUFx12f_ASAP7_75t_L g625 ( .A(n_419), .Y(n_625) );
AND2x4_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g452 ( .A(n_421), .B(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g451 ( .A(n_422), .B(n_452), .Y(n_451) );
NAND2x1p5_ASAP7_75t_L g456 ( .A(n_422), .B(n_457), .Y(n_456) );
AND2x4_ASAP7_75t_L g515 ( .A(n_422), .B(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_SL g504 ( .A(n_428), .Y(n_504) );
BUFx2_ASAP7_75t_SL g800 ( .A(n_428), .Y(n_800) );
INVx1_ASAP7_75t_L g585 ( .A(n_429), .Y(n_585) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B1(n_441), .B2(n_442), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_433), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_568) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_435), .A2(n_444), .B1(n_645), .B2(n_646), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_435), .A2(n_612), .B1(n_923), .B2(n_924), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_435), .A2(n_571), .B1(n_1038), .B2(n_1039), .Y(n_1037) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g672 ( .A(n_436), .Y(n_672) );
BUFx3_ASAP7_75t_L g887 ( .A(n_436), .Y(n_887) );
OAI221xp5_ASAP7_75t_L g999 ( .A1(n_436), .A2(n_444), .B1(n_1000), .B2(n_1001), .C(n_1002), .Y(n_999) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
INVx2_ASAP7_75t_L g464 ( .A(n_437), .Y(n_464) );
AND2x2_ASAP7_75t_L g468 ( .A(n_438), .B(n_453), .Y(n_468) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2x1p5_ASAP7_75t_L g445 ( .A(n_440), .B(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_L g488 ( .A(n_440), .B(n_468), .Y(n_488) );
AND2x4_ASAP7_75t_L g509 ( .A(n_440), .B(n_464), .Y(n_509) );
AND2x6_ASAP7_75t_L g512 ( .A(n_440), .B(n_446), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_442), .A2(n_670), .B1(n_671), .B2(n_673), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_442), .A2(n_830), .B1(n_831), .B2(n_832), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_442), .A2(n_787), .B1(n_861), .B2(n_862), .Y(n_860) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_442), .A2(n_887), .B1(n_1111), .B2(n_1112), .Y(n_1110) );
OAI22xp5_ASAP7_75t_L g1143 ( .A1(n_442), .A2(n_831), .B1(n_1144), .B2(n_1145), .Y(n_1143) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx3_ASAP7_75t_L g789 ( .A(n_444), .Y(n_789) );
BUFx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g572 ( .A(n_445), .Y(n_572) );
AND2x2_ASAP7_75t_L g485 ( .A(n_446), .B(n_467), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_446), .B(n_467), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B1(n_454), .B2(n_455), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_450), .Y(n_549) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx4f_ASAP7_75t_SL g514 ( .A(n_451), .Y(n_514) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_451), .Y(n_615) );
BUFx2_ASAP7_75t_L g650 ( .A(n_451), .Y(n_650) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_451), .Y(n_677) );
INVx1_ASAP7_75t_L g457 ( .A(n_453), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_455), .A2(n_582), .B1(n_930), .B2(n_931), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_455), .A2(n_582), .B1(n_978), .B2(n_979), .Y(n_977) );
BUFx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_456), .Y(n_656) );
INVx4_ASAP7_75t_L g683 ( .A(n_456), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g893 ( .A1(n_456), .A2(n_894), .B1(n_895), .B2(n_896), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_456), .A2(n_871), .B1(n_949), .B2(n_950), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_456), .A2(n_871), .B1(n_1029), .B2(n_1030), .Y(n_1028) );
AND2x2_ASAP7_75t_L g533 ( .A(n_457), .B(n_475), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_477), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_469), .Y(n_459) );
INVx2_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVx4_ASAP7_75t_L g554 ( .A(n_462), .Y(n_554) );
INVx4_ASAP7_75t_L g844 ( .A(n_462), .Y(n_844) );
OAI21xp33_ASAP7_75t_SL g1071 ( .A1(n_462), .A2(n_1072), .B(n_1073), .Y(n_1071) );
INVx11_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx11_ASAP7_75t_L g521 ( .A(n_463), .Y(n_521) );
INVx1_ASAP7_75t_L g773 ( .A(n_465), .Y(n_773) );
BUFx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx3_ASAP7_75t_L g522 ( .A(n_466), .Y(n_522) );
BUFx3_ASAP7_75t_L g640 ( .A(n_466), .Y(n_640) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_467), .B(n_468), .Y(n_720) );
AND2x4_ASAP7_75t_L g474 ( .A(n_468), .B(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx3_ASAP7_75t_L g621 ( .A(n_471), .Y(n_621) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_472), .Y(n_524) );
BUFx2_ASAP7_75t_SL g556 ( .A(n_472), .Y(n_556) );
BUFx2_ASAP7_75t_SL g815 ( .A(n_472), .Y(n_815) );
BUFx2_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g525 ( .A(n_474), .Y(n_525) );
BUFx3_ASAP7_75t_L g622 ( .A(n_474), .Y(n_622) );
BUFx3_ASAP7_75t_L g692 ( .A(n_474), .Y(n_692) );
BUFx2_ASAP7_75t_SL g707 ( .A(n_474), .Y(n_707) );
BUFx3_ASAP7_75t_L g769 ( .A(n_474), .Y(n_769) );
BUFx2_ASAP7_75t_L g901 ( .A(n_474), .Y(n_901) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OR2x6_ASAP7_75t_L g491 ( .A(n_476), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_486), .Y(n_477) );
INVx2_ASAP7_75t_L g1019 ( .A(n_479), .Y(n_1019) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g528 ( .A(n_480), .Y(n_528) );
INVx2_ASAP7_75t_L g539 ( .A(n_480), .Y(n_539) );
INVx3_ASAP7_75t_L g589 ( .A(n_480), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_480), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_715) );
INVx6_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx3_ASAP7_75t_L g638 ( .A(n_481), .Y(n_638) );
BUFx3_ASAP7_75t_L g751 ( .A(n_481), .Y(n_751) );
BUFx3_ASAP7_75t_L g880 ( .A(n_481), .Y(n_880) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_L g1160 ( .A(n_483), .Y(n_1160) );
INVx5_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx3_ASAP7_75t_L g529 ( .A(n_484), .Y(n_529) );
INVx4_ASAP7_75t_L g541 ( .A(n_484), .Y(n_541) );
BUFx3_ASAP7_75t_L g606 ( .A(n_484), .Y(n_606) );
INVx2_ASAP7_75t_L g920 ( .A(n_484), .Y(n_920) );
INVx1_ASAP7_75t_L g1016 ( .A(n_484), .Y(n_1016) );
INVx8_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g532 ( .A(n_488), .Y(n_532) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_488), .Y(n_596) );
BUFx3_ASAP7_75t_L g608 ( .A(n_488), .Y(n_608) );
BUFx3_ASAP7_75t_L g690 ( .A(n_488), .Y(n_690) );
BUFx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_L g609 ( .A(n_490), .Y(n_609) );
BUFx4f_ASAP7_75t_SL g642 ( .A(n_490), .Y(n_642) );
BUFx2_ASAP7_75t_L g709 ( .A(n_490), .Y(n_709) );
BUFx2_ASAP7_75t_L g846 ( .A(n_490), .Y(n_846) );
INVx6_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_SL g543 ( .A(n_491), .Y(n_543) );
INVx1_ASAP7_75t_L g876 ( .A(n_491), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_491), .A2(n_583), .B1(n_1075), .B2(n_1076), .Y(n_1074) );
INVx1_ASAP7_75t_L g516 ( .A(n_492), .Y(n_516) );
INVx1_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B1(n_535), .B2(n_560), .Y(n_495) );
OAI22xp5_ASAP7_75t_SL g663 ( .A1(n_496), .A2(n_664), .B1(n_665), .B2(n_697), .Y(n_663) );
INVx2_ASAP7_75t_SL g697 ( .A(n_496), .Y(n_697) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
XOR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_534), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_499), .B(n_517), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_505), .Y(n_499) );
INVx2_ASAP7_75t_L g559 ( .A(n_503), .Y(n_559) );
BUFx3_ASAP7_75t_L g653 ( .A(n_503), .Y(n_653) );
BUFx2_ASAP7_75t_L g1036 ( .A(n_503), .Y(n_1036) );
NAND3xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_510), .C(n_513), .Y(n_505) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g546 ( .A(n_508), .Y(n_546) );
INVx2_ASAP7_75t_L g755 ( .A(n_508), .Y(n_755) );
INVx5_ASAP7_75t_L g806 ( .A(n_508), .Y(n_806) );
INVx4_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx4f_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx2_ASAP7_75t_L g547 ( .A(n_512), .Y(n_547) );
BUFx2_ASAP7_75t_L g803 ( .A(n_512), .Y(n_803) );
INVx1_ASAP7_75t_SL g1053 ( .A(n_512), .Y(n_1053) );
INVx1_ASAP7_75t_L g974 ( .A(n_514), .Y(n_974) );
INVx1_ASAP7_75t_L g551 ( .A(n_515), .Y(n_551) );
BUFx2_ASAP7_75t_L g579 ( .A(n_515), .Y(n_579) );
BUFx3_ASAP7_75t_L g616 ( .A(n_515), .Y(n_616) );
BUFx2_ASAP7_75t_L g808 ( .A(n_515), .Y(n_808) );
NOR2x1_ASAP7_75t_L g517 ( .A(n_518), .B(n_526), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
INVx4_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g619 ( .A(n_521), .Y(n_619) );
INVx5_ASAP7_75t_SL g713 ( .A(n_521), .Y(n_713) );
INVx2_ASAP7_75t_SL g747 ( .A(n_521), .Y(n_747) );
INVx2_ASAP7_75t_L g957 ( .A(n_521), .Y(n_957) );
INVx1_ASAP7_75t_L g918 ( .A(n_522), .Y(n_918) );
BUFx3_ASAP7_75t_L g634 ( .A(n_524), .Y(n_634) );
BUFx3_ASAP7_75t_L g688 ( .A(n_524), .Y(n_688) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_524), .Y(n_706) );
INVx3_ASAP7_75t_L g737 ( .A(n_524), .Y(n_737) );
INVx2_ASAP7_75t_L g598 ( .A(n_525), .Y(n_598) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_525), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_530), .Y(n_526) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g560 ( .A(n_535), .Y(n_560) );
NAND4xp75_ASAP7_75t_L g536 ( .A(n_537), .B(n_544), .C(n_552), .D(n_557), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_542), .Y(n_537) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g592 ( .A(n_541), .Y(n_592) );
AND2x2_ASAP7_75t_SL g544 ( .A(n_545), .B(n_548), .Y(n_544) );
INVx2_ASAP7_75t_SL g895 ( .A(n_549), .Y(n_895) );
INVx2_ASAP7_75t_SL g1033 ( .A(n_549), .Y(n_1033) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OAI22xp5_ASAP7_75t_SL g580 ( .A1(n_559), .A2(n_581), .B1(n_582), .B2(n_586), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B1(n_627), .B2(n_698), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
XNOR2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_600), .Y(n_563) );
XNOR2x1_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_587), .Y(n_566) );
NOR3xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_573), .C(n_580), .Y(n_567) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_SL g612 ( .A(n_572), .Y(n_612) );
INVx1_ASAP7_75t_L g889 ( .A(n_572), .Y(n_889) );
OAI21xp33_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_577), .B(n_578), .Y(n_573) );
OAI221xp5_ASAP7_75t_SL g647 ( .A1(n_574), .A2(n_648), .B1(n_649), .B2(n_651), .C(n_652), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_574), .A2(n_675), .B1(n_676), .B2(n_678), .C(n_679), .Y(n_674) );
OAI221xp5_ASAP7_75t_SL g833 ( .A1(n_574), .A2(n_834), .B1(n_835), .B2(n_836), .C(n_837), .Y(n_833) );
OAI221xp5_ASAP7_75t_L g925 ( .A1(n_574), .A2(n_676), .B1(n_926), .B2(n_927), .C(n_928), .Y(n_925) );
OAI221xp5_ASAP7_75t_SL g944 ( .A1(n_574), .A2(n_649), .B1(n_945), .B2(n_946), .C(n_947), .Y(n_944) );
OAI221xp5_ASAP7_75t_L g1031 ( .A1(n_574), .A2(n_1032), .B1(n_1033), .B2(n_1034), .C(n_1035), .Y(n_1031) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx4_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
BUFx2_ASAP7_75t_L g865 ( .A(n_576), .Y(n_865) );
OAI21xp5_ASAP7_75t_SL g890 ( .A1(n_576), .A2(n_891), .B(n_892), .Y(n_890) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_582), .A2(n_681), .B1(n_682), .B2(n_684), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g1117 ( .A1(n_582), .A2(n_778), .B1(n_1118), .B2(n_1119), .Y(n_1117) );
BUFx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
CKINVDCx16_ASAP7_75t_R g659 ( .A(n_583), .Y(n_659) );
OR2x6_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
AND4x1_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .C(n_593), .D(n_599), .Y(n_587) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx4_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_595), .A2(n_711), .B1(n_712), .B2(n_714), .Y(n_710) );
INVx4_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
XNOR2x2_ASAP7_75t_L g793 ( .A(n_601), .B(n_794), .Y(n_793) );
XOR2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_626), .Y(n_601) );
NAND4xp75_ASAP7_75t_L g602 ( .A(n_603), .B(n_610), .C(n_617), .D(n_623), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_607), .Y(n_603) );
INVx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OA211x2_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B(n_613), .C(n_614), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g1068 ( .A1(n_612), .A2(n_887), .B1(n_1069), .B2(n_1070), .Y(n_1068) );
CKINVDCx20_ASAP7_75t_R g835 ( .A(n_615), .Y(n_835) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVxp67_ASAP7_75t_L g1026 ( .A(n_622), .Y(n_1026) );
BUFx4f_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g698 ( .A(n_627), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B1(n_662), .B2(n_663), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g661 ( .A(n_630), .Y(n_661) );
AND2x2_ASAP7_75t_SL g630 ( .A(n_631), .B(n_643), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_636), .Y(n_631) );
NAND2xp33_ASAP7_75t_SL g632 ( .A(n_633), .B(n_635), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_641), .Y(n_636) );
BUFx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g643 ( .A(n_644), .B(n_647), .C(n_654), .Y(n_643) );
OAI221xp5_ASAP7_75t_SL g780 ( .A1(n_649), .A2(n_781), .B1(n_782), .B2(n_783), .C(n_784), .Y(n_780) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B1(n_657), .B2(n_658), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g1150 ( .A1(n_656), .A2(n_658), .B1(n_1151), .B2(n_1152), .Y(n_1150) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_658), .A2(n_682), .B1(n_757), .B2(n_758), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_658), .A2(n_777), .B1(n_778), .B2(n_779), .Y(n_776) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_658), .A2(n_778), .B1(n_839), .B2(n_840), .Y(n_838) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g871 ( .A(n_659), .Y(n_871) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_SL g667 ( .A(n_668), .B(n_685), .Y(n_667) );
NOR3xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_674), .C(n_680), .Y(n_668) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g787 ( .A(n_672), .Y(n_787) );
INVx2_ASAP7_75t_L g831 ( .A(n_672), .Y(n_831) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx4_ASAP7_75t_L g727 ( .A(n_677), .Y(n_727) );
BUFx2_ASAP7_75t_L g867 ( .A(n_677), .Y(n_867) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx3_ASAP7_75t_SL g778 ( .A(n_683), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_693), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_687), .B(n_691), .Y(n_686) );
BUFx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g1024 ( .A(n_690), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_732), .B1(n_820), .B2(n_821), .Y(n_700) );
INVx2_ASAP7_75t_L g821 ( .A(n_701), .Y(n_821) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_703), .B(n_721), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_710), .C(n_715), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_708), .Y(n_704) );
INVx1_ASAP7_75t_L g743 ( .A(n_709), .Y(n_743) );
INVx2_ASAP7_75t_L g911 ( .A(n_712), .Y(n_911) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_718), .A2(n_749), .B1(n_750), .B2(n_752), .Y(n_748) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g1021 ( .A(n_719), .Y(n_1021) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_729), .Y(n_721) );
OAI21xp5_ASAP7_75t_SL g722 ( .A1(n_723), .A2(n_724), .B(n_725), .Y(n_722) );
INVx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g820 ( .A(n_732), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_762), .B1(n_818), .B2(n_819), .Y(n_732) );
INVx1_ASAP7_75t_L g818 ( .A(n_733), .Y(n_818) );
INVx1_ASAP7_75t_L g761 ( .A(n_734), .Y(n_761) );
AND4x1_ASAP7_75t_L g734 ( .A(n_735), .B(n_744), .C(n_753), .D(n_759), .Y(n_734) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_740), .B1(n_742), .B2(n_743), .Y(n_738) );
BUFx2_ASAP7_75t_R g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g916 ( .A(n_750), .Y(n_916) );
INVx3_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
BUFx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g819 ( .A(n_762), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_792), .B1(n_793), .B2(n_817), .Y(n_762) );
INVx1_ASAP7_75t_L g817 ( .A(n_763), .Y(n_817) );
INVx1_ASAP7_75t_SL g791 ( .A(n_764), .Y(n_791) );
AND2x2_ASAP7_75t_SL g764 ( .A(n_765), .B(n_775), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_770), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
BUFx2_ASAP7_75t_L g913 ( .A(n_769), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_774), .Y(n_770) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NOR3xp33_ASAP7_75t_SL g775 ( .A(n_776), .B(n_780), .C(n_785), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_778), .A2(n_869), .B1(n_870), .B2(n_871), .Y(n_868) );
OAI21xp5_ASAP7_75t_SL g797 ( .A1(n_781), .A2(n_798), .B(n_799), .Y(n_797) );
OAI221xp5_ASAP7_75t_L g1113 ( .A1(n_781), .A2(n_895), .B1(n_1114), .B2(n_1115), .C(n_1116), .Y(n_1113) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_787), .B1(n_788), .B2(n_789), .Y(n_785) );
INVx2_ASAP7_75t_SL g792 ( .A(n_793), .Y(n_792) );
XOR2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_816), .Y(n_794) );
NAND3x1_ASAP7_75t_L g795 ( .A(n_796), .B(n_809), .C(n_812), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_801), .Y(n_796) );
NAND3xp33_ASAP7_75t_L g801 ( .A(n_802), .B(n_804), .C(n_807), .Y(n_801) );
BUFx6f_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
AND2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
AND2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
INVx1_ASAP7_75t_L g1092 ( .A(n_823), .Y(n_1092) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_825), .B1(n_936), .B2(n_1090), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_852), .B1(n_853), .B2(n_935), .Y(n_825) );
INVx1_ASAP7_75t_L g935 ( .A(n_826), .Y(n_935) );
INVx2_ASAP7_75t_L g851 ( .A(n_827), .Y(n_851) );
AND2x2_ASAP7_75t_L g827 ( .A(n_828), .B(n_841), .Y(n_827) );
NOR3xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_833), .C(n_838), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_831), .A2(n_889), .B1(n_942), .B2(n_943), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g968 ( .A1(n_831), .A2(n_889), .B1(n_969), .B2(n_970), .Y(n_968) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_847), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_845), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_848), .B(n_849), .Y(n_847) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_856), .B1(n_906), .B2(n_934), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
XNOR2xp5_ASAP7_75t_L g856 ( .A(n_857), .B(n_882), .Y(n_856) );
XOR2x2_ASAP7_75t_L g857 ( .A(n_858), .B(n_881), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_872), .Y(n_858) );
NOR3xp33_ASAP7_75t_L g859 ( .A(n_860), .B(n_863), .C(n_868), .Y(n_859) );
OAI21xp33_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_865), .B(n_866), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g872 ( .A(n_873), .B(n_877), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_878), .B(n_879), .Y(n_877) );
XOR2x2_ASAP7_75t_L g882 ( .A(n_883), .B(n_905), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_884), .B(n_897), .Y(n_883) );
NOR3xp33_ASAP7_75t_L g884 ( .A(n_885), .B(n_890), .C(n_893), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_887), .B1(n_888), .B2(n_889), .Y(n_885) );
NOR2xp33_ASAP7_75t_L g897 ( .A(n_898), .B(n_902), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_899), .B(n_900), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
INVx1_ASAP7_75t_L g934 ( .A(n_906), .Y(n_934) );
INVx2_ASAP7_75t_L g933 ( .A(n_907), .Y(n_933) );
AND2x2_ASAP7_75t_SL g907 ( .A(n_908), .B(n_921), .Y(n_907) );
NOR2xp33_ASAP7_75t_L g908 ( .A(n_909), .B(n_914), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_910), .B(n_912), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_915), .B(n_919), .Y(n_914) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
NOR3xp33_ASAP7_75t_L g921 ( .A(n_922), .B(n_925), .C(n_929), .Y(n_921) );
INVx2_ASAP7_75t_L g1090 ( .A(n_936), .Y(n_1090) );
AOI22xp5_ASAP7_75t_L g936 ( .A1(n_937), .A2(n_961), .B1(n_1088), .B2(n_1089), .Y(n_936) );
INVxp67_ASAP7_75t_L g1088 ( .A(n_937), .Y(n_1088) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx1_ASAP7_75t_SL g959 ( .A(n_939), .Y(n_959) );
AND2x2_ASAP7_75t_SL g939 ( .A(n_940), .B(n_951), .Y(n_939) );
NOR3xp33_ASAP7_75t_L g940 ( .A(n_941), .B(n_944), .C(n_948), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_952), .B(n_955), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_953), .B(n_954), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_956), .B(n_958), .Y(n_955) );
INVx1_ASAP7_75t_L g1089 ( .A(n_961), .Y(n_1089) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_962), .A2(n_963), .B1(n_1008), .B2(n_1087), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g963 ( .A1(n_964), .A2(n_965), .B1(n_989), .B2(n_990), .Y(n_963) );
INVx2_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx2_ASAP7_75t_SL g988 ( .A(n_966), .Y(n_988) );
AND2x2_ASAP7_75t_L g966 ( .A(n_967), .B(n_980), .Y(n_966) );
NOR3xp33_ASAP7_75t_L g967 ( .A(n_968), .B(n_971), .C(n_977), .Y(n_967) );
OAI221xp5_ASAP7_75t_SL g971 ( .A1(n_972), .A2(n_973), .B1(n_974), .B2(n_975), .C(n_976), .Y(n_971) );
OAI221xp5_ASAP7_75t_L g1146 ( .A1(n_972), .A2(n_974), .B1(n_1147), .B2(n_1148), .C(n_1149), .Y(n_1146) );
NOR2xp33_ASAP7_75t_L g980 ( .A(n_981), .B(n_984), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_982), .B(n_983), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_985), .B(n_986), .Y(n_984) );
INVx2_ASAP7_75t_SL g989 ( .A(n_990), .Y(n_989) );
XNOR2x2_ASAP7_75t_L g990 ( .A(n_991), .B(n_992), .Y(n_990) );
NOR4xp75_ASAP7_75t_L g992 ( .A(n_993), .B(n_996), .C(n_999), .D(n_1003), .Y(n_992) );
NAND2xp5_ASAP7_75t_SL g993 ( .A(n_994), .B(n_995), .Y(n_993) );
NAND2xp5_ASAP7_75t_SL g996 ( .A(n_997), .B(n_998), .Y(n_996) );
OAI21xp5_ASAP7_75t_SL g1003 ( .A1(n_1004), .A2(n_1006), .B(n_1007), .Y(n_1003) );
OAI21xp5_ASAP7_75t_SL g1047 ( .A1(n_1004), .A2(n_1048), .B(n_1049), .Y(n_1047) );
INVx3_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx2_ASAP7_75t_SL g1087 ( .A(n_1008), .Y(n_1087) );
OA22x2_ASAP7_75t_L g1008 ( .A1(n_1009), .A2(n_1042), .B1(n_1085), .B2(n_1086), .Y(n_1008) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1009), .Y(n_1085) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1010), .Y(n_1041) );
AND2x2_ASAP7_75t_SL g1010 ( .A(n_1011), .B(n_1027), .Y(n_1010) );
NOR3xp33_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1017), .C(n_1022), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1014), .Y(n_1012) );
HB1xp67_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_1018), .A2(n_1019), .B1(n_1020), .B2(n_1021), .Y(n_1017) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_1023), .A2(n_1024), .B1(n_1025), .B2(n_1026), .Y(n_1022) );
NOR3xp33_ASAP7_75t_SL g1027 ( .A(n_1028), .B(n_1031), .C(n_1037), .Y(n_1027) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1042), .Y(n_1086) );
XOR2x2_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1064), .Y(n_1042) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1045), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1056), .Y(n_1045) );
NOR2xp67_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1050), .Y(n_1046) );
NAND3xp33_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1054), .C(n_1055), .Y(n_1050) );
INVx1_ASAP7_75t_SL g1052 ( .A(n_1053), .Y(n_1052) );
NOR2x1_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1060), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1059), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1062), .Y(n_1060) );
INVx2_ASAP7_75t_L g1084 ( .A(n_1066), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1077), .Y(n_1066) );
NOR3xp33_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1071), .C(n_1074), .Y(n_1067) );
NOR2xp33_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1081), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1080), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1083), .Y(n_1081) );
INVx1_ASAP7_75t_SL g1093 ( .A(n_1094), .Y(n_1093) );
NOR2x1_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1099), .Y(n_1094) );
OR2x2_ASAP7_75t_SL g1164 ( .A(n_1095), .B(n_1100), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1098), .Y(n_1095) );
CKINVDCx20_ASAP7_75t_R g1131 ( .A(n_1096), .Y(n_1131) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_1097), .B(n_1134), .Y(n_1138) );
CKINVDCx16_ASAP7_75t_R g1134 ( .A(n_1098), .Y(n_1134) );
CKINVDCx20_ASAP7_75t_R g1099 ( .A(n_1100), .Y(n_1099) );
NAND2xp5_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1102), .Y(n_1100) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1105), .Y(n_1103) );
OAI322xp33_ASAP7_75t_L g1106 ( .A1(n_1107), .A2(n_1130), .A3(n_1132), .B1(n_1135), .B2(n_1139), .C1(n_1140), .C2(n_1162), .Y(n_1106) );
INVx2_ASAP7_75t_L g1129 ( .A(n_1108), .Y(n_1129) );
AND2x2_ASAP7_75t_SL g1108 ( .A(n_1109), .B(n_1120), .Y(n_1108) );
NOR3xp33_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1113), .C(n_1117), .Y(n_1109) );
NOR2xp33_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1124), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1123), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1126), .Y(n_1124) );
HB1xp67_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
HB1xp67_ASAP7_75t_L g1132 ( .A(n_1133), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
CKINVDCx20_ASAP7_75t_R g1136 ( .A(n_1137), .Y(n_1136) );
INVx2_ASAP7_75t_L g1161 ( .A(n_1141), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1153), .Y(n_1141) );
NOR3xp33_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1146), .C(n_1150), .Y(n_1142) );
NOR2xp33_ASAP7_75t_L g1153 ( .A(n_1154), .B(n_1157), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1156), .Y(n_1154) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1159), .Y(n_1157) );
CKINVDCx20_ASAP7_75t_R g1162 ( .A(n_1163), .Y(n_1162) );
CKINVDCx20_ASAP7_75t_R g1163 ( .A(n_1164), .Y(n_1163) );
endmodule