module fake_jpeg_22680_n_290 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_29),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_47),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_20),
.B(n_0),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_54),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_27),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_66),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_18),
.B1(n_21),
.B2(n_31),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_67),
.B1(n_69),
.B2(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_74),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_27),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_21),
.B1(n_31),
.B2(n_33),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_21),
.B1(n_31),
.B2(n_33),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_33),
.B(n_35),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_24),
.B(n_25),
.C(n_40),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_30),
.B1(n_22),
.B2(n_26),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_28),
.B1(n_22),
.B2(n_26),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_39),
.B1(n_38),
.B2(n_34),
.Y(n_96)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_39),
.B1(n_28),
.B2(n_30),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_84),
.B1(n_87),
.B2(n_72),
.Y(n_105)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_78),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_23),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_37),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_45),
.Y(n_79)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_83),
.A2(n_53),
.B1(n_71),
.B2(n_68),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_20),
.B1(n_37),
.B2(n_36),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_36),
.C(n_32),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_1),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_42),
.A2(n_32),
.B1(n_35),
.B2(n_34),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_57),
.A2(n_39),
.B1(n_46),
.B2(n_35),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_94),
.A2(n_104),
.B1(n_119),
.B2(n_103),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_97),
.B1(n_114),
.B2(n_84),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_39),
.B1(n_46),
.B2(n_38),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_55),
.A2(n_41),
.B1(n_40),
.B2(n_46),
.Y(n_100)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_54),
.A3(n_59),
.B1(n_56),
.B2(n_61),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_66),
.A2(n_34),
.B1(n_25),
.B2(n_24),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_105),
.B1(n_51),
.B2(n_60),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_75),
.C(n_78),
.Y(n_126)
);

AO22x2_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_41),
.B1(n_40),
.B2(n_25),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_24),
.B1(n_23),
.B2(n_5),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_64),
.A2(n_86),
.B1(n_71),
.B2(n_68),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_6),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_69),
.A2(n_41),
.B1(n_4),
.B2(n_5),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_80),
.B(n_41),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_1),
.C(n_4),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_91),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_130),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_126),
.A2(n_138),
.B(n_94),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_133),
.B1(n_134),
.B2(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_64),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_129),
.B(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_135),
.Y(n_180)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_41),
.B(n_89),
.C(n_82),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_136),
.B(n_138),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_54),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_65),
.B(n_4),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_144),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_65),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_146),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_118),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_5),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_145),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_93),
.Y(n_146)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_148),
.A2(n_149),
.B1(n_92),
.B2(n_112),
.Y(n_174)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_150),
.B(n_100),
.Y(n_178)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_98),
.B(n_7),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_104),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_11),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_96),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_154),
.A2(n_93),
.B1(n_121),
.B2(n_112),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_156),
.A2(n_170),
.B(n_172),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_142),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_159),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_115),
.Y(n_160)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_160),
.B(n_150),
.C(n_13),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_154),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_164),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_99),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_176),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_100),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_173),
.B(n_181),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

AND2x4_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_100),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_178),
.C(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_130),
.B(n_8),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_179),
.B(n_12),
.Y(n_186)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_182),
.A2(n_133),
.B1(n_124),
.B2(n_153),
.Y(n_187)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_185),
.B(n_135),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_186),
.B(n_205),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_193),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_163),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_180),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_202),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_176),
.A2(n_132),
.B1(n_127),
.B2(n_125),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_207),
.B1(n_156),
.B2(n_175),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_149),
.C(n_140),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_206),
.C(n_181),
.Y(n_210)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_150),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_204),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_179),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_169),
.B1(n_162),
.B2(n_168),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_101),
.C(n_120),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_161),
.A2(n_127),
.B1(n_125),
.B2(n_92),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_201),
.Y(n_223)
);

A2O1A1O1Ixp25_ASAP7_75t_L g217 ( 
.A1(n_209),
.A2(n_160),
.B(n_178),
.C(n_175),
.D(n_182),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_206),
.C(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_185),
.B1(n_171),
.B2(n_110),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_167),
.B1(n_161),
.B2(n_166),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_224),
.B1(n_227),
.B2(n_195),
.Y(n_236)
);

NOR3xp33_ASAP7_75t_SL g231 ( 
.A(n_217),
.B(n_221),
.C(n_200),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_220),
.A2(n_223),
.B1(n_110),
.B2(n_107),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_201),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_226),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_191),
.A2(n_166),
.B1(n_175),
.B2(n_172),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_157),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_190),
.A2(n_172),
.B1(n_173),
.B2(n_155),
.Y(n_227)
);

OAI322xp33_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_203),
.A3(n_198),
.B1(n_188),
.B2(n_200),
.C1(n_189),
.C2(n_197),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_SL g252 ( 
.A(n_229),
.B(n_227),
.C(n_228),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_196),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_228),
.Y(n_249)
);

AOI31xp67_ASAP7_75t_L g247 ( 
.A1(n_231),
.A2(n_243),
.A3(n_217),
.B(n_214),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_198),
.A3(n_190),
.B1(n_187),
.B2(n_203),
.C1(n_202),
.C2(n_208),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g253 ( 
.A(n_233),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_242),
.C(n_244),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_236),
.B(n_238),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_193),
.B1(n_194),
.B2(n_155),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_186),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_219),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_107),
.C(n_120),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_108),
.C(n_13),
.Y(n_244)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_231),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_215),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_251),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_234),
.C(n_241),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_254),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_216),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_212),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_255),
.B(n_230),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_212),
.C(n_225),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_257),
.B(n_258),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_108),
.C(n_14),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_260),
.B(n_262),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_240),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_268),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_236),
.B(n_252),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_256),
.B(n_232),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_245),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_272),
.C(n_273),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_271),
.B(n_274),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_245),
.B1(n_243),
.B2(n_246),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_253),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_12),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_260),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_278),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_267),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_279),
.A2(n_275),
.B(n_264),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_259),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_280),
.B(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_14),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_14),
.B(n_15),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_281),
.C(n_15),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_285),
.A2(n_287),
.B(n_286),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_16),
.B(n_17),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_17),
.Y(n_290)
);


endmodule