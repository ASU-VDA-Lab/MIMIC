module real_aes_4520_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_919;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_908;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_918;
wire n_478;
wire n_356;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_892;
wire n_372;
wire n_528;
wire n_202;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_906;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_931;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_298;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_926;
wire n_922;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g546 ( .A(n_0), .B(n_219), .Y(n_546) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_1), .Y(n_559) );
O2A1O1Ixp33_ASAP7_75t_SL g595 ( .A1(n_2), .A2(n_134), .B(n_596), .C(n_597), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g551 ( .A1(n_3), .A2(n_79), .B1(n_123), .B2(n_202), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_4), .A2(n_29), .B1(n_177), .B2(n_180), .Y(n_176) );
INVx1_ASAP7_75t_L g530 ( .A(n_5), .Y(n_530) );
INVx1_ASAP7_75t_L g895 ( .A(n_5), .Y(n_895) );
INVxp67_ASAP7_75t_L g918 ( .A(n_5), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_6), .A2(n_86), .B1(n_260), .B2(n_261), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_7), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_8), .A2(n_67), .B1(n_179), .B2(n_202), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g151 ( .A1(n_9), .A2(n_30), .B1(n_132), .B2(n_152), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g612 ( .A(n_10), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_11), .A2(n_100), .B1(n_934), .B2(n_942), .Y(n_99) );
INVx2_ASAP7_75t_L g233 ( .A(n_12), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_13), .A2(n_60), .B1(n_123), .B2(n_153), .Y(n_587) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_14), .A2(n_66), .B(n_114), .Y(n_113) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_14), .A2(n_66), .B(n_114), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_15), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_SL g231 ( .A(n_16), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_17), .B(n_140), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_18), .Y(n_573) );
BUFx3_ASAP7_75t_L g924 ( .A(n_19), .Y(n_924) );
O2A1O1Ixp33_ASAP7_75t_L g600 ( .A1(n_20), .A2(n_155), .B(n_291), .C(n_601), .Y(n_600) );
OAI22xp33_ASAP7_75t_SL g549 ( .A1(n_21), .A2(n_44), .B1(n_123), .B2(n_130), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_22), .A2(n_28), .B1(n_130), .B2(n_162), .Y(n_639) );
CKINVDCx5p33_ASAP7_75t_R g908 ( .A(n_23), .Y(n_908) );
O2A1O1Ixp5_ASAP7_75t_L g281 ( .A1(n_24), .A2(n_157), .B(n_282), .C(n_285), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_25), .B(n_122), .Y(n_121) );
O2A1O1Ixp5_ASAP7_75t_L g675 ( .A1(n_26), .A2(n_134), .B(n_225), .C(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g535 ( .A(n_27), .Y(n_535) );
AND2x2_ASAP7_75t_L g939 ( .A(n_31), .B(n_940), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_32), .B(n_187), .Y(n_643) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_33), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_34), .A2(n_38), .B1(n_183), .B2(n_184), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_35), .A2(n_65), .B1(n_184), .B2(n_201), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g117 ( .A(n_36), .B(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g210 ( .A(n_37), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_39), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_40), .B(n_167), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_41), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_42), .A2(n_155), .B(n_228), .C(n_229), .Y(n_227) );
INVx1_ASAP7_75t_L g251 ( .A(n_43), .Y(n_251) );
INVx2_ASAP7_75t_L g292 ( .A(n_45), .Y(n_292) );
INVx1_ASAP7_75t_L g114 ( .A(n_46), .Y(n_114) );
AND2x4_ASAP7_75t_L g137 ( .A(n_47), .B(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g216 ( .A(n_47), .B(n_138), .Y(n_216) );
INVx2_ASAP7_75t_L g203 ( .A(n_48), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_49), .B(n_187), .Y(n_607) );
INVxp67_ASAP7_75t_SL g630 ( .A(n_49), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_49), .A2(n_64), .B1(n_187), .B2(n_651), .Y(n_650) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_50), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g914 ( .A(n_51), .Y(n_914) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_52), .Y(n_557) );
O2A1O1Ixp33_ASAP7_75t_L g574 ( .A1(n_53), .A2(n_134), .B(n_575), .C(n_576), .Y(n_574) );
INVx2_ASAP7_75t_L g617 ( .A(n_54), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g683 ( .A(n_55), .Y(n_683) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_56), .Y(n_556) );
INVx1_ASAP7_75t_SL g286 ( .A(n_57), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_58), .A2(n_929), .B1(n_930), .B2(n_931), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_58), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_59), .B(n_140), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_61), .A2(n_76), .B1(n_178), .B2(n_641), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_62), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_63), .Y(n_560) );
NAND2xp33_ASAP7_75t_R g590 ( .A(n_64), .B(n_113), .Y(n_590) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_68), .A2(n_155), .B(n_177), .C(n_206), .Y(n_205) );
OR2x6_ASAP7_75t_L g532 ( .A(n_69), .B(n_533), .Y(n_532) );
NAND3xp33_ASAP7_75t_L g938 ( .A(n_69), .B(n_918), .C(n_939), .Y(n_938) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_70), .Y(n_237) );
INVx1_ASAP7_75t_L g247 ( .A(n_71), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_72), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_73), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_74), .B(n_132), .Y(n_131) );
NOR2xp67_ASAP7_75t_L g224 ( .A(n_75), .B(n_225), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_77), .A2(n_134), .B(n_198), .C(n_200), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_77), .A2(n_134), .B(n_198), .C(n_200), .Y(n_330) );
INVx1_ASAP7_75t_L g534 ( .A(n_78), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_80), .A2(n_90), .B1(n_160), .B2(n_164), .Y(n_159) );
INVx1_ASAP7_75t_L g940 ( .A(n_81), .Y(n_940) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_82), .Y(n_120) );
BUFx5_ASAP7_75t_L g123 ( .A(n_82), .Y(n_123) );
INVx1_ASAP7_75t_L g163 ( .A(n_82), .Y(n_163) );
INVx2_ASAP7_75t_L g605 ( .A(n_83), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_84), .B(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g579 ( .A(n_85), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_87), .Y(n_602) );
INVx2_ASAP7_75t_SL g138 ( .A(n_88), .Y(n_138) );
INVx1_ASAP7_75t_L g681 ( .A(n_89), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_91), .B(n_113), .Y(n_248) );
INVx1_ASAP7_75t_SL g191 ( .A(n_92), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_93), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g685 ( .A(n_94), .Y(n_685) );
AND2x2_ASAP7_75t_L g168 ( .A(n_95), .B(n_169), .Y(n_168) );
OAI21xp33_ASAP7_75t_SL g571 ( .A1(n_96), .A2(n_123), .B(n_572), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g102 ( .A1(n_97), .A2(n_103), .B1(n_896), .B2(n_906), .C(n_907), .Y(n_102) );
INVx1_ASAP7_75t_L g906 ( .A(n_97), .Y(n_906) );
INVx1_ASAP7_75t_SL g290 ( .A(n_98), .Y(n_290) );
AO21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_919), .B(n_925), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_102), .B(n_912), .Y(n_101) );
OAI22xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_529), .B1(n_536), .B2(n_892), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g901 ( .A(n_104), .B(n_902), .Y(n_901) );
NAND2x1p5_ASAP7_75t_L g104 ( .A(n_105), .B(n_410), .Y(n_104) );
NOR2x1_ASAP7_75t_L g105 ( .A(n_106), .B(n_344), .Y(n_105) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_306), .Y(n_106) );
OAI21xp5_ASAP7_75t_SL g107 ( .A1(n_108), .A2(n_143), .B(n_267), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_108), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g321 ( .A(n_110), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g405 ( .A(n_110), .B(n_235), .Y(n_405) );
AND2x2_ASAP7_75t_L g430 ( .A(n_110), .B(n_402), .Y(n_430) );
OAI21x1_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_115), .B(n_139), .Y(n_110) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_111), .A2(n_257), .B(n_266), .Y(n_256) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_112), .B(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
BUFx3_ASAP7_75t_L g169 ( .A(n_113), .Y(n_169) );
INVx2_ASAP7_75t_L g190 ( .A(n_113), .Y(n_190) );
INVx1_ASAP7_75t_L g569 ( .A(n_113), .Y(n_569) );
INVx1_ASAP7_75t_L g686 ( .A(n_113), .Y(n_686) );
OAI21x1_ASAP7_75t_L g275 ( .A1(n_115), .A2(n_139), .B(n_253), .Y(n_275) );
OAI21x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_127), .B(n_135), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_121), .B(n_124), .Y(n_116) );
INVx1_ASAP7_75t_L g180 ( .A(n_118), .Y(n_180) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g225 ( .A(n_119), .Y(n_225) );
INVx2_ASAP7_75t_L g261 ( .A(n_119), .Y(n_261) );
INVx1_ASAP7_75t_L g575 ( .A(n_119), .Y(n_575) );
INVx1_ASAP7_75t_L g679 ( .A(n_119), .Y(n_679) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx6_ASAP7_75t_L g130 ( .A(n_120), .Y(n_130) );
INVx2_ASAP7_75t_L g153 ( .A(n_120), .Y(n_153) );
INVx2_ASAP7_75t_L g202 ( .A(n_120), .Y(n_202) );
INVx1_ASAP7_75t_L g183 ( .A(n_122), .Y(n_183) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g132 ( .A(n_123), .Y(n_132) );
INVx2_ASAP7_75t_L g164 ( .A(n_123), .Y(n_164) );
INVx1_ASAP7_75t_L g199 ( .A(n_123), .Y(n_199) );
NAND2xp33_ASAP7_75t_L g222 ( .A(n_123), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g260 ( .A(n_123), .Y(n_260) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_123), .A2(n_130), .B1(n_556), .B2(n_557), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_123), .A2(n_153), .B1(n_559), .B2(n_560), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_123), .B(n_573), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_123), .A2(n_130), .B1(n_612), .B2(n_613), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_123), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_123), .B(n_683), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_124), .A2(n_571), .B(n_574), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_124), .A2(n_215), .B1(n_610), .B2(n_614), .C(n_618), .Y(n_609) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
O2A1O1Ixp5_ASAP7_75t_SL g236 ( .A1(n_125), .A2(n_237), .B(n_238), .C(n_241), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_125), .A2(n_134), .B1(n_587), .B2(n_588), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g628 ( .A1(n_125), .A2(n_134), .B1(n_611), .B2(n_615), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_125), .A2(n_679), .B1(n_680), .B2(n_682), .Y(n_678) );
INVx4_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_126), .Y(n_134) );
INVx3_ASAP7_75t_L g155 ( .A(n_126), .Y(n_155) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_126), .Y(n_158) );
INVxp67_ASAP7_75t_L g263 ( .A(n_126), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_126), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g642 ( .A(n_126), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_126), .B(n_681), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_131), .B(n_133), .Y(n_127) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g230 ( .A(n_130), .Y(n_230) );
INVx1_ASAP7_75t_L g240 ( .A(n_130), .Y(n_240) );
INVx2_ASAP7_75t_L g284 ( .A(n_130), .Y(n_284) );
INVx2_ASAP7_75t_SL g641 ( .A(n_130), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_133), .A2(n_221), .B(n_224), .Y(n_220) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_134), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_134), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_SL g265 ( .A(n_134), .Y(n_265) );
OAI221xp5_ASAP7_75t_L g554 ( .A1(n_134), .A2(n_137), .B1(n_155), .B2(n_555), .C(n_558), .Y(n_554) );
INVx1_ASAP7_75t_L g618 ( .A(n_134), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_135), .B(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_136), .A2(n_248), .B(n_253), .Y(n_252) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g165 ( .A(n_137), .B(n_166), .Y(n_165) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_137), .Y(n_194) );
INVx1_ASAP7_75t_L g294 ( .A(n_137), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_137), .B(n_188), .Y(n_552) );
NOR2xp67_ASAP7_75t_L g589 ( .A(n_140), .B(n_294), .Y(n_589) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_141), .B(n_233), .Y(n_232) );
BUFx3_ASAP7_75t_L g254 ( .A(n_141), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_141), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx3_ASAP7_75t_L g167 ( .A(n_142), .Y(n_167) );
INVx4_ASAP7_75t_L g188 ( .A(n_142), .Y(n_188) );
NAND3xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_211), .C(n_255), .Y(n_143) );
AOI222xp33_ASAP7_75t_L g475 ( .A1(n_144), .A2(n_353), .B1(n_476), .B2(n_478), .C1(n_480), .C2(n_483), .Y(n_475) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OR2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_170), .Y(n_145) );
OR2x2_ASAP7_75t_L g432 ( .A(n_146), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g440 ( .A(n_146), .B(n_370), .Y(n_440) );
BUFx2_ASAP7_75t_SL g146 ( .A(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_147), .B(n_313), .Y(n_312) );
AND2x4_ASAP7_75t_L g327 ( .A(n_147), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g347 ( .A(n_147), .B(n_192), .Y(n_347) );
INVx1_ASAP7_75t_L g451 ( .A(n_147), .Y(n_451) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NAND2x1_ASAP7_75t_L g304 ( .A(n_148), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g334 ( .A(n_149), .Y(n_334) );
AO31x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_156), .A3(n_165), .B(n_168), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_154), .Y(n_150) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVxp67_ASAP7_75t_SL g228 ( .A(n_153), .Y(n_228) );
INVx1_ASAP7_75t_L g291 ( .A(n_153), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_153), .A2(n_162), .B1(n_616), .B2(n_617), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_154), .A2(n_182), .B(n_185), .Y(n_181) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_155), .A2(n_551), .B(n_552), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_159), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_157), .B(n_176), .Y(n_175) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
OA22x2_ASAP7_75t_L g638 ( .A1(n_158), .A2(n_639), .B1(n_640), .B2(n_642), .Y(n_638) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g184 ( .A(n_162), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_162), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_162), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g179 ( .A(n_163), .Y(n_179) );
INVx2_ASAP7_75t_L g245 ( .A(n_164), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_166), .B(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_166), .A2(n_696), .B(n_697), .Y(n_695) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_167), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g627 ( .A(n_169), .Y(n_627) );
OAI221xp5_ASAP7_75t_L g413 ( .A1(n_170), .A2(n_414), .B1(n_415), .B2(n_417), .C(n_421), .Y(n_413) );
NOR2x1_ASAP7_75t_L g428 ( .A(n_170), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g477 ( .A(n_170), .B(n_312), .Y(n_477) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NAND2x1p5_ASAP7_75t_L g442 ( .A(n_171), .B(n_303), .Y(n_442) );
AND2x4_ASAP7_75t_L g171 ( .A(n_172), .B(n_192), .Y(n_171) );
OR2x2_ASAP7_75t_L g326 ( .A(n_172), .B(n_314), .Y(n_326) );
AND2x2_ASAP7_75t_L g408 ( .A(n_172), .B(n_256), .Y(n_408) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g362 ( .A(n_173), .Y(n_362) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g305 ( .A(n_174), .Y(n_305) );
AOI21x1_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_181), .B(n_189), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_177), .B(n_286), .Y(n_285) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g596 ( .A(n_178), .Y(n_596) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AOI21x1_ASAP7_75t_L g314 ( .A1(n_186), .A2(n_315), .B(n_316), .Y(n_314) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g219 ( .A(n_188), .Y(n_219) );
NOR2xp33_ASAP7_75t_SL g604 ( .A(n_188), .B(n_605), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
INVx1_ASAP7_75t_L g296 ( .A(n_190), .Y(n_296) );
INVx1_ASAP7_75t_L g651 ( .A(n_190), .Y(n_651) );
NOR2x1_ASAP7_75t_L g317 ( .A(n_192), .B(n_305), .Y(n_317) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_195), .B(n_208), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_194), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_194), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_204), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_203), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_201), .B(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g289 ( .A(n_201), .Y(n_289) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g242 ( .A(n_202), .Y(n_242) );
INVxp67_ASAP7_75t_SL g204 ( .A(n_205), .Y(n_204) );
NOR4xp25_ASAP7_75t_L g329 ( .A(n_205), .B(n_215), .C(n_296), .D(n_330), .Y(n_329) );
INVxp67_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g328 ( .A(n_209), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_211), .B(n_308), .Y(n_307) );
OAI32xp33_ASAP7_75t_L g388 ( .A1(n_211), .A2(n_389), .A3(n_390), .B1(n_392), .B2(n_395), .Y(n_388) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g270 ( .A(n_212), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g375 ( .A(n_212), .B(n_376), .Y(n_375) );
NOR2xp67_ASAP7_75t_L g437 ( .A(n_212), .B(n_389), .Y(n_437) );
AND2x2_ASAP7_75t_L g460 ( .A(n_212), .B(n_393), .Y(n_460) );
AND2x2_ASAP7_75t_L g489 ( .A(n_212), .B(n_420), .Y(n_489) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_234), .Y(n_212) );
OR2x2_ASAP7_75t_L g297 ( .A(n_213), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g319 ( .A(n_213), .Y(n_319) );
AND2x2_ASAP7_75t_L g353 ( .A(n_213), .B(n_298), .Y(n_353) );
INVx2_ASAP7_75t_L g384 ( .A(n_213), .Y(n_384) );
OR2x2_ASAP7_75t_L g394 ( .A(n_213), .B(n_234), .Y(n_394) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_213), .Y(n_468) );
AO31x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_220), .A3(n_226), .B(n_232), .Y(n_213) );
NOR2x1_ASAP7_75t_SL g214 ( .A(n_215), .B(n_217), .Y(n_214) );
NOR2xp33_ASAP7_75t_SL g603 ( .A(n_215), .B(n_219), .Y(n_603) );
NOR3xp33_ASAP7_75t_L g674 ( .A(n_215), .B(n_675), .C(n_678), .Y(n_674) );
INVx4_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g568 ( .A(n_216), .B(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_216), .B(n_627), .Y(n_637) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_217), .A2(n_554), .B(n_561), .Y(n_553) );
OA21x2_ASAP7_75t_L g657 ( .A1(n_217), .A2(n_554), .B(n_561), .Y(n_657) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g629 ( .A(n_218), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_230), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g349 ( .A(n_234), .B(n_279), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_234), .B(n_273), .Y(n_515) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g368 ( .A(n_235), .B(n_274), .Y(n_368) );
OAI21x1_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_243), .B(n_252), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g298 ( .A1(n_236), .A2(n_243), .B(n_252), .Y(n_298) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_239), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND3x1_ASAP7_75t_L g243 ( .A(n_244), .B(n_248), .C(n_249), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_254), .B(n_609), .Y(n_608) );
AO21x2_ASAP7_75t_L g673 ( .A1(n_254), .A2(n_674), .B(n_684), .Y(n_673) );
OAI32xp33_ASAP7_75t_L g351 ( .A1(n_255), .A2(n_352), .A3(n_353), .B1(n_354), .B2(n_355), .Y(n_351) );
INVx1_ASAP7_75t_L g429 ( .A(n_255), .Y(n_429) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_256), .Y(n_303) );
INVx1_ASAP7_75t_L g336 ( .A(n_256), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_256), .B(n_334), .Y(n_359) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_258), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_262), .B1(n_264), .B2(n_265), .Y(n_258) );
OAI21xp5_ASAP7_75t_SL g287 ( .A1(n_262), .A2(n_288), .B(n_293), .Y(n_287) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g316 ( .A(n_266), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_299), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_276), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_269), .A2(n_354), .B1(n_378), .B2(n_381), .Y(n_377) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2x1p5_ASAP7_75t_L g414 ( .A(n_272), .B(n_349), .Y(n_414) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx2_ASAP7_75t_SL g343 ( .A(n_273), .Y(n_343) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_273), .Y(n_350) );
AND2x2_ASAP7_75t_L g403 ( .A(n_273), .B(n_384), .Y(n_403) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g278 ( .A(n_274), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g420 ( .A(n_274), .B(n_402), .Y(n_420) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_297), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
BUFx2_ASAP7_75t_L g308 ( .A(n_278), .Y(n_308) );
NAND2x1_ASAP7_75t_SL g479 ( .A(n_278), .B(n_468), .Y(n_479) );
INVx2_ASAP7_75t_SL g340 ( .A(n_279), .Y(n_340) );
BUFx2_ASAP7_75t_L g386 ( .A(n_279), .Y(n_386) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx3_ASAP7_75t_L g322 ( .A(n_280), .Y(n_322) );
INVx1_ASAP7_75t_L g357 ( .A(n_280), .Y(n_357) );
OA21x2_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_287), .B(n_295), .Y(n_280) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_290), .B1(n_291), .B2(n_292), .Y(n_288) );
OR2x2_ASAP7_75t_L g452 ( .A(n_297), .B(n_453), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_297), .B(n_352), .C(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g505 ( .A(n_297), .B(n_365), .Y(n_505) );
INVx1_ASAP7_75t_L g517 ( .A(n_297), .Y(n_517) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_298), .Y(n_418) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_300), .A2(n_446), .B1(n_450), .B2(n_452), .Y(n_445) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g500 ( .A(n_301), .B(n_463), .Y(n_500) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g462 ( .A(n_302), .B(n_463), .Y(n_462) );
NOR2x1p5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx2_ASAP7_75t_L g398 ( .A(n_303), .Y(n_398) );
INVx2_ASAP7_75t_L g511 ( .A(n_303), .Y(n_511) );
OR2x2_ASAP7_75t_L g484 ( .A(n_304), .B(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g370 ( .A(n_305), .B(n_314), .Y(n_370) );
INVx1_ASAP7_75t_L g426 ( .A(n_305), .Y(n_426) );
OAI222xp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_309), .B1(n_318), .B2(n_323), .C1(n_331), .C2(n_337), .Y(n_306) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_317), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g494 ( .A(n_313), .B(n_362), .Y(n_494) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_317), .B(n_333), .Y(n_380) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx2_ASAP7_75t_SL g342 ( .A(n_319), .Y(n_342) );
AND2x4_ASAP7_75t_L g423 ( .A(n_319), .B(n_405), .Y(n_423) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g389 ( .A(n_321), .Y(n_389) );
INVx2_ASAP7_75t_L g402 ( .A(n_322), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_322), .B(n_449), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_323), .A2(n_502), .B(n_504), .C(n_505), .Y(n_501) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
AND2x4_ASAP7_75t_L g346 ( .A(n_325), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g450 ( .A(n_326), .B(n_451), .Y(n_450) );
AND2x4_ASAP7_75t_L g369 ( .A(n_327), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_327), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_SL g409 ( .A(n_327), .Y(n_409) );
AND2x2_ASAP7_75t_L g496 ( .A(n_327), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g503 ( .A(n_327), .Y(n_503) );
NOR2x1_ASAP7_75t_L g335 ( .A(n_328), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_328), .B(n_361), .Y(n_360) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_328), .Y(n_391) );
INVx1_ASAP7_75t_L g396 ( .A(n_328), .Y(n_396) );
INVx1_ASAP7_75t_L g472 ( .A(n_328), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_331), .B(n_373), .Y(n_372) );
OAI22xp33_ASAP7_75t_L g431 ( .A1(n_331), .A2(n_363), .B1(n_432), .B2(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g455 ( .A(n_332), .B(n_426), .Y(n_455) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_333), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g492 ( .A(n_333), .Y(n_492) );
BUFx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g485 ( .A(n_335), .Y(n_485) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
NOR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g365 ( .A(n_340), .Y(n_365) );
AND2x2_ASAP7_75t_L g367 ( .A(n_340), .B(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_340), .B(n_470), .Y(n_469) );
OR2x6_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g376 ( .A(n_343), .Y(n_376) );
NAND3xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_371), .C(n_387), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_348), .B1(n_351), .B2(n_363), .C(n_366), .Y(n_345) );
INVx1_ASAP7_75t_L g354 ( .A(n_347), .Y(n_354) );
AND2x2_ASAP7_75t_L g416 ( .A(n_347), .B(n_370), .Y(n_416) );
AND2x2_ASAP7_75t_L g424 ( .A(n_347), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g510 ( .A(n_347), .B(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g364 ( .A(n_353), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
BUFx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_R g393 ( .A(n_357), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g519 ( .A(n_359), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_360), .Y(n_520) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g374 ( .A(n_362), .Y(n_374) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_362), .Y(n_497) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
AND2x2_ASAP7_75t_L g467 ( .A(n_367), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g435 ( .A(n_368), .Y(n_435) );
AND2x2_ASAP7_75t_L g499 ( .A(n_368), .B(n_384), .Y(n_499) );
AND2x2_ASAP7_75t_L g385 ( .A(n_370), .B(n_386), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_375), .B(n_377), .Y(n_371) );
OAI221xp5_ASAP7_75t_L g507 ( .A1(n_378), .A2(n_508), .B1(n_509), .B2(n_512), .C(n_516), .Y(n_507) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g528 ( .A(n_380), .Y(n_528) );
NAND2x1_ASAP7_75t_L g381 ( .A(n_382), .B(n_385), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g434 ( .A(n_384), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g449 ( .A(n_384), .Y(n_449) );
INVx1_ASAP7_75t_L g481 ( .A(n_386), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_397), .B(n_399), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI222xp33_ASAP7_75t_L g487 ( .A1(n_392), .A2(n_488), .B1(n_490), .B2(n_495), .C1(n_498), .C2(n_500), .Y(n_487) );
OR2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
AND2x2_ASAP7_75t_L g422 ( .A(n_393), .B(n_405), .Y(n_422) );
AND2x2_ASAP7_75t_L g513 ( .A(n_393), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g482 ( .A(n_394), .Y(n_482) );
INVx1_ASAP7_75t_L g526 ( .A(n_394), .Y(n_526) );
INVx1_ASAP7_75t_L g463 ( .A(n_396), .Y(n_463) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g474 ( .A(n_398), .Y(n_474) );
AOI21xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_404), .B(n_406), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g433 ( .A(n_408), .Y(n_433) );
INVx1_ASAP7_75t_L g504 ( .A(n_408), .Y(n_504) );
NOR2x1p5_ASAP7_75t_L g410 ( .A(n_411), .B(n_464), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_436), .C(n_454), .Y(n_411) );
NOR3xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_427), .C(n_431), .Y(n_412) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_414), .A2(n_444), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AO22x1_ASAP7_75t_L g427 ( .A1(n_416), .A2(n_422), .B1(n_428), .B2(n_430), .Y(n_427) );
OR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g444 ( .A(n_420), .Y(n_444) );
INVx1_ASAP7_75t_L g453 ( .A(n_420), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B(n_424), .Y(n_421) );
INVx2_ASAP7_75t_L g470 ( .A(n_423), .Y(n_470) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g461 ( .A(n_430), .Y(n_461) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_435), .B(n_448), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_441), .B2(n_443), .C(n_445), .Y(n_436) );
INVxp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_448), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B1(n_458), .B2(n_462), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND4xp75_ASAP7_75t_L g464 ( .A(n_465), .B(n_486), .C(n_506), .D(n_521), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_475), .Y(n_465) );
OAI21xp33_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_469), .B(n_471), .Y(n_466) );
INVx1_ASAP7_75t_L g523 ( .A(n_468), .Y(n_523) );
NOR2xp33_ASAP7_75t_SL g471 ( .A(n_472), .B(n_473), .Y(n_471) );
AND2x4_ASAP7_75t_L g527 ( .A(n_473), .B(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g508 ( .A(n_479), .Y(n_508) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NOR2x1_ASAP7_75t_L g486 ( .A(n_487), .B(n_501), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_524), .B(n_527), .Y(n_521) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g905 ( .A(n_529), .Y(n_905) );
OR2x6_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_531), .B(n_918), .Y(n_917) );
INVx8_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g894 ( .A(n_532), .B(n_895), .Y(n_894) );
OR2x6_ASAP7_75t_L g911 ( .A(n_532), .B(n_895), .Y(n_911) );
HB1xp67_ASAP7_75t_L g941 ( .A(n_533), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g900 ( .A(n_536), .Y(n_900) );
INVx2_ASAP7_75t_L g933 ( .A(n_536), .Y(n_933) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_806), .Y(n_536) );
NAND4xp25_ASAP7_75t_L g537 ( .A(n_538), .B(n_703), .C(n_758), .D(n_787), .Y(n_537) );
NOR2xp67_ASAP7_75t_L g538 ( .A(n_539), .B(n_619), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_580), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI221xp5_ASAP7_75t_SL g704 ( .A1(n_541), .A2(n_705), .B1(n_711), .B2(n_713), .C(n_716), .Y(n_704) );
OR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_562), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g788 ( .A(n_543), .B(n_789), .Y(n_788) );
OAI21xp33_ASAP7_75t_L g888 ( .A1(n_543), .A2(n_889), .B(n_891), .Y(n_888) );
AND2x4_ASAP7_75t_L g543 ( .A(n_544), .B(n_553), .Y(n_543) );
AND2x2_ASAP7_75t_L g692 ( .A(n_544), .B(n_566), .Y(n_692) );
INVx1_ASAP7_75t_L g783 ( .A(n_544), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_544), .B(n_671), .Y(n_825) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_545), .Y(n_654) );
INVx2_ASAP7_75t_L g665 ( .A(n_545), .Y(n_665) );
NAND2xp33_ASAP7_75t_R g721 ( .A(n_545), .B(n_566), .Y(n_721) );
INVx1_ASAP7_75t_L g744 ( .A(n_545), .Y(n_744) );
AND2x2_ASAP7_75t_L g751 ( .A(n_545), .B(n_553), .Y(n_751) );
AND2x2_ASAP7_75t_L g763 ( .A(n_545), .B(n_566), .Y(n_763) );
AND2x4_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
AND2x2_ASAP7_75t_L g634 ( .A(n_553), .B(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g694 ( .A(n_553), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g731 ( .A(n_553), .B(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g785 ( .A(n_562), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2x1p5_ASAP7_75t_L g663 ( .A(n_563), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_563), .B(n_712), .Y(n_795) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g645 ( .A(n_565), .Y(n_645) );
AND2x2_ASAP7_75t_L g866 ( .A(n_565), .B(n_751), .Y(n_866) );
AND2x2_ASAP7_75t_L g889 ( .A(n_565), .B(n_890), .Y(n_889) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g658 ( .A(n_566), .Y(n_658) );
INVx2_ASAP7_75t_L g671 ( .A(n_566), .Y(n_671) );
OR2x2_ASAP7_75t_L g756 ( .A(n_566), .B(n_665), .Y(n_756) );
AND2x2_ASAP7_75t_L g803 ( .A(n_566), .B(n_656), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_566), .B(n_657), .Y(n_821) );
BUFx2_ASAP7_75t_L g853 ( .A(n_566), .Y(n_853) );
INVx3_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AOI21x1_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_570), .B(n_578), .Y(n_567) );
AOI221xp5_ASAP7_75t_L g787 ( .A1(n_580), .A2(n_788), .B1(n_790), .B2(n_793), .C(n_796), .Y(n_787) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_591), .Y(n_581) );
OR2x2_ASAP7_75t_L g622 ( .A(n_582), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_582), .B(n_624), .Y(n_815) );
OR2x2_ASAP7_75t_L g848 ( .A(n_582), .B(n_723), .Y(n_848) );
INVx2_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g662 ( .A(n_584), .B(n_625), .Y(n_662) );
INVx2_ASAP7_75t_L g710 ( .A(n_584), .Y(n_710) );
AND2x2_ASAP7_75t_L g754 ( .A(n_584), .B(n_715), .Y(n_754) );
INVx1_ASAP7_75t_L g768 ( .A(n_584), .Y(n_768) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_590), .Y(n_584) );
AND2x2_ASAP7_75t_L g649 ( .A(n_585), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
INVxp67_ASAP7_75t_SL g811 ( .A(n_591), .Y(n_811) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g805 ( .A(n_592), .B(n_709), .Y(n_805) );
AND2x2_ASAP7_75t_L g878 ( .A(n_592), .B(n_767), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_592), .B(n_882), .Y(n_881) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_606), .Y(n_592) );
AND2x4_ASAP7_75t_L g624 ( .A(n_593), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g661 ( .A(n_593), .Y(n_661) );
INVx1_ASAP7_75t_L g708 ( .A(n_593), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_593), .B(n_673), .Y(n_719) );
INVx2_ASAP7_75t_L g725 ( .A(n_593), .Y(n_725) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_593), .Y(n_771) );
OR2x2_ASAP7_75t_L g792 ( .A(n_593), .B(n_606), .Y(n_792) );
HB1xp67_ASAP7_75t_L g886 ( .A(n_593), .Y(n_886) );
AO31x2_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_599), .A3(n_603), .B(n_604), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g688 ( .A(n_606), .B(n_661), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_606), .B(n_672), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_606), .B(n_841), .Y(n_840) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
AND2x2_ASAP7_75t_L g648 ( .A(n_608), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_667), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_631), .B(n_646), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
OAI21xp33_ASAP7_75t_L g772 ( .A1(n_624), .A2(n_773), .B(n_775), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_624), .B(n_767), .Y(n_775) );
AND2x2_ASAP7_75t_L g867 ( .A(n_624), .B(n_709), .Y(n_867) );
AND2x2_ASAP7_75t_L g891 ( .A(n_624), .B(n_754), .Y(n_891) );
INVx1_ASAP7_75t_L g699 ( .A(n_625), .Y(n_699) );
OAI21x1_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_628), .B(n_629), .Y(n_625) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_644), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_634), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_634), .B(n_739), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g842 ( .A1(n_634), .A2(n_755), .B(n_801), .Y(n_842) );
INVx1_ASAP7_75t_L g732 ( .A(n_635), .Y(n_732) );
INVx3_ASAP7_75t_L g750 ( .A(n_635), .Y(n_750) );
AND2x2_ASAP7_75t_L g890 ( .A(n_635), .B(n_665), .Y(n_890) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g746 ( .A(n_636), .Y(n_746) );
OAI21x1_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_638), .B(n_643), .Y(n_636) );
INVx1_ASAP7_75t_L g696 ( .A(n_638), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_643), .Y(n_697) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_645), .B(n_788), .Y(n_870) );
OAI22x1_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_652), .B1(n_659), .B2(n_663), .Y(n_646) );
OR2x2_ASAP7_75t_L g713 ( .A(n_647), .B(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g780 ( .A(n_647), .B(n_781), .Y(n_780) );
OR2x2_ASAP7_75t_L g835 ( .A(n_647), .B(n_719), .Y(n_835) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g757 ( .A(n_648), .B(n_715), .Y(n_757) );
INVx1_ASAP7_75t_L g885 ( .A(n_648), .Y(n_885) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_654), .B(n_746), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g666 ( .A(n_657), .Y(n_666) );
INVx1_ASAP7_75t_L g729 ( .A(n_658), .Y(n_729) );
OAI221xp5_ASAP7_75t_L g829 ( .A1(n_659), .A2(n_760), .B1(n_775), .B2(n_830), .C(n_832), .Y(n_829) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
AND2x4_ASAP7_75t_L g717 ( .A(n_662), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g741 ( .A(n_662), .B(n_742), .Y(n_741) );
AND2x4_ASAP7_75t_L g761 ( .A(n_664), .B(n_745), .Y(n_761) );
NAND2x1p5_ASAP7_75t_L g876 ( .A(n_664), .B(n_853), .Y(n_876) );
AND2x4_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
AND2x4_ASAP7_75t_L g764 ( .A(n_666), .B(n_695), .Y(n_764) );
OA21x2_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_687), .B(n_689), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
BUFx2_ASAP7_75t_L g739 ( .A(n_671), .Y(n_739) );
AND2x4_ASAP7_75t_L g709 ( .A(n_672), .B(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_673), .Y(n_702) );
INVx2_ASAP7_75t_L g715 ( .A(n_673), .Y(n_715) );
AND2x2_ASAP7_75t_L g742 ( .A(n_673), .B(n_725), .Y(n_742) );
AND2x2_ASAP7_75t_L g767 ( .A(n_673), .B(n_768), .Y(n_767) );
BUFx2_ASAP7_75t_R g882 ( .A(n_673), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_688), .B(n_767), .Y(n_797) );
NAND4xp75_ASAP7_75t_L g689 ( .A(n_690), .B(n_693), .C(n_698), .D(n_700), .Y(n_689) );
INVx2_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g711 ( .A(n_691), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_692), .B(n_750), .Y(n_831) );
OAI32xp33_ASAP7_75t_L g779 ( .A1(n_693), .A2(n_780), .A3(n_782), .B1(n_784), .B2(n_785), .Y(n_779) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g712 ( .A(n_694), .Y(n_712) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND3x1_ASAP7_75t_L g827 ( .A(n_701), .B(n_810), .C(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_733), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
INVx2_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g861 ( .A(n_708), .Y(n_861) );
AND2x2_ASAP7_75t_L g809 ( .A(n_709), .B(n_729), .Y(n_809) );
AND2x2_ASAP7_75t_L g736 ( .A(n_710), .B(n_725), .Y(n_736) );
INVx1_ASAP7_75t_L g864 ( .A(n_710), .Y(n_864) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_712), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g817 ( .A(n_712), .B(n_783), .Y(n_817) );
AND2x2_ASAP7_75t_L g859 ( .A(n_712), .B(n_755), .Y(n_859) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g841 ( .A(n_715), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_720), .B1(n_722), .B2(n_727), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g784 ( .A(n_722), .Y(n_784) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
INVx1_ASAP7_75t_L g753 ( .A(n_724), .Y(n_753) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g737 ( .A(n_726), .Y(n_737) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_728), .B(n_730), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OR2x2_ASAP7_75t_L g777 ( .A(n_729), .B(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_729), .B(n_730), .Y(n_837) );
INVxp67_ASAP7_75t_SL g833 ( .A(n_730), .Y(n_833) );
INVx3_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g828 ( .A(n_731), .B(n_739), .Y(n_828) );
NOR3xp33_ASAP7_75t_L g850 ( .A(n_731), .B(n_846), .C(n_851), .Y(n_850) );
OAI221xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_738), .B1(n_740), .B2(n_743), .C(n_747), .Y(n_733) );
INVxp67_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
AND2x2_ASAP7_75t_L g839 ( .A(n_736), .B(n_840), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_740), .A2(n_837), .B1(n_838), .B2(n_842), .Y(n_836) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g781 ( .A(n_742), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVx1_ASAP7_75t_L g802 ( .A(n_744), .Y(n_802) );
NOR2xp67_ASAP7_75t_L g820 ( .A(n_744), .B(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_745), .B(n_820), .Y(n_819) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_752), .B1(n_755), .B2(n_757), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx3_ASAP7_75t_L g789 ( .A(n_750), .Y(n_789) );
AND2x2_ASAP7_75t_L g873 ( .A(n_750), .B(n_866), .Y(n_873) );
AND2x2_ASAP7_75t_L g887 ( .A(n_750), .B(n_763), .Y(n_887) );
AND2x2_ASAP7_75t_L g799 ( .A(n_751), .B(n_789), .Y(n_799) );
AND2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
OR2x2_ASAP7_75t_L g855 ( .A(n_753), .B(n_766), .Y(n_855) );
BUFx2_ASAP7_75t_L g774 ( .A(n_754), .Y(n_774) );
AND2x2_ASAP7_75t_L g857 ( .A(n_755), .B(n_764), .Y(n_857) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_765), .B1(n_772), .B2(n_776), .C(n_779), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_762), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx2_ASAP7_75t_L g778 ( .A(n_764), .Y(n_778) );
INVx2_ASAP7_75t_SL g847 ( .A(n_764), .Y(n_847) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_769), .Y(n_765) );
OR2x2_ASAP7_75t_L g822 ( .A(n_766), .B(n_769), .Y(n_822) );
INVx2_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
AND2x4_ASAP7_75t_L g790 ( .A(n_767), .B(n_791), .Y(n_790) );
INVxp67_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVxp67_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
BUFx3_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_784), .B(n_813), .Y(n_812) );
AND2x2_ASAP7_75t_L g808 ( .A(n_789), .B(n_809), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_789), .B(n_852), .Y(n_851) );
OAI21xp5_ASAP7_75t_L g823 ( .A1(n_790), .A2(n_805), .B(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
BUFx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_798), .B1(n_800), .B2(n_804), .Y(n_796) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
AND2x4_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NAND4xp25_ASAP7_75t_L g806 ( .A(n_807), .B(n_826), .C(n_843), .D(n_868), .Y(n_806) );
AOI221x1_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_810), .B1(n_812), .B2(n_816), .C(n_818), .Y(n_807) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
OAI21xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_822), .B(n_823), .Y(n_818) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
NOR3xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_829), .C(n_836), .Y(n_826) );
BUFx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
OAI21xp33_ASAP7_75t_SL g844 ( .A1(n_838), .A2(n_845), .B(n_848), .Y(n_844) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_840), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_841), .B(n_864), .Y(n_863) );
AOI21xp33_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_849), .B(n_854), .Y(n_843) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVxp67_ASAP7_75t_SL g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
OAI221xp5_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_856), .B1(n_858), .B2(n_860), .C(n_865), .Y(n_854) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx2_ASAP7_75t_SL g858 ( .A(n_859), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .Y(n_860) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
O2A1O1Ixp5_ASAP7_75t_L g868 ( .A1(n_869), .A2(n_871), .B(n_874), .C(n_875), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
OAI211xp5_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_877), .B(n_879), .C(n_888), .Y(n_875) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
OAI21xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_883), .B(n_887), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
OR2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_886), .Y(n_884) );
INVx2_ASAP7_75t_SL g892 ( .A(n_893), .Y(n_892) );
BUFx8_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_894), .Y(n_899) );
NAND2x1p5_ASAP7_75t_SL g896 ( .A(n_897), .B(n_901), .Y(n_896) );
OR2x2_ASAP7_75t_L g897 ( .A(n_898), .B(n_900), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
BUFx12f_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
CKINVDCx11_ASAP7_75t_R g904 ( .A(n_905), .Y(n_904) );
NOR2xp33_ASAP7_75t_L g907 ( .A(n_908), .B(n_909), .Y(n_907) );
CKINVDCx5p33_ASAP7_75t_R g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVxp67_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
AOI21xp5_ASAP7_75t_L g926 ( .A1(n_913), .A2(n_927), .B(n_928), .Y(n_926) );
NOR2xp33_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .Y(n_913) );
BUFx6f_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
BUFx8_ASAP7_75t_SL g927 ( .A(n_916), .Y(n_927) );
BUFx6f_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
CKINVDCx20_ASAP7_75t_R g919 ( .A(n_920), .Y(n_919) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_921), .Y(n_920) );
NOR2xp67_ASAP7_75t_L g925 ( .A(n_921), .B(n_926), .Y(n_925) );
BUFx8_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
CKINVDCx6p67_ASAP7_75t_R g923 ( .A(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx1_ASAP7_75t_SL g934 ( .A(n_935), .Y(n_934) );
BUFx5_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
INVx1_ASAP7_75t_L g943 ( .A(n_936), .Y(n_943) );
BUFx3_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
OR2x2_ASAP7_75t_L g937 ( .A(n_938), .B(n_941), .Y(n_937) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
endmodule