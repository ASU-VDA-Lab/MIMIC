module real_jpeg_24962_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_0),
.A2(n_26),
.B1(n_31),
.B2(n_73),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_0),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_0),
.A2(n_54),
.B1(n_55),
.B2(n_73),
.Y(n_86)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_2),
.B(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_2),
.B(n_55),
.C(n_57),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_2),
.A2(n_40),
.B1(n_44),
.B2(n_50),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_2),
.B(n_81),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_2),
.A2(n_44),
.B1(n_54),
.B2(n_55),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_2),
.B(n_26),
.C(n_89),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_2),
.A2(n_25),
.B(n_152),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_3),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_4),
.A2(n_40),
.B1(n_50),
.B2(n_61),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_4),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_4),
.A2(n_54),
.B1(n_55),
.B2(n_61),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_4),
.A2(n_26),
.B1(n_31),
.B2(n_61),
.Y(n_165)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_7),
.A2(n_40),
.B1(n_50),
.B2(n_83),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_7),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_7),
.A2(n_54),
.B1(n_55),
.B2(n_83),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_7),
.A2(n_26),
.B1(n_31),
.B2(n_83),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_10),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_12),
.A2(n_26),
.B1(n_31),
.B2(n_36),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_13),
.A2(n_40),
.B1(n_50),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_13),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_13),
.A2(n_54),
.B1(n_55),
.B2(n_64),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_13),
.A2(n_64),
.B1(n_101),
.B2(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_13),
.A2(n_26),
.B1(n_31),
.B2(n_64),
.Y(n_124)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_14),
.Y(n_122)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_14),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_127),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_125),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_105),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_18),
.B(n_105),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_76),
.B2(n_77),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_51),
.B1(n_74),
.B2(n_75),
.Y(n_20)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_37),
.B2(n_38),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_33),
.B2(n_35),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_24),
.A2(n_164),
.B1(n_166),
.B2(n_168),
.Y(n_163)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_25),
.A2(n_30),
.B1(n_34),
.B2(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_25),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_25),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_26),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_26),
.A2(n_31),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_28),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_28),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_31),
.B(n_179),
.Y(n_178)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_34),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B(n_43),
.C(n_47),
.Y(n_38)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_40),
.B1(n_48),
.B2(n_50),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_39),
.A2(n_48),
.B1(n_49),
.B2(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_50),
.B1(n_57),
.B2(n_58),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_40),
.B(n_118),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_SL g100 ( 
.A1(n_43),
.A2(n_44),
.B(n_101),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_44),
.B(n_87),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_44),
.B(n_180),
.Y(n_179)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.C(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_68),
.C(n_71),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_59),
.B(n_62),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_55),
.B1(n_88),
.B2(n_89),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_55),
.B(n_160),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_65),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_63),
.B(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_66),
.A2(n_136),
.B(n_137),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_71),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_94),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_90),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_87),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_87),
.A2(n_90),
.B(n_133),
.Y(n_149)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_113),
.B1(n_115),
.B2(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_100),
.B(n_102),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_116),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_107),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_116),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B(n_114),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_111),
.A2(n_114),
.B(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_119),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B(n_123),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_124),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_141),
.B(n_192),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_138),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_129),
.B(n_138),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.C(n_134),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_130),
.B(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_131),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_186),
.B(n_191),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_161),
.B(n_185),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_155),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_155),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_150),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_149),
.C(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_171),
.B(n_184),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_169),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_169),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_177),
.B(n_183),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_174),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.Y(n_177)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_190),
.Y(n_191)
);


endmodule