module fake_jpeg_13866_n_210 (n_13, n_21, n_57, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_56, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_210);

input n_13;
input n_21;
input n_57;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_56;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_210;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_21),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_11),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_14),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_3),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_28),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_3),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_42),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_31),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_30),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_72),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_94),
.A2(n_77),
.B1(n_68),
.B2(n_65),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_92),
.B1(n_90),
.B2(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_104),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_59),
.B1(n_85),
.B2(n_62),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_65),
.B1(n_68),
.B2(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_79),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_74),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_92),
.B1(n_90),
.B2(n_87),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_80),
.B(n_71),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_125),
.B1(n_129),
.B2(n_130),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_101),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_114),
.Y(n_136)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_118),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_72),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_81),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_121),
.Y(n_145)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_69),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_106),
.A2(n_59),
.B1(n_85),
.B2(n_62),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_84),
.B1(n_82),
.B2(n_67),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_61),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_138),
.C(n_147),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_130),
.A2(n_63),
.B1(n_78),
.B2(n_76),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_141),
.B1(n_0),
.B2(n_1),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_64),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_86),
.B1(n_75),
.B2(n_70),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_128),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_66),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_143),
.B(n_149),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_114),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_23),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_0),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_150),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_22),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_152),
.A2(n_125),
.B1(n_80),
.B2(n_2),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_164),
.B1(n_167),
.B2(n_8),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_157),
.Y(n_181)
);

AO22x1_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_32),
.B1(n_55),
.B2(n_54),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_57),
.B(n_53),
.C(n_52),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_34),
.B(n_33),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_148),
.A2(n_51),
.B1(n_48),
.B2(n_47),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_160),
.A2(n_145),
.B1(n_39),
.B2(n_36),
.Y(n_176)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_166),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_140),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_160),
.Y(n_177)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_147),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_151),
.B(n_144),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_168),
.A2(n_171),
.B(n_35),
.Y(n_179)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_133),
.A2(n_45),
.B1(n_43),
.B2(n_40),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_173),
.A2(n_138),
.B1(n_10),
.B2(n_11),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_131),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_175),
.B(n_180),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_176),
.A2(n_177),
.B1(n_182),
.B2(n_158),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_185),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_9),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_187),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_12),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_12),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_161),
.B1(n_157),
.B2(n_171),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_190),
.A2(n_187),
.B1(n_185),
.B2(n_184),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_178),
.A2(n_163),
.B1(n_174),
.B2(n_157),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_163),
.B(n_174),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_183),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_176),
.B1(n_186),
.B2(n_16),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_197),
.B(n_199),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_194),
.B(n_191),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_194),
.C(n_198),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_202),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_196),
.C(n_198),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_196),
.B(n_189),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_192),
.C(n_15),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_13),
.C(n_17),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_208),
.A2(n_17),
.B(n_18),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_209),
.B(n_18),
.Y(n_210)
);


endmodule