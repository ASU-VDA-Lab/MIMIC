module fake_jpeg_16872_n_267 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_267);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_267;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_11),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_41),
.B(n_60),
.Y(n_97)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_66),
.Y(n_67)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_29),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_18),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_22),
.B1(n_36),
.B2(n_32),
.Y(n_85)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_4),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_4),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_34),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_68),
.B(n_75),
.Y(n_145)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_82),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_66),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_101),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_22),
.B1(n_36),
.B2(n_32),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_20),
.B1(n_8),
.B2(n_9),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_31),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_85),
.A2(n_93),
.B1(n_9),
.B2(n_10),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_35),
.B1(n_38),
.B2(n_31),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_86),
.A2(n_106),
.B1(n_24),
.B2(n_21),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_34),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_91),
.Y(n_121)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_30),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_99),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_30),
.B1(n_27),
.B2(n_26),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

CKINVDCx6p67_ASAP7_75t_R g98 ( 
.A(n_42),
.Y(n_98)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_46),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_19),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_56),
.B(n_19),
.Y(n_102)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_39),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_107),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_13),
.B(n_14),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_50),
.A2(n_38),
.B1(n_35),
.B2(n_23),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_24),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_123),
.Y(n_146)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_113),
.A2(n_134),
.B1(n_143),
.B2(n_140),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_38),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_140),
.B1(n_79),
.B2(n_100),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_38),
.C(n_21),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_115),
.B(n_126),
.Y(n_151)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_119),
.A2(n_127),
.B(n_108),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_68),
.Y(n_123)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_130),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_86),
.A2(n_106),
.B1(n_77),
.B2(n_81),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_141),
.B1(n_109),
.B2(n_111),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_71),
.C(n_74),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_80),
.B(n_5),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_83),
.B(n_20),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_73),
.B(n_75),
.Y(n_150)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_8),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_132),
.Y(n_149)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_138),
.Y(n_167)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_95),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_84),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_15),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_78),
.B(n_104),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_79),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_108),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_147),
.B(n_155),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_100),
.B1(n_73),
.B2(n_88),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_148),
.A2(n_153),
.B1(n_158),
.B2(n_162),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_157),
.B(n_162),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_154),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_125),
.A2(n_88),
.B1(n_123),
.B2(n_122),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_161),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_116),
.B(n_109),
.Y(n_161)
);

OAI22x1_ASAP7_75t_SL g162 ( 
.A1(n_114),
.A2(n_143),
.B1(n_113),
.B2(n_128),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_170),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_114),
.B1(n_137),
.B2(n_139),
.Y(n_166)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_121),
.Y(n_170)
);

O2A1O1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_114),
.A2(n_144),
.B(n_135),
.C(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_115),
.B1(n_118),
.B2(n_126),
.Y(n_172)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_116),
.B1(n_120),
.B2(n_132),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_158),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_110),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_176),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_112),
.A2(n_138),
.B1(n_124),
.B2(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_112),
.B(n_117),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_117),
.B(n_116),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_161),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_196),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_174),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_191),
.C(n_175),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_148),
.B1(n_160),
.B2(n_176),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_169),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_187),
.B(n_188),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_146),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_189),
.A2(n_195),
.B(n_164),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_159),
.C(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_170),
.C(n_149),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_149),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_197),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_171),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_199),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_160),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_153),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_202),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_152),
.B(n_150),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_154),
.B1(n_157),
.B2(n_166),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_186),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_200),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_219),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_167),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_211),
.C(n_218),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_165),
.B1(n_156),
.B2(n_167),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_214),
.C(n_204),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_165),
.C(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_180),
.B(n_201),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_221),
.A2(n_180),
.B(n_198),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_182),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_204),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_190),
.C(n_182),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_190),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_231),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_235),
.C(n_211),
.Y(n_244)
);

AO22x1_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_181),
.B1(n_203),
.B2(n_185),
.Y(n_229)
);

BUFx24_ASAP7_75t_SL g231 ( 
.A(n_224),
.Y(n_231)
);

OAI322xp33_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_195),
.A3(n_187),
.B1(n_178),
.B2(n_181),
.C1(n_203),
.C2(n_193),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_216),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_193),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_234),
.B(n_240),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_183),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_238),
.B(n_226),
.Y(n_243)
);

BUFx12_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_239),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_243),
.C(n_246),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_247),
.C(n_227),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_218),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_222),
.C(n_220),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_217),
.B(n_209),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_229),
.B(n_228),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_250),
.A2(n_252),
.B(n_255),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_237),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_254),
.C(n_256),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_244),
.C(n_247),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_230),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_248),
.A2(n_235),
.B1(n_213),
.B2(n_210),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_239),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_259),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_255),
.A2(n_243),
.B(n_241),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_245),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_212),
.B(n_239),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_253),
.C(n_254),
.Y(n_262)
);

AND2x4_ASAP7_75t_SL g265 ( 
.A(n_262),
.B(n_263),
.Y(n_265)
);

AO21x1_ASAP7_75t_L g266 ( 
.A1(n_265),
.A2(n_264),
.B(n_260),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_266),
.Y(n_267)
);


endmodule