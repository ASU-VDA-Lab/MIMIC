module fake_jpeg_3417_n_109 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_1),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_17),
.B1(n_21),
.B2(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_28),
.Y(n_43)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_16),
.Y(n_38)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_36),
.B1(n_41),
.B2(n_26),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_38),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_17),
.B1(n_15),
.B2(n_13),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_21),
.B1(n_14),
.B2(n_13),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_29),
.A2(n_11),
.B1(n_18),
.B2(n_19),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_48),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_23),
.B1(n_26),
.B2(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_54),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_52),
.Y(n_59)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_26),
.B1(n_30),
.B2(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_58),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_30),
.A3(n_28),
.B1(n_16),
.B2(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_11),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_33),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_33),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_24),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_25),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_34),
.C(n_27),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_24),
.C(n_27),
.Y(n_81)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_54),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_72),
.B(n_75),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_57),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_44),
.B(n_59),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_80),
.B1(n_82),
.B2(n_42),
.Y(n_87)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_84),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_50),
.B1(n_62),
.B2(n_40),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_72),
.A3(n_69),
.B1(n_73),
.B2(n_66),
.C(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_5),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_86),
.B1(n_18),
.B2(n_37),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_76),
.B1(n_78),
.B2(n_37),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_42),
.C(n_37),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_91),
.C(n_81),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_37),
.C(n_25),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_93),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_37),
.A3(n_12),
.B1(n_6),
.B2(n_8),
.C1(n_10),
.C2(n_5),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_88),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_96),
.C(n_97),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_12),
.C(n_18),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_4),
.Y(n_103)
);

AOI21x1_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_91),
.B(n_12),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_100),
.B(n_101),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_97),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_104),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_12),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_12),
.Y(n_107)
);

AOI21x1_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_105),
.B(n_100),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_102),
.Y(n_109)
);


endmodule