module fake_jpeg_512_n_512 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_512);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_512;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_20),
.B(n_14),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_47),
.B(n_58),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_20),
.B(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_51),
.B(n_82),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_31),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_53),
.B(n_60),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_56),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_28),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_31),
.Y(n_59)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_30),
.B(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_19),
.B(n_0),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_62),
.B(n_77),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_68),
.Y(n_154)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_72),
.Y(n_140)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_18),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_13),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_83),
.B(n_91),
.Y(n_144)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_34),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_87),
.B(n_92),
.Y(n_142)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_16),
.Y(n_88)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_90),
.Y(n_128)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_41),
.B(n_29),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_94),
.Y(n_107)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_34),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_97),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_24),
.B(n_13),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_98),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_29),
.B(n_13),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_29),
.C(n_34),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_100),
.B(n_59),
.C(n_66),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_19),
.B1(n_45),
.B2(n_42),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_101),
.A2(n_126),
.B1(n_130),
.B2(n_137),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_69),
.A2(n_46),
.B1(n_45),
.B2(n_42),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_105),
.A2(n_135),
.B1(n_152),
.B2(n_76),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_60),
.B(n_22),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_106),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_85),
.B(n_46),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_117),
.B(n_145),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_84),
.A2(n_19),
.B1(n_45),
.B2(n_42),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_88),
.A2(n_46),
.B1(n_36),
.B2(n_15),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g134 ( 
.A1(n_50),
.A2(n_56),
.A3(n_62),
.B1(n_53),
.B2(n_94),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_83),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_74),
.A2(n_36),
.B1(n_15),
.B2(n_44),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_48),
.A2(n_36),
.B1(n_15),
.B2(n_44),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_147),
.B1(n_22),
.B2(n_25),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_77),
.A2(n_17),
.B1(n_43),
.B2(n_39),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_52),
.A2(n_44),
.B1(n_17),
.B2(n_22),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_156),
.B1(n_32),
.B2(n_37),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_86),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_54),
.A2(n_17),
.B1(n_39),
.B2(n_38),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_75),
.A2(n_43),
.B1(n_39),
.B2(n_38),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_71),
.A2(n_34),
.B1(n_38),
.B2(n_37),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_32),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_61),
.A2(n_43),
.B1(n_37),
.B2(n_32),
.Y(n_156)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_159),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_150),
.Y(n_214)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_162),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_142),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_183),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_106),
.B(n_89),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_164),
.B(n_173),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_165),
.A2(n_166),
.B1(n_178),
.B2(n_205),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_72),
.B1(n_68),
.B2(n_63),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_65),
.B1(n_78),
.B2(n_90),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_167),
.A2(n_168),
.B1(n_200),
.B2(n_129),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_113),
.Y(n_169)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_107),
.B(n_67),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_171),
.B(n_172),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_121),
.B(n_49),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_106),
.B(n_25),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

AO22x1_ASAP7_75t_L g232 ( 
.A1(n_175),
.A2(n_203),
.B1(n_122),
.B2(n_140),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_100),
.B(n_25),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_177),
.B(n_187),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_120),
.A2(n_81),
.B1(n_70),
.B2(n_79),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_120),
.B(n_83),
.Y(n_179)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_179),
.B(n_118),
.Y(n_234)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_184),
.A2(n_186),
.B(n_198),
.Y(n_224)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_127),
.A2(n_73),
.B(n_57),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_120),
.B(n_1),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_153),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_190),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_127),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_124),
.B(n_151),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_191),
.B(n_202),
.Y(n_216)
);

BUFx4f_ASAP7_75t_SL g192 ( 
.A(n_148),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_196),
.Y(n_228)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_193),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_99),
.B(n_64),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_194),
.B(n_195),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_108),
.B(n_55),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_144),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_144),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_197),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_144),
.A2(n_73),
.B(n_27),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_199),
.A2(n_201),
.B1(n_119),
.B2(n_169),
.Y(n_219)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_104),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_103),
.B(n_97),
.Y(n_202)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_155),
.A2(n_23),
.B1(n_92),
.B2(n_27),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_1),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_204),
.B(n_1),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_134),
.A2(n_23),
.B1(n_27),
.B2(n_12),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_186),
.A2(n_114),
.B(n_128),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_206),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_179),
.C(n_190),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_175),
.A2(n_156),
.B1(n_139),
.B2(n_149),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_215),
.A2(n_217),
.B1(n_230),
.B2(n_239),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_161),
.B(n_138),
.CI(n_149),
.CON(n_218),
.SN(n_218)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_214),
.C(n_164),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_219),
.A2(n_225),
.B1(n_178),
.B2(n_176),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_175),
.A2(n_112),
.B1(n_123),
.B2(n_115),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_222),
.A2(n_166),
.B1(n_217),
.B2(n_225),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_196),
.A2(n_122),
.B1(n_111),
.B2(n_139),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_131),
.B1(n_154),
.B2(n_146),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_234),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_233),
.B(n_204),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_160),
.A2(n_133),
.B(n_157),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_203),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_184),
.A2(n_131),
.B1(n_154),
.B2(n_146),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_177),
.B(n_157),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_173),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_214),
.C(n_234),
.Y(n_273)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_245),
.B(n_248),
.Y(n_286)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_246),
.Y(n_299)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_247),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_213),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_253),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_237),
.B(n_182),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_250),
.B(n_252),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_171),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_251),
.B(n_263),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_170),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_170),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_240),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_163),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_258),
.Y(n_277)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_213),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_197),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_261),
.Y(n_288)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_260),
.Y(n_302)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_262),
.A2(n_269),
.B(n_236),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_228),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_221),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_264),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_241),
.B(n_182),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_240),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_210),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_267),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_179),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_272),
.B1(n_232),
.B2(n_224),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_209),
.A2(n_184),
.B1(n_168),
.B2(n_194),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_271),
.A2(n_209),
.B1(n_211),
.B2(n_222),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_217),
.A2(n_165),
.B1(n_203),
.B2(n_198),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_284),
.C(n_290),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_276),
.A2(n_280),
.B1(n_282),
.B2(n_287),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_278),
.B(n_281),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_279),
.A2(n_289),
.B(n_296),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_222),
.B1(n_230),
.B2(n_211),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_242),
.A2(n_218),
.B1(n_232),
.B2(n_226),
.Y(n_282)
);

OAI32xp33_ASAP7_75t_L g283 ( 
.A1(n_251),
.A2(n_226),
.A3(n_218),
.B1(n_231),
.B2(n_215),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_255),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_243),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_270),
.A2(n_258),
.B(n_249),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_231),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_272),
.A2(n_232),
.B1(n_224),
.B2(n_215),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_294),
.A2(n_303),
.B1(n_239),
.B2(n_203),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_263),
.A2(n_256),
.B(n_261),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_250),
.B(n_216),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_298),
.C(n_300),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_218),
.C(n_216),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_245),
.B(n_187),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_242),
.A2(n_239),
.B1(n_236),
.B2(n_233),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_304),
.B(n_309),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_259),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_316),
.C(n_318),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_256),
.B(n_262),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_307),
.A2(n_313),
.B(n_317),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_253),
.Y(n_308)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_293),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_310),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_SL g313 ( 
.A1(n_282),
.A2(n_256),
.B(n_268),
.C(n_259),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_248),
.Y(n_314)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_314),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_293),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_322),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_273),
.B(n_259),
.C(n_267),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_289),
.A2(n_256),
.B(n_206),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_267),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_274),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_319),
.B(n_181),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_288),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_278),
.B(n_267),
.C(n_234),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_323),
.B(n_330),
.C(n_291),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_295),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_324),
.Y(n_366)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_299),
.Y(n_325)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_325),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_279),
.A2(n_206),
.B(n_223),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_326),
.Y(n_352)
);

OAI21xp33_ASAP7_75t_L g327 ( 
.A1(n_292),
.A2(n_252),
.B(n_191),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_327),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_286),
.B(n_221),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_328),
.B(n_302),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_329),
.A2(n_212),
.B1(n_208),
.B2(n_192),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_290),
.B(n_195),
.C(n_202),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_299),
.Y(n_331)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_301),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_332),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_287),
.A2(n_223),
.B(n_219),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_333),
.Y(n_350)
);

MAJx2_ASAP7_75t_L g334 ( 
.A(n_297),
.B(n_172),
.C(n_244),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_334),
.B(n_291),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_288),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_335),
.B(n_266),
.Y(n_358)
);

FAx1_ASAP7_75t_SL g338 ( 
.A(n_307),
.B(n_292),
.CI(n_281),
.CON(n_338),
.SN(n_338)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_338),
.B(n_343),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_320),
.A2(n_276),
.B1(n_303),
.B2(n_294),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_339),
.A2(n_351),
.B1(n_357),
.B2(n_363),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_320),
.A2(n_283),
.B1(n_286),
.B2(n_288),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_341),
.A2(n_348),
.B1(n_359),
.B2(n_364),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_314),
.B(n_300),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_344),
.B(n_347),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_308),
.B(n_280),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_329),
.A2(n_291),
.B1(n_285),
.B2(n_302),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_321),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_353),
.B(n_355),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_333),
.A2(n_285),
.B1(n_301),
.B2(n_246),
.Y(n_357)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_358),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_304),
.A2(n_266),
.B1(n_264),
.B2(n_203),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_305),
.B(n_235),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_360),
.B(n_362),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_305),
.B(n_235),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_326),
.A2(n_264),
.B1(n_260),
.B2(n_247),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_365),
.A2(n_343),
.B1(n_346),
.B2(n_336),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_350),
.A2(n_322),
.B1(n_335),
.B2(n_321),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_370),
.A2(n_373),
.B1(n_376),
.B2(n_379),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_344),
.B(n_330),
.Y(n_371)
);

NAND3xp33_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_388),
.C(n_392),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_362),
.B(n_318),
.C(n_316),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_382),
.C(n_394),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_339),
.A2(n_317),
.B1(n_313),
.B2(n_315),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_345),
.Y(n_374)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_374),
.Y(n_398)
);

OAI21xp33_ASAP7_75t_L g375 ( 
.A1(n_336),
.A2(n_323),
.B(n_311),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_375),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_352),
.A2(n_313),
.B1(n_332),
.B2(n_310),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_361),
.B(n_331),
.Y(n_378)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_378),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_347),
.A2(n_313),
.B1(n_325),
.B2(n_306),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_311),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_380),
.B(n_338),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_342),
.B(n_312),
.C(n_334),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_345),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_383),
.B(n_393),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_361),
.B(n_324),
.Y(n_385)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_385),
.Y(n_408)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_349),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_386),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_354),
.A2(n_313),
.B(n_312),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_387),
.A2(n_338),
.B(n_355),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_346),
.B(n_212),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_390),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_340),
.A2(n_257),
.B1(n_208),
.B2(n_201),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_391),
.B(n_378),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_353),
.B(n_207),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_227),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_174),
.C(n_185),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_352),
.A2(n_201),
.B1(n_188),
.B2(n_199),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_395),
.A2(n_359),
.B1(n_348),
.B2(n_366),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_381),
.B(n_389),
.Y(n_399)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_399),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_368),
.A2(n_357),
.B1(n_367),
.B2(n_363),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_401),
.A2(n_405),
.B1(n_406),
.B2(n_419),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_383),
.A2(n_367),
.B1(n_337),
.B2(n_356),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_385),
.B(n_337),
.Y(n_407)
);

INVxp33_ASAP7_75t_L g437 ( 
.A(n_407),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_410),
.A2(n_386),
.B1(n_376),
.B2(n_370),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_416),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_356),
.Y(n_414)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_414),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_396),
.B(n_349),
.Y(n_415)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_415),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_380),
.B(n_227),
.Y(n_417)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_417),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_394),
.B(n_227),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_418),
.B(n_377),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_368),
.A2(n_192),
.B1(n_123),
.B2(n_115),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_369),
.B(n_207),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_404),
.Y(n_439)
);

FAx1_ASAP7_75t_SL g421 ( 
.A(n_387),
.B(n_192),
.CI(n_210),
.CON(n_421),
.SN(n_421)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_421),
.A2(n_180),
.B1(n_116),
.B2(n_193),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_372),
.C(n_369),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_423),
.B(n_425),
.Y(n_459)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_424),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_403),
.B(n_377),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_416),
.C(n_420),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_428),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_409),
.A2(n_374),
.B1(n_384),
.B2(n_373),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_427),
.A2(n_429),
.B1(n_431),
.B2(n_435),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_382),
.C(n_379),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_395),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_430),
.B(n_102),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_401),
.A2(n_104),
.B1(n_112),
.B2(n_140),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_162),
.C(n_159),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_434),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_133),
.C(n_111),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_398),
.A2(n_176),
.B(n_118),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_439),
.B(n_442),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_433),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_443),
.B(n_453),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_423),
.B(n_407),
.C(n_408),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_447),
.C(n_450),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_407),
.C(n_408),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_441),
.A2(n_404),
.B1(n_398),
.B2(n_397),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_448),
.A2(n_452),
.B1(n_456),
.B2(n_442),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_405),
.C(n_412),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_436),
.A2(n_397),
.B1(n_411),
.B2(n_421),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_412),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_439),
.B(n_419),
.C(n_421),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_454),
.B(n_458),
.C(n_3),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_422),
.B(n_102),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_455),
.B(n_461),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_427),
.A2(n_183),
.B1(n_193),
.B2(n_110),
.Y(n_457)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_457),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_183),
.C(n_110),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_440),
.B(n_183),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_444),
.A2(n_437),
.B(n_432),
.Y(n_462)
);

OAI21x1_ASAP7_75t_SL g482 ( 
.A1(n_462),
.A2(n_475),
.B(n_476),
.Y(n_482)
);

XNOR2x1_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_7),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_431),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_465),
.B(n_467),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_448),
.A2(n_434),
.B1(n_435),
.B2(n_23),
.Y(n_466)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_466),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_23),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_452),
.A2(n_1),
.B(n_2),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_469),
.A2(n_472),
.B(n_473),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_451),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_470)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_470),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_460),
.A2(n_2),
.B(n_3),
.Y(n_472)
);

NAND3xp33_ASAP7_75t_SL g473 ( 
.A(n_445),
.B(n_3),
.C(n_4),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_7),
.Y(n_489)
);

OAI321xp33_ASAP7_75t_L g475 ( 
.A1(n_459),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_9),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_446),
.A2(n_5),
.B(n_7),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_454),
.C(n_444),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_484),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_468),
.B(n_449),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_480),
.B(n_490),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g483 ( 
.A(n_471),
.Y(n_483)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_483),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_474),
.B(n_458),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_469),
.A2(n_7),
.B(n_9),
.Y(n_487)
);

OAI31xp33_ASAP7_75t_L g493 ( 
.A1(n_487),
.A2(n_470),
.A3(n_463),
.B(n_11),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_488),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_489),
.B(n_9),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_477),
.B(n_9),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_481),
.A2(n_462),
.B(n_476),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_492),
.A2(n_486),
.B(n_489),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_493),
.B(n_488),
.Y(n_505)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_494),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_479),
.A2(n_465),
.B(n_467),
.Y(n_498)
);

AOI21x1_ASAP7_75t_L g500 ( 
.A1(n_498),
.A2(n_486),
.B(n_485),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_482),
.A2(n_10),
.B(n_11),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_499),
.B(n_478),
.Y(n_502)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_500),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_495),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_501),
.A2(n_502),
.B(n_505),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_504),
.A2(n_496),
.B(n_497),
.Y(n_508)
);

NAND3xp33_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_491),
.C(n_503),
.Y(n_509)
);

OAI211xp5_ASAP7_75t_L g511 ( 
.A1(n_509),
.A2(n_510),
.B(n_506),
.C(n_10),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_507),
.A2(n_494),
.B(n_10),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_511),
.B(n_11),
.Y(n_512)
);


endmodule