module fake_jpeg_10229_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_40),
.Y(n_48)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_43),
.Y(n_53)
);

HAxp5_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_0),
.CON(n_42),
.SN(n_42)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_19),
.B(n_16),
.Y(n_68)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_58),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_31),
.B1(n_22),
.B2(n_27),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_67),
.B1(n_28),
.B2(n_41),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_42),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_31),
.B1(n_22),
.B2(n_20),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_65),
.A2(n_35),
.B1(n_40),
.B2(n_28),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_46),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_36),
.A2(n_31),
.B1(n_22),
.B2(n_20),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_16),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_43),
.B1(n_39),
.B2(n_31),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_76),
.B1(n_94),
.B2(n_96),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_38),
.B1(n_36),
.B2(n_41),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_35),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_85),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_79),
.A2(n_19),
.B(n_23),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_28),
.B1(n_44),
.B2(n_37),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_87),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_86),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_40),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_53),
.B(n_38),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_38),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_95),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_47),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_46),
.C(n_40),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_17),
.C(n_60),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_46),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_48),
.A2(n_35),
.B1(n_37),
.B2(n_44),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_98),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_57),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_78),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_54),
.Y(n_123)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_106),
.Y(n_139)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

OAI32xp33_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_57),
.A3(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_110)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_110),
.A2(n_17),
.A3(n_73),
.B1(n_32),
.B2(n_18),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_0),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_85),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_119),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_110),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_117),
.C(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_59),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_95),
.C(n_76),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_82),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_84),
.B(n_55),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_74),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_86),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_87),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_117),
.C(n_115),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_132),
.B(n_137),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_85),
.B1(n_75),
.B2(n_55),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_134),
.A2(n_147),
.B1(n_149),
.B2(n_158),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_116),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_136),
.A2(n_138),
.B1(n_21),
.B2(n_32),
.Y(n_192)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_103),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_146),
.Y(n_186)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_148),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_101),
.A2(n_55),
.B1(n_64),
.B2(n_94),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_77),
.B1(n_91),
.B2(n_37),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_74),
.Y(n_150)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_152),
.A2(n_153),
.B(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_73),
.Y(n_154)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_155),
.A2(n_30),
.B1(n_127),
.B2(n_18),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_157),
.B(n_161),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_106),
.A2(n_108),
.B1(n_126),
.B2(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_89),
.Y(n_159)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_109),
.B(n_23),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_164),
.C(n_165),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_133),
.C(n_138),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_107),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_104),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_170),
.B(n_143),
.Y(n_204)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_145),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_107),
.B(n_113),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_107),
.B(n_111),
.Y(n_171)
);

HB1xp67_ASAP7_75t_SL g209 ( 
.A(n_171),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_111),
.C(n_120),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_174),
.C(n_177),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_114),
.C(n_83),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_44),
.C(n_37),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_134),
.A2(n_77),
.B1(n_44),
.B2(n_91),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_178),
.A2(n_183),
.B1(n_190),
.B2(n_191),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_18),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_181),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_147),
.A2(n_59),
.B1(n_127),
.B2(n_29),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_180),
.A2(n_187),
.B1(n_194),
.B2(n_137),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_125),
.C(n_72),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_182),
.A2(n_192),
.B1(n_151),
.B2(n_32),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_141),
.A2(n_30),
.B1(n_34),
.B2(n_125),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_141),
.A2(n_80),
.B1(n_71),
.B2(n_34),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_130),
.A2(n_80),
.B1(n_71),
.B2(n_33),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_130),
.A2(n_71),
.B1(n_33),
.B2(n_24),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_193),
.B(n_195),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_152),
.A2(n_33),
.B1(n_24),
.B2(n_122),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_140),
.B(n_25),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_139),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_196),
.B(n_148),
.Y(n_220)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_203),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_204),
.B(n_186),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_184),
.Y(n_205)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_132),
.Y(n_206)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_206),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_146),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_162),
.C(n_173),
.Y(n_239)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_212),
.Y(n_250)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_213),
.A2(n_216),
.B1(n_221),
.B2(n_182),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_167),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_215),
.Y(n_235)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_170),
.A2(n_155),
.B(n_144),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_217),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_222),
.B1(n_223),
.B2(n_226),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_169),
.A2(n_180),
.B1(n_189),
.B2(n_188),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_163),
.B(n_21),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_178),
.A2(n_146),
.B1(n_122),
.B2(n_33),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_187),
.B1(n_172),
.B2(n_185),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_169),
.A2(n_135),
.B1(n_24),
.B2(n_21),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_231),
.B(n_245),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_234),
.A2(n_237),
.B1(n_246),
.B2(n_247),
.Y(n_273)
);

AOI21x1_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_186),
.B(n_179),
.Y(n_238)
);

AOI22x1_ASAP7_75t_L g263 ( 
.A1(n_238),
.A2(n_231),
.B1(n_216),
.B2(n_235),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_241),
.C(n_251),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_165),
.C(n_177),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_174),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_197),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_212),
.A2(n_183),
.B(n_14),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_213),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_201),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_204),
.A2(n_25),
.B(n_1),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_248),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_25),
.C(n_1),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_210),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_261),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_210),
.C(n_197),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_264),
.C(n_266),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_228),
.B(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_259),
.Y(n_278)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_263),
.B(n_9),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_238),
.C(n_252),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_206),
.C(n_223),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_225),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_269),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_199),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_268),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_226),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_240),
.A2(n_214),
.B1(n_203),
.B2(n_211),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_237),
.B1(n_247),
.B2(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_232),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_230),
.B(n_233),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_218),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_25),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_273),
.A2(n_250),
.B1(n_242),
.B2(n_249),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_274),
.A2(n_286),
.B1(n_8),
.B2(n_2),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_275),
.B(n_280),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_217),
.C(n_214),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_282),
.C(n_283),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_217),
.C(n_236),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_217),
.C(n_236),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_245),
.B1(n_13),
.B2(n_12),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_253),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_25),
.C(n_2),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_253),
.C(n_266),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_288),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_278),
.Y(n_291)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_279),
.A2(n_265),
.B(n_264),
.Y(n_293)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_254),
.C(n_267),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_282),
.C(n_284),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_302),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_283),
.B(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_296),
.B(n_301),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_269),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_303),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_300),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_8),
.Y(n_300)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_0),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_2),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_311),
.A2(n_292),
.B(n_300),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_285),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_3),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_290),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_314),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_277),
.Y(n_314)
);

OAI21xp33_ASAP7_75t_L g316 ( 
.A1(n_295),
.A2(n_285),
.B(n_4),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_316),
.B(n_3),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_318),
.B(n_319),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_301),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_292),
.B(n_4),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_320),
.A2(n_325),
.B(n_5),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_321),
.A2(n_326),
.B1(n_308),
.B2(n_6),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_324),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_4),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_4),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_315),
.A2(n_307),
.B1(n_316),
.B2(n_310),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_328),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_322),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_329),
.A2(n_332),
.B(n_325),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g335 ( 
.A(n_330),
.B(n_5),
.CI(n_6),
.CON(n_335),
.SN(n_335)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_323),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_335),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_331),
.B1(n_333),
.B2(n_332),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_310),
.Y(n_338)
);

AOI322xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_312),
.C1(n_327),
.C2(n_331),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_7),
.B(n_319),
.Y(n_340)
);


endmodule