module fake_netlist_1_12470_n_760 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_760);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_760;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_384;
wire n_227;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_711;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g107 ( .A(n_91), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_7), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_70), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_25), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_84), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_42), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_65), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_34), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_41), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_73), .Y(n_116) );
CKINVDCx14_ASAP7_75t_R g117 ( .A(n_90), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_15), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_104), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_44), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_39), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_5), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_76), .Y(n_123) );
BUFx2_ASAP7_75t_L g124 ( .A(n_71), .Y(n_124) );
CKINVDCx14_ASAP7_75t_R g125 ( .A(n_37), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_100), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_56), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_2), .Y(n_128) );
BUFx3_ASAP7_75t_L g129 ( .A(n_48), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_93), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_72), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_63), .B(n_97), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_12), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_87), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_89), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_9), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_13), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_62), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_46), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_106), .Y(n_140) );
CKINVDCx16_ASAP7_75t_R g141 ( .A(n_49), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_9), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_38), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_53), .Y(n_144) );
INVx1_ASAP7_75t_SL g145 ( .A(n_57), .Y(n_145) );
INVxp33_ASAP7_75t_SL g146 ( .A(n_68), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_103), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_15), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_30), .Y(n_149) );
INVx1_ASAP7_75t_SL g150 ( .A(n_19), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_107), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_119), .B(n_0), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_119), .B(n_124), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_108), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_107), .Y(n_155) );
CKINVDCx6p67_ASAP7_75t_R g156 ( .A(n_141), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_107), .Y(n_157) );
CKINVDCx11_ASAP7_75t_R g158 ( .A(n_111), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_107), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_107), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_107), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_126), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_114), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_128), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_164) );
INVx6_ASAP7_75t_L g165 ( .A(n_114), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_114), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_126), .Y(n_167) );
AND2x6_ASAP7_75t_L g168 ( .A(n_115), .B(n_22), .Y(n_168) );
BUFx12f_ASAP7_75t_L g169 ( .A(n_124), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_120), .Y(n_170) );
NOR3xp33_ASAP7_75t_L g171 ( .A(n_152), .B(n_150), .C(n_122), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_161), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_155), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_155), .Y(n_174) );
NOR2x1p5_ASAP7_75t_L g175 ( .A(n_169), .B(n_118), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_170), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_170), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_157), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_157), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_170), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_163), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_153), .B(n_169), .Y(n_185) );
INVxp67_ASAP7_75t_L g186 ( .A(n_162), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_163), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_163), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_162), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_156), .B(n_141), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_157), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_167), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_167), .A2(n_142), .B1(n_118), .B2(n_108), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_169), .B(n_109), .Y(n_194) );
INVx5_ASAP7_75t_L g195 ( .A(n_168), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_157), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_154), .B(n_110), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_165), .B(n_120), .Y(n_198) );
BUFx4f_ASAP7_75t_L g199 ( .A(n_168), .Y(n_199) );
BUFx4f_ASAP7_75t_L g200 ( .A(n_168), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_199), .B(n_131), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_186), .B(n_156), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_199), .B(n_131), .Y(n_203) );
OAI22xp5_ASAP7_75t_SL g204 ( .A1(n_193), .A2(n_164), .B1(n_130), .B2(n_112), .Y(n_204) );
NAND2xp33_ASAP7_75t_SL g205 ( .A(n_190), .B(n_133), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_186), .B(n_146), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_189), .A2(n_149), .B(n_135), .C(n_143), .Y(n_207) );
INVx8_ASAP7_75t_L g208 ( .A(n_195), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_195), .Y(n_209) );
INVxp67_ASAP7_75t_L g210 ( .A(n_190), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_175), .A2(n_164), .B1(n_136), .B2(n_137), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_197), .B(n_154), .Y(n_212) );
INVxp33_ASAP7_75t_L g213 ( .A(n_171), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_178), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_189), .B(n_168), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_178), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_179), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_192), .B(n_168), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_199), .B(n_116), .Y(n_219) );
OR2x6_ASAP7_75t_L g220 ( .A(n_175), .B(n_142), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_179), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_192), .B(n_168), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_183), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_185), .B(n_154), .Y(n_224) );
OR2x2_ASAP7_75t_L g225 ( .A(n_194), .B(n_148), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_183), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_184), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_198), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_198), .A2(n_154), .B(n_149), .C(n_147), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_184), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_184), .Y(n_231) );
NOR2xp33_ASAP7_75t_SL g232 ( .A(n_199), .B(n_168), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_184), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_200), .B(n_135), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_200), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_195), .B(n_113), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_187), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_200), .A2(n_143), .B(n_144), .C(n_147), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_195), .B(n_165), .Y(n_239) );
O2A1O1Ixp5_ASAP7_75t_L g240 ( .A1(n_200), .A2(n_144), .B(n_138), .C(n_140), .Y(n_240) );
BUFx3_ASAP7_75t_L g241 ( .A(n_195), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_213), .B(n_195), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_228), .B(n_195), .Y(n_243) );
AOI21x1_ASAP7_75t_L g244 ( .A1(n_215), .A2(n_196), .B(n_191), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_223), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_207), .A2(n_117), .B(n_125), .C(n_140), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_218), .A2(n_187), .B(n_188), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_222), .A2(n_187), .B(n_188), .Y(n_248) );
NOR3xp33_ASAP7_75t_L g249 ( .A(n_204), .B(n_158), .C(n_145), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_232), .A2(n_187), .B(n_188), .Y(n_250) );
NAND3xp33_ASAP7_75t_L g251 ( .A(n_206), .B(n_134), .C(n_139), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_210), .A2(n_138), .B(n_121), .C(n_129), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_223), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_214), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_206), .B(n_165), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_202), .B(n_165), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_224), .B(n_123), .Y(n_257) );
O2A1O1Ixp5_ASAP7_75t_L g258 ( .A1(n_240), .A2(n_188), .B(n_132), .C(n_196), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_201), .A2(n_196), .B(n_191), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_225), .B(n_127), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_224), .B(n_163), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_216), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_201), .A2(n_191), .B(n_182), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_217), .A2(n_115), .B1(n_121), .B2(n_129), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_235), .B(n_163), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_203), .A2(n_182), .B(n_181), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_221), .B(n_166), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_238), .A2(n_115), .B(n_121), .C(n_129), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g269 ( .A(n_226), .B(n_166), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_212), .B(n_166), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_203), .A2(n_182), .B(n_181), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_212), .B(n_166), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_211), .A2(n_166), .B1(n_151), .B2(n_157), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_234), .A2(n_219), .B(n_239), .Y(n_274) );
AO32x1_ASAP7_75t_L g275 ( .A1(n_230), .A2(n_151), .A3(n_181), .B1(n_177), .B2(n_176), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_220), .B(n_1), .Y(n_276) );
AO22x2_ASAP7_75t_L g277 ( .A1(n_249), .A2(n_234), .B1(n_220), .B2(n_205), .Y(n_277) );
AND2x2_ASAP7_75t_SL g278 ( .A(n_262), .B(n_235), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_253), .B(n_220), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g280 ( .A1(n_252), .A2(n_229), .B(n_236), .C(n_237), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_262), .B(n_236), .Y(n_281) );
OA21x2_ASAP7_75t_L g282 ( .A1(n_258), .A2(n_151), .B(n_176), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_245), .Y(n_283) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_246), .A2(n_231), .B(n_233), .C(n_227), .Y(n_284) );
BUFx2_ASAP7_75t_L g285 ( .A(n_254), .Y(n_285) );
OAI21xp5_ASAP7_75t_L g286 ( .A1(n_268), .A2(n_233), .B(n_227), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_267), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_270), .Y(n_288) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_260), .A2(n_208), .B1(n_209), .B2(n_241), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_247), .A2(n_208), .B(n_241), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_244), .Y(n_291) );
BUFx12f_ASAP7_75t_L g292 ( .A(n_269), .Y(n_292) );
OAI21x1_ASAP7_75t_L g293 ( .A1(n_250), .A2(n_174), .B(n_180), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_272), .Y(n_294) );
AO21x1_ASAP7_75t_L g295 ( .A1(n_261), .A2(n_174), .B(n_177), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_269), .A2(n_174), .B(n_180), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_260), .B(n_276), .Y(n_297) );
AOI21xp5_ASAP7_75t_SL g298 ( .A1(n_264), .A2(n_209), .B(n_161), .Y(n_298) );
CKINVDCx16_ASAP7_75t_R g299 ( .A(n_273), .Y(n_299) );
OAI21x1_ASAP7_75t_SL g300 ( .A1(n_274), .A2(n_208), .B(n_4), .Y(n_300) );
O2A1O1Ixp33_ASAP7_75t_L g301 ( .A1(n_255), .A2(n_177), .B(n_176), .C(n_173), .Y(n_301) );
NAND2x1p5_ASAP7_75t_L g302 ( .A(n_283), .B(n_265), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_297), .B(n_242), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_285), .Y(n_304) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_293), .A2(n_271), .B(n_266), .Y(n_305) );
OAI21x1_ASAP7_75t_L g306 ( .A1(n_293), .A2(n_263), .B(n_259), .Y(n_306) );
AO31x2_ASAP7_75t_L g307 ( .A1(n_295), .A2(n_256), .A3(n_242), .B(n_248), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_297), .B(n_256), .Y(n_308) );
OAI21xp5_ASAP7_75t_L g309 ( .A1(n_288), .A2(n_265), .B(n_243), .Y(n_309) );
OA21x2_ASAP7_75t_L g310 ( .A1(n_291), .A2(n_275), .B(n_173), .Y(n_310) );
OA21x2_ASAP7_75t_L g311 ( .A1(n_291), .A2(n_275), .B(n_173), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_283), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_283), .Y(n_313) );
AOI22x1_ASAP7_75t_L g314 ( .A1(n_300), .A2(n_160), .B1(n_159), .B2(n_161), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_283), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_292), .Y(n_316) );
OAI21x1_ASAP7_75t_L g317 ( .A1(n_295), .A2(n_275), .B(n_180), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_285), .B(n_251), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_279), .B(n_257), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_288), .Y(n_320) );
NAND3xp33_ASAP7_75t_SL g321 ( .A(n_280), .B(n_3), .C(n_4), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_292), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_294), .B(n_3), .Y(n_323) );
NAND2x1p5_ASAP7_75t_L g324 ( .A(n_278), .B(n_161), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_310), .Y(n_325) );
INVxp67_ASAP7_75t_SL g326 ( .A(n_324), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_303), .B(n_279), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_320), .B(n_294), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_320), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_312), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_310), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_310), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_310), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_312), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_304), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_313), .B(n_282), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_313), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_311), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_303), .A2(n_277), .B1(n_300), .B2(n_287), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_315), .B(n_287), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_324), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_315), .B(n_282), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_323), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_323), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_311), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_311), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_324), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_311), .Y(n_348) );
AO21x2_ASAP7_75t_L g349 ( .A1(n_321), .A2(n_298), .B(n_286), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_308), .B(n_299), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_307), .Y(n_351) );
OAI21x1_ASAP7_75t_L g352 ( .A1(n_317), .A2(n_282), .B(n_298), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_307), .Y(n_353) );
INVx2_ASAP7_75t_SL g354 ( .A(n_316), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_329), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_329), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_328), .B(n_308), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_350), .A2(n_319), .B1(n_277), .B2(n_321), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_328), .B(n_343), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_325), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_328), .B(n_307), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_345), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_351), .B(n_307), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_351), .B(n_307), .Y(n_364) );
AOI22xp33_ASAP7_75t_SL g365 ( .A1(n_350), .A2(n_314), .B1(n_277), .B2(n_322), .Y(n_365) );
INVxp67_ASAP7_75t_L g366 ( .A(n_335), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_345), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_325), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_353), .B(n_307), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_353), .B(n_335), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_330), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_330), .B(n_316), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_325), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_327), .A2(n_277), .B1(n_319), .B2(n_318), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_334), .Y(n_375) );
OR2x2_ASAP7_75t_L g376 ( .A(n_334), .B(n_322), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_336), .B(n_317), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_337), .B(n_309), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_337), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_327), .A2(n_319), .B1(n_322), .B2(n_318), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_336), .B(n_309), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_331), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_331), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_336), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_343), .B(n_319), .Y(n_385) );
INVx3_ASAP7_75t_L g386 ( .A(n_347), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_342), .B(n_317), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_347), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_342), .B(n_302), .Y(n_389) );
NOR2x1_ASAP7_75t_L g390 ( .A(n_347), .B(n_322), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_331), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_347), .Y(n_392) );
AND2x4_ASAP7_75t_SL g393 ( .A(n_341), .B(n_318), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_342), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_332), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_332), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_332), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_344), .B(n_302), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_344), .B(n_302), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_339), .A2(n_318), .B1(n_299), .B2(n_278), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_333), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_347), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_354), .Y(n_403) );
NOR2xp67_ASAP7_75t_L g404 ( .A(n_366), .B(n_354), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_362), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_384), .B(n_333), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_384), .B(n_333), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_403), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_394), .B(n_338), .Y(n_409) );
INVx4_ASAP7_75t_R g410 ( .A(n_402), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_372), .B(n_354), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_360), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_360), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_360), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_369), .B(n_338), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_366), .Y(n_416) );
AOI22xp33_ASAP7_75t_SL g417 ( .A1(n_393), .A2(n_326), .B1(n_341), .B2(n_314), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_394), .B(n_338), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_370), .B(n_346), .Y(n_419) );
NAND2x1_ASAP7_75t_L g420 ( .A(n_362), .B(n_346), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_368), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_377), .B(n_387), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_368), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_377), .B(n_346), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_367), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_359), .B(n_340), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_377), .B(n_348), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_359), .B(n_340), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_370), .B(n_348), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_367), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_357), .B(n_340), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_355), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_387), .B(n_348), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_368), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_355), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_357), .B(n_340), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_356), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_372), .B(n_5), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_387), .B(n_369), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_369), .B(n_339), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_385), .B(n_340), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_361), .B(n_326), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_376), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_390), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_363), .B(n_352), .Y(n_445) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_383), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_385), .B(n_349), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_363), .B(n_352), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_373), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_356), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_364), .B(n_352), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_371), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_371), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_364), .B(n_349), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_361), .B(n_349), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_373), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_381), .B(n_349), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_373), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_389), .B(n_349), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_381), .B(n_383), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_375), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_375), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_389), .B(n_282), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_379), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_391), .B(n_159), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_391), .B(n_159), .Y(n_466) );
NAND2x1_ASAP7_75t_L g467 ( .A(n_386), .B(n_161), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_379), .B(n_6), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_395), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_395), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_382), .B(n_159), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_382), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_382), .B(n_159), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_396), .B(n_160), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_396), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_396), .B(n_6), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_439), .B(n_378), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_416), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_439), .B(n_393), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_422), .B(n_424), .Y(n_480) );
INVxp67_ASAP7_75t_L g481 ( .A(n_446), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_422), .B(n_393), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_432), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_424), .B(n_398), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_440), .B(n_378), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_427), .B(n_398), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_442), .B(n_397), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_427), .B(n_399), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_432), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_435), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_440), .B(n_397), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_435), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_433), .B(n_399), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_433), .B(n_443), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_405), .B(n_397), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_415), .B(n_402), .Y(n_496) );
NOR2x1_ASAP7_75t_SL g497 ( .A(n_476), .B(n_376), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_408), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_405), .B(n_401), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_437), .Y(n_500) );
INVx3_ASAP7_75t_SL g501 ( .A(n_476), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_415), .B(n_402), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_438), .A2(n_374), .B1(n_358), .B2(n_380), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_437), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_425), .B(n_401), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_450), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
AND2x4_ASAP7_75t_SL g508 ( .A(n_415), .B(n_386), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_452), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_442), .B(n_401), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_452), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_453), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_460), .B(n_380), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_468), .B(n_411), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_425), .B(n_430), .Y(n_515) );
BUFx3_ASAP7_75t_L g516 ( .A(n_467), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_431), .A2(n_358), .B1(n_365), .B2(n_400), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_453), .Y(n_518) );
INVxp67_ASAP7_75t_L g519 ( .A(n_420), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_415), .B(n_386), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_420), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_430), .B(n_365), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_461), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_460), .B(n_386), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_404), .B(n_388), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_444), .B(n_388), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_461), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_444), .B(n_388), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_462), .B(n_392), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_413), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_436), .B(n_392), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_462), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_406), .B(n_388), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_464), .Y(n_534) );
NAND2x1p5_ASAP7_75t_L g535 ( .A(n_467), .B(n_390), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_464), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_409), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_406), .B(n_392), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_409), .B(n_392), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_413), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_469), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_407), .B(n_7), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_426), .B(n_8), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_407), .B(n_8), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_413), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_469), .Y(n_546) );
INVx3_ASAP7_75t_L g547 ( .A(n_475), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_470), .B(n_160), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_470), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_419), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_418), .B(n_10), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_457), .B(n_160), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_418), .B(n_305), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_475), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_428), .B(n_10), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_419), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_475), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_457), .B(n_160), .Y(n_558) );
NAND2x1_ASAP7_75t_L g559 ( .A(n_410), .B(n_161), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_429), .B(n_11), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_445), .B(n_11), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_445), .B(n_12), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_429), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_448), .B(n_451), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_480), .B(n_448), .Y(n_565) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_481), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_515), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_485), .B(n_454), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_564), .B(n_451), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_485), .B(n_477), .Y(n_570) );
INVxp67_ASAP7_75t_L g571 ( .A(n_552), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_530), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_494), .B(n_459), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_530), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_515), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_478), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_508), .B(n_459), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_483), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_477), .B(n_455), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_489), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_490), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_491), .B(n_487), .Y(n_582) );
O2A1O1Ixp33_ASAP7_75t_SL g583 ( .A1(n_498), .A2(n_441), .B(n_455), .C(n_447), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_516), .B(n_417), .Y(n_584) );
INVx2_ASAP7_75t_SL g585 ( .A(n_508), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_482), .B(n_459), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_479), .Y(n_587) );
OAI21xp5_ASAP7_75t_L g588 ( .A1(n_561), .A2(n_466), .B(n_465), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_492), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_500), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_484), .B(n_486), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_504), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_506), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_488), .B(n_459), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_514), .B(n_454), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_507), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_522), .B(n_465), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_522), .B(n_466), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_509), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_550), .B(n_463), .Y(n_600) );
OAI221xp5_ASAP7_75t_L g601 ( .A1(n_517), .A2(n_423), .B1(n_412), .B2(n_472), .C(n_414), .Y(n_601) );
AND2x4_ASAP7_75t_SL g602 ( .A(n_496), .B(n_412), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_511), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_493), .B(n_463), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_512), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_556), .B(n_414), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_502), .B(n_520), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_563), .B(n_421), .Y(n_608) );
INVx2_ASAP7_75t_SL g609 ( .A(n_516), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_562), .B(n_491), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_533), .B(n_538), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_518), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_523), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_527), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_532), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_513), .B(n_421), .Y(n_616) );
AND2x4_ASAP7_75t_SL g617 ( .A(n_525), .B(n_423), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_537), .B(n_434), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_481), .B(n_434), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_501), .B(n_449), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_510), .B(n_449), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_501), .B(n_456), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_534), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_536), .Y(n_624) );
NAND2x2_ASAP7_75t_L g625 ( .A(n_559), .B(n_13), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_542), .B(n_456), .Y(n_626) );
OAI21xp33_ASAP7_75t_L g627 ( .A1(n_517), .A2(n_474), .B(n_473), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_541), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_546), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_544), .B(n_458), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_549), .Y(n_631) );
INVxp67_ASAP7_75t_L g632 ( .A(n_552), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_535), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_503), .A2(n_514), .B1(n_543), .B2(n_555), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_548), .Y(n_635) );
INVx1_ASAP7_75t_SL g636 ( .A(n_551), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_560), .B(n_458), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_524), .B(n_472), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_529), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_548), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_529), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_495), .Y(n_642) );
INVx2_ASAP7_75t_SL g643 ( .A(n_602), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_566), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_627), .A2(n_503), .B1(n_553), .B2(n_558), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_636), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_595), .B(n_531), .Y(n_647) );
AOI322xp5_ASAP7_75t_L g648 ( .A1(n_634), .A2(n_558), .A3(n_521), .B1(n_553), .B2(n_519), .C1(n_557), .C2(n_540), .Y(n_648) );
NOR2xp33_ASAP7_75t_SL g649 ( .A(n_609), .B(n_521), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_595), .A2(n_526), .B1(n_528), .B2(n_525), .Y(n_650) );
OAI21xp33_ASAP7_75t_SL g651 ( .A1(n_584), .A2(n_519), .B(n_540), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_639), .B(n_557), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_566), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_641), .B(n_497), .Y(n_654) );
AOI21x1_ASAP7_75t_L g655 ( .A1(n_584), .A2(n_471), .B(n_473), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_571), .B(n_495), .Y(n_656) );
BUFx2_ASAP7_75t_L g657 ( .A(n_585), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_570), .B(n_526), .Y(n_658) );
OAI222xp33_ASAP7_75t_L g659 ( .A1(n_601), .A2(n_535), .B1(n_539), .B2(n_547), .C1(n_528), .C2(n_505), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_571), .B(n_499), .Y(n_660) );
OA21x2_ASAP7_75t_L g661 ( .A1(n_572), .A2(n_505), .B(n_499), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_567), .Y(n_662) );
INVx1_ASAP7_75t_SL g663 ( .A(n_602), .Y(n_663) );
INVxp67_ASAP7_75t_L g664 ( .A(n_576), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_572), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_587), .B(n_547), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_575), .Y(n_667) );
INVxp67_ASAP7_75t_SL g668 ( .A(n_619), .Y(n_668) );
AOI322xp5_ASAP7_75t_L g669 ( .A1(n_634), .A2(n_554), .A3(n_545), .B1(n_474), .B2(n_471), .C1(n_278), .C2(n_20), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_632), .A2(n_305), .B1(n_306), .B2(n_284), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_632), .B(n_14), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_583), .A2(n_275), .B(n_305), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_L g673 ( .A1(n_583), .A2(n_281), .B(n_289), .C(n_301), .Y(n_673) );
OAI31xp33_ASAP7_75t_SL g674 ( .A1(n_577), .A2(n_14), .A3(n_16), .B(n_17), .Y(n_674) );
AOI32xp33_ASAP7_75t_L g675 ( .A1(n_617), .A2(n_306), .A3(n_296), .B1(n_18), .B2(n_19), .Y(n_675) );
INVx1_ASAP7_75t_SL g676 ( .A(n_617), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_642), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_590), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_590), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_569), .B(n_306), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_610), .B(n_16), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_568), .B(n_17), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_603), .Y(n_683) );
OAI21xp33_ASAP7_75t_L g684 ( .A1(n_579), .A2(n_296), .B(n_290), .Y(n_684) );
OAI21xp33_ASAP7_75t_L g685 ( .A1(n_616), .A2(n_18), .B(n_20), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_597), .A2(n_172), .B1(n_21), .B2(n_24), .Y(n_686) );
OAI22xp33_ASAP7_75t_L g687 ( .A1(n_625), .A2(n_21), .B1(n_172), .B2(n_26), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_637), .B(n_23), .Y(n_688) );
INVx1_ASAP7_75t_SL g689 ( .A(n_620), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_L g690 ( .A1(n_633), .A2(n_27), .B(n_28), .C(n_29), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_633), .A2(n_172), .B(n_32), .Y(n_691) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_585), .A2(n_31), .B(n_33), .C(n_35), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_656), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_660), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_651), .A2(n_609), .B(n_633), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_659), .A2(n_637), .B1(n_592), .B2(n_578), .C(n_631), .Y(n_696) );
AOI31xp33_ASAP7_75t_L g697 ( .A1(n_676), .A2(n_588), .A3(n_625), .B(n_622), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_677), .Y(n_698) );
INVxp67_ASAP7_75t_L g699 ( .A(n_681), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_646), .B(n_582), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g701 ( .A(n_648), .B(n_605), .C(n_580), .Y(n_701) );
AOI322xp5_ASAP7_75t_L g702 ( .A1(n_647), .A2(n_565), .A3(n_591), .B1(n_604), .B2(n_573), .C1(n_594), .C2(n_598), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_662), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_649), .B(n_577), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_657), .A2(n_577), .B1(n_640), .B2(n_635), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_667), .Y(n_706) );
OAI332xp33_ASAP7_75t_L g707 ( .A1(n_682), .A2(n_630), .A3(n_626), .B1(n_600), .B2(n_606), .B3(n_608), .C1(n_628), .C2(n_629), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_645), .A2(n_586), .B1(n_581), .B2(n_614), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_668), .Y(n_709) );
AOI221x1_ASAP7_75t_L g710 ( .A1(n_644), .A2(n_615), .B1(n_599), .B2(n_596), .C(n_612), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_664), .A2(n_589), .B1(n_593), .B2(n_604), .C(n_624), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_663), .A2(n_607), .B1(n_611), .B2(n_618), .Y(n_712) );
OAI221xp5_ASAP7_75t_L g713 ( .A1(n_674), .A2(n_603), .B1(n_624), .B2(n_623), .C(n_613), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_649), .A2(n_613), .B(n_623), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_663), .A2(n_621), .B1(n_638), .B2(n_635), .Y(n_715) );
OAI221xp5_ASAP7_75t_SL g716 ( .A1(n_675), .A2(n_640), .B1(n_574), .B2(n_43), .C(n_45), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_676), .A2(n_574), .B1(n_172), .B2(n_47), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_653), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_652), .Y(n_719) );
AOI332xp33_ASAP7_75t_L g720 ( .A1(n_650), .A2(n_36), .A3(n_40), .B1(n_50), .B2(n_51), .B3(n_52), .C1(n_54), .C2(n_55), .Y(n_720) );
O2A1O1Ixp5_ASAP7_75t_L g721 ( .A1(n_695), .A2(n_655), .B(n_687), .C(n_671), .Y(n_721) );
AOI211xp5_ASAP7_75t_L g722 ( .A1(n_713), .A2(n_685), .B(n_643), .C(n_666), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_707), .B(n_658), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_709), .B(n_680), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_697), .A2(n_654), .B1(n_689), .B2(n_679), .C(n_678), .Y(n_725) );
AOI221x1_ASAP7_75t_SL g726 ( .A1(n_701), .A2(n_683), .B1(n_688), .B2(n_665), .C(n_684), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_693), .B(n_669), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g728 ( .A1(n_704), .A2(n_690), .B(n_692), .Y(n_728) );
AOI222xp33_ASAP7_75t_L g729 ( .A1(n_696), .A2(n_661), .B1(n_686), .B2(n_673), .C1(n_670), .C2(n_672), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_694), .B(n_661), .Y(n_730) );
NOR2xp67_ASAP7_75t_L g731 ( .A(n_714), .B(n_691), .Y(n_731) );
INVxp67_ASAP7_75t_L g732 ( .A(n_700), .Y(n_732) );
NOR4xp25_ASAP7_75t_SL g733 ( .A(n_716), .B(n_58), .C(n_59), .D(n_60), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_719), .B(n_61), .Y(n_734) );
AOI222xp33_ASAP7_75t_L g735 ( .A1(n_732), .A2(n_699), .B1(n_711), .B2(n_715), .C1(n_718), .C2(n_703), .Y(n_735) );
NAND4xp25_ASAP7_75t_L g736 ( .A(n_721), .B(n_716), .C(n_699), .D(n_708), .Y(n_736) );
NOR3x1_ASAP7_75t_L g737 ( .A(n_728), .B(n_717), .C(n_706), .Y(n_737) );
NAND3xp33_ASAP7_75t_SL g738 ( .A(n_733), .B(n_720), .C(n_702), .Y(n_738) );
NAND4xp25_ASAP7_75t_L g739 ( .A(n_726), .B(n_705), .C(n_710), .D(n_712), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g740 ( .A1(n_723), .A2(n_698), .B1(n_172), .B2(n_67), .C(n_69), .Y(n_740) );
NAND4xp25_ASAP7_75t_SL g741 ( .A(n_725), .B(n_64), .C(n_66), .D(n_74), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_738), .A2(n_729), .B1(n_731), .B2(n_727), .Y(n_742) );
AOI211xp5_ASAP7_75t_L g743 ( .A1(n_736), .A2(n_722), .B(n_730), .C(n_734), .Y(n_743) );
NAND3xp33_ASAP7_75t_SL g744 ( .A(n_735), .B(n_724), .C(n_77), .Y(n_744) );
OR2x2_ASAP7_75t_L g745 ( .A(n_739), .B(n_75), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g746 ( .A1(n_742), .A2(n_737), .B(n_740), .C(n_741), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_743), .B(n_78), .Y(n_747) );
NOR3xp33_ASAP7_75t_L g748 ( .A(n_745), .B(n_79), .C(n_80), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_747), .Y(n_749) );
AO22x2_ASAP7_75t_L g750 ( .A1(n_748), .A2(n_744), .B1(n_82), .B2(n_83), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_749), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g752 ( .A1(n_750), .A2(n_746), .B1(n_172), .B2(n_86), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_752), .B(n_751), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_751), .B(n_81), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_753), .A2(n_85), .B1(n_88), .B2(n_92), .Y(n_755) );
OAI21xp5_ASAP7_75t_L g756 ( .A1(n_754), .A2(n_94), .B(n_95), .Y(n_756) );
OR2x2_ASAP7_75t_L g757 ( .A(n_755), .B(n_96), .Y(n_757) );
AO21x2_ASAP7_75t_L g758 ( .A1(n_757), .A2(n_756), .B(n_99), .Y(n_758) );
OR2x6_ASAP7_75t_L g759 ( .A(n_758), .B(n_98), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_759), .A2(n_101), .B1(n_102), .B2(n_105), .Y(n_760) );
endmodule