module real_jpeg_702_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_75),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_1),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_75),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_75),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_75),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_2),
.A2(n_52),
.B1(n_63),
.B2(n_64),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_3),
.A2(n_41),
.B1(n_42),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_3),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_122),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_122),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_3),
.A2(n_63),
.B1(n_64),
.B2(n_122),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_4),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_5),
.B(n_53),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_5),
.B(n_26),
.C(n_28),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_5),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_5),
.B(n_25),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_5),
.B(n_60),
.C(n_63),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_211),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_5),
.B(n_112),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_5),
.B(n_65),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_211),
.Y(n_276)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_8),
.A2(n_37),
.B1(n_63),
.B2(n_64),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_44),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_44),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_10),
.A2(n_44),
.B1(n_63),
.B2(n_64),
.Y(n_169)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_13),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_144),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_144),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_144),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_14),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_83),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_83),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_14),
.A2(n_63),
.B1(n_64),
.B2(n_83),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_15),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_176),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_176),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_15),
.A2(n_63),
.B1(n_64),
.B2(n_176),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_89),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_88),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_76),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_56),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_38),
.B1(n_54),
.B2(n_55),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_23),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B(n_35),
.Y(n_23)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_24),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_25),
.B(n_173),
.Y(n_277)
);

AO22x1_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_25)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_27),
.A2(n_28),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_28),
.B(n_250),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_33),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_32),
.B(n_201),
.Y(n_200)
);

NAND2xp33_ASAP7_75t_SL g225 ( 
.A(n_32),
.B(n_48),
.Y(n_225)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

AOI32xp33_ASAP7_75t_L g223 ( 
.A1(n_33),
.A2(n_42),
.A3(n_47),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_36),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_45),
.B1(n_51),
.B2(n_53),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_46),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_50)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_42),
.A2(n_73),
.B(n_211),
.C(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_42),
.B(n_211),
.Y(n_212)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_45),
.B(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_45),
.A2(n_53),
.B1(n_143),
.B2(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_73),
.B1(n_74),
.B2(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_46),
.A2(n_82),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_46),
.B(n_121),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_46),
.A2(n_119),
.B(n_297),
.Y(n_296)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_68),
.C(n_72),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_68),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_81),
.C(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_57),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_65),
.B(n_66),
.Y(n_57)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_58),
.A2(n_65),
.B1(n_117),
.B2(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_58),
.A2(n_65),
.B1(n_138),
.B2(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_58),
.A2(n_193),
.B(n_195),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_58),
.B(n_197),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_67),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_62),
.A2(n_98),
.B1(n_99),
.B2(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_62),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_62),
.A2(n_218),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_62),
.A2(n_98),
.B1(n_194),
.B2(n_244),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_63),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_63),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_65),
.B(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_71),
.B1(n_87),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_69),
.A2(n_71),
.B1(n_96),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_69),
.A2(n_71),
.B1(n_184),
.B2(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_69),
.A2(n_276),
.B(n_277),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_69),
.A2(n_215),
.B(n_277),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_71),
.A2(n_140),
.B(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_71),
.A2(n_172),
.B(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_73),
.A2(n_142),
.B(n_145),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.C(n_84),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_77),
.A2(n_81),
.B1(n_101),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_84),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AO21x1_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_152),
.B(n_325),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_147),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_123),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_92),
.B(n_123),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_104),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_95),
.B(n_97),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_94),
.B(n_100),
.C(n_104),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_98),
.A2(n_196),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B(n_118),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_106),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_115),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_108),
.B1(n_118),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_107),
.A2(n_108),
.B1(n_115),
.B2(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_112),
.B(n_113),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_109),
.A2(n_112),
.B1(n_135),
.B2(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_109),
.A2(n_211),
.B(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_110),
.A2(n_111),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_110),
.B(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_110),
.A2(n_111),
.B1(n_191),
.B2(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_110),
.A2(n_236),
.B(n_237),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_110),
.A2(n_111),
.B1(n_236),
.B2(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_111),
.A2(n_190),
.B(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_111),
.B(n_205),
.Y(n_238)
);

INVx3_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_112),
.A2(n_204),
.B(n_261),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_115),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_118),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.C(n_130),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_125),
.B1(n_129),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_139),
.C(n_141),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_132),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_133),
.A2(n_136),
.B1(n_137),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_133),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_141),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_146),
.B(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_147),
.A2(n_326),
.B(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_148),
.B(n_151),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_177),
.B(n_324),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_154),
.B(n_157),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_163),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_158),
.B(n_161),
.Y(n_322)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_163),
.B(n_322),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.C(n_174),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_164),
.A2(n_165),
.B1(n_312),
.B2(n_314),
.Y(n_311)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_166),
.B(n_168),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_167),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_169),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_174),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_175),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_319),
.B(n_323),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_288),
.B(n_316),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_230),
.B(n_287),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_206),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_181),
.B(n_206),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_192),
.C(n_198),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_182),
.B(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_186),
.C(n_189),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_192),
.B(n_198),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_202),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_220),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_207),
.B(n_221),
.C(n_229),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_213),
.B2(n_219),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_208),
.B(n_214),
.C(n_216),
.Y(n_301)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_212),
.Y(n_224)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_222),
.B(n_227),
.Y(n_292)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_282),
.B(n_286),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_271),
.B(n_281),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_253),
.B(n_270),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_247),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_247),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_239),
.B1(n_245),
.B2(n_246),
.Y(n_234)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_239),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_242),
.C(n_245),
.Y(n_272)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_248),
.A2(n_249),
.B1(n_251),
.B2(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_251),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_264),
.B(n_269),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_259),
.B(n_263),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_262),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_261),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_267),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_273),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_279),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_278),
.C(n_279),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_285),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_303),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_302),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_302),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_299),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_300),
.C(n_301),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_294),
.C(n_298),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_298),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_296),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_315),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_315),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_305),
.B(n_309),
.C(n_311),
.Y(n_320)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_312),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_321),
.Y(n_323)
);


endmodule