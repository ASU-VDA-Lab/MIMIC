module fake_jpeg_31166_n_177 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_17),
.A2(n_25),
.B1(n_29),
.B2(n_32),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_36),
.B1(n_35),
.B2(n_26),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_42),
.Y(n_51)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_0),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_7),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_1),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_21),
.Y(n_61)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_53),
.Y(n_82)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_30),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_15),
.B1(n_23),
.B2(n_19),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_21),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_29),
.B1(n_26),
.B2(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_28),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_28),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_69),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_70),
.B(n_16),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_43),
.Y(n_72)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_4),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_70),
.A2(n_39),
.B(n_44),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_67),
.B(n_57),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_51),
.A2(n_15),
.B1(n_23),
.B2(n_22),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_80),
.A2(n_83),
.B1(n_57),
.B2(n_58),
.Y(n_115)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_92),
.B(n_96),
.C(n_72),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_89),
.B(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_93),
.Y(n_102)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_50),
.A2(n_32),
.B1(n_26),
.B2(n_16),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_32),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_62),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_66),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_13),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_14),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_7),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_77),
.B1(n_93),
.B2(n_87),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_108),
.A2(n_85),
.B1(n_76),
.B2(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_59),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_86),
.B(n_11),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_113),
.B(n_114),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_12),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_49),
.B1(n_59),
.B2(n_85),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_89),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_124),
.C(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_121),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_122),
.B(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_90),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_95),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_83),
.B(n_79),
.C(n_78),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_127),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_81),
.B(n_77),
.C(n_79),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_103),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_49),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_133),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_101),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_127),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_138),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_110),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_110),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_140),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_144),
.B1(n_107),
.B2(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_143),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_135),
.C(n_124),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_149),
.C(n_154),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_SL g147 ( 
.A(n_139),
.B(n_108),
.C(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_147),
.B(n_125),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_151),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_125),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_141),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_112),
.C(n_98),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_144),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_158),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_141),
.B1(n_108),
.B2(n_125),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_160),
.B(n_153),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_153),
.A2(n_108),
.B1(n_65),
.B2(n_58),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_146),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_154),
.B(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_157),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_164),
.B(n_165),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_165),
.C(n_163),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_162),
.A2(n_157),
.B1(n_98),
.B2(n_73),
.Y(n_169)
);

AOI31xp67_ASAP7_75t_SL g173 ( 
.A1(n_169),
.A2(n_4),
.A3(n_6),
.B(n_168),
.Y(n_173)
);

AOI222xp33_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_78),
.B1(n_72),
.B2(n_12),
.C1(n_65),
.C2(n_91),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_169),
.B(n_6),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

AOI31xp33_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_171),
.A3(n_6),
.B(n_170),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_175),
.Y(n_177)
);


endmodule