module fake_jpeg_23708_n_324 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_13),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_32),
.A2(n_23),
.B1(n_13),
.B2(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_13),
.B1(n_14),
.B2(n_36),
.Y(n_66)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_54),
.A2(n_31),
.B1(n_33),
.B2(n_30),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_31),
.A2(n_27),
.B1(n_13),
.B2(n_14),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_56),
.B(n_27),
.C(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_17),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_58),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_42),
.B1(n_61),
.B2(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_61),
.Y(n_82)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_47),
.B1(n_41),
.B2(n_44),
.Y(n_96)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_23),
.B1(n_13),
.B2(n_37),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_72),
.B1(n_76),
.B2(n_78),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_42),
.B1(n_40),
.B2(n_52),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_23),
.B1(n_29),
.B2(n_30),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_43),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_75),
.B(n_44),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_39),
.A2(n_27),
.B1(n_34),
.B2(n_23),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_39),
.A2(n_21),
.B1(n_26),
.B2(n_25),
.Y(n_78)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_84),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_66),
.B1(n_72),
.B2(n_47),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_75),
.B(n_64),
.Y(n_107)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_97),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_53),
.B1(n_74),
.B2(n_62),
.Y(n_119)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_54),
.B1(n_47),
.B2(n_49),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_98),
.A2(n_65),
.B1(n_67),
.B2(n_57),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_57),
.B(n_41),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_91),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_64),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_103),
.A2(n_105),
.B(n_107),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_111),
.B1(n_117),
.B2(n_93),
.Y(n_125)
);

NAND2xp67_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_58),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_68),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_116),
.B1(n_97),
.B2(n_79),
.Y(n_135)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_113),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_85),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_115),
.C(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_100),
.B(n_78),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_60),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_71),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_71),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_71),
.B1(n_62),
.B2(n_49),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_123),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_82),
.B1(n_93),
.B2(n_89),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_87),
.Y(n_138)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_71),
.B1(n_46),
.B2(n_27),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_124),
.A2(n_80),
.B1(n_84),
.B2(n_101),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_141),
.B1(n_104),
.B2(n_109),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_135),
.B1(n_144),
.B2(n_147),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_128),
.B(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_137),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_116),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_82),
.Y(n_134)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_112),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_106),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_140),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_79),
.Y(n_139)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_101),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_148),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_95),
.B1(n_17),
.B2(n_18),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_0),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_0),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_91),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_95),
.B1(n_83),
.B2(n_26),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_108),
.A2(n_26),
.B1(n_21),
.B2(n_20),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_149),
.A2(n_117),
.B1(n_107),
.B2(n_124),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_91),
.Y(n_150)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_151),
.A2(n_22),
.B1(n_19),
.B2(n_25),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_174),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_164),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_109),
.Y(n_157)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_150),
.B1(n_146),
.B2(n_143),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_141),
.B1(n_134),
.B2(n_145),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_115),
.B(n_116),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_160),
.A2(n_178),
.B(n_25),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_118),
.C(n_113),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_137),
.C(n_144),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_165),
.A2(n_18),
.B(n_20),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_135),
.A2(n_122),
.B1(n_123),
.B2(n_26),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_172),
.B1(n_175),
.B2(n_176),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_126),
.B(n_17),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_133),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_77),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_22),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_130),
.A2(n_122),
.B1(n_21),
.B2(n_16),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g174 ( 
.A(n_142),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_130),
.A2(n_122),
.B1(n_21),
.B2(n_16),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_127),
.A2(n_16),
.B1(n_25),
.B2(n_24),
.Y(n_176)
);

AO21x1_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_20),
.B(n_18),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_173),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_179),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_156),
.B(n_136),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_185),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_126),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_183),
.C(n_193),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_149),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_171),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_187),
.B(n_192),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_140),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_198),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_190),
.A2(n_204),
.B1(n_169),
.B2(n_159),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_133),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_145),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_194),
.B(n_202),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_165),
.B(n_24),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_174),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_166),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_94),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_199),
.C(n_154),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_94),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_77),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_178),
.B(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_9),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_212),
.B1(n_225),
.B2(n_191),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_184),
.B(n_153),
.Y(n_207)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_176),
.Y(n_208)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_211),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_167),
.B1(n_166),
.B2(n_162),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_213),
.A2(n_218),
.B(n_222),
.Y(n_229)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_167),
.B(n_151),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_215),
.A2(n_224),
.B1(n_221),
.B2(n_218),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_162),
.B(n_153),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_182),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_175),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_221),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_172),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_224),
.A2(n_7),
.B1(n_11),
.B2(n_10),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_200),
.B(n_152),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_239),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_197),
.B1(n_183),
.B2(n_188),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_228),
.A2(n_232),
.B1(n_238),
.B2(n_241),
.Y(n_257)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_193),
.B1(n_185),
.B2(n_191),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_195),
.B1(n_165),
.B2(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_180),
.C(n_22),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_240),
.C(n_242),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_180),
.B1(n_24),
.B2(n_16),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_19),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_22),
.C(n_19),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_24),
.B1(n_22),
.B2(n_2),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_0),
.C(n_1),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_7),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_246),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_7),
.C(n_11),
.Y(n_244)
);

AOI21x1_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_229),
.B(n_222),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_223),
.B(n_214),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_247),
.A2(n_207),
.B1(n_217),
.B2(n_209),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_228),
.B(n_225),
.Y(n_248)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

OAI321xp33_ASAP7_75t_L g270 ( 
.A1(n_249),
.A2(n_238),
.A3(n_247),
.B1(n_258),
.B2(n_241),
.C(n_265),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_246),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_253),
.B(n_254),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_233),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_216),
.Y(n_256)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_226),
.C(n_206),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_260),
.C(n_264),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_219),
.C(n_217),
.Y(n_260)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_211),
.B(n_8),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_0),
.C(n_1),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_1),
.C(n_2),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_250),
.C(n_252),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_239),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_279),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_231),
.B(n_235),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_269),
.A2(n_270),
.B(n_277),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_251),
.A2(n_242),
.B1(n_2),
.B2(n_3),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_9),
.B1(n_11),
.B2(n_10),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_1),
.Y(n_275)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_2),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_276),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_257),
.B(n_12),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_8),
.Y(n_279)
);

INVx11_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_280),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_8),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_250),
.C(n_255),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_289),
.C(n_292),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_274),
.A2(n_255),
.B1(n_9),
.B2(n_10),
.Y(n_284)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_294),
.C(n_272),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_8),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_287),
.B(n_288),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_271),
.B(n_9),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_276),
.C(n_275),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_10),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_2),
.C(n_3),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_267),
.B(n_278),
.Y(n_295)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

NOR2x1_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_280),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_296),
.B(n_305),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_302),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_268),
.C(n_279),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_301),
.C(n_291),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_273),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_283),
.B(n_6),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_6),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_290),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_307),
.Y(n_316)
);

NAND4xp25_ASAP7_75t_SL g307 ( 
.A(n_296),
.B(n_293),
.C(n_284),
.D(n_292),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_310),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_299),
.B(n_301),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_299),
.B(n_300),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_313),
.B(n_312),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_304),
.B1(n_297),
.B2(n_11),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_12),
.Y(n_318)
);

OAI21x1_ASAP7_75t_SL g319 ( 
.A1(n_317),
.A2(n_318),
.B(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_314),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_311),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_3),
.C(n_5),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);


endmodule