module fake_jpeg_15150_n_249 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_32),
.B(n_35),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_0),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_28),
.B1(n_19),
.B2(n_18),
.Y(n_45)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_45),
.A2(n_46),
.B1(n_52),
.B2(n_53),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_28),
.B1(n_19),
.B2(n_30),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_18),
.B1(n_23),
.B2(n_20),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_58),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_30),
.B1(n_20),
.B2(n_23),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_18),
.B1(n_23),
.B2(n_26),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_25),
.B1(n_29),
.B2(n_27),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_24),
.B1(n_29),
.B2(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_70),
.Y(n_95)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_62),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_69),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_34),
.B1(n_41),
.B2(n_25),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_64),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_24),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_72),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_32),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_21),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_71),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_21),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_35),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_87),
.Y(n_105)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_34),
.B1(n_41),
.B2(n_18),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_39),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_48),
.B(n_17),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_83),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_45),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_21),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_85),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_49),
.B(n_17),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_43),
.B(n_33),
.C(n_54),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_34),
.B1(n_41),
.B2(n_26),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_39),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_39),
.C(n_38),
.Y(n_97)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_43),
.B(n_33),
.Y(n_109)
);

OAI32xp33_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_26),
.A3(n_17),
.B1(n_31),
.B2(n_16),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_93),
.B(n_43),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_89),
.C(n_61),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_98),
.A2(n_109),
.B(n_33),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_1),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_99),
.B(n_1),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_124),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_38),
.C(n_36),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_82),
.B1(n_73),
.B2(n_70),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_129),
.B1(n_102),
.B2(n_93),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_83),
.B1(n_86),
.B2(n_65),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_95),
.B1(n_101),
.B2(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_59),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_130),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_65),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_135),
.B(n_138),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_81),
.B1(n_68),
.B2(n_74),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_81),
.B1(n_72),
.B2(n_90),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_63),
.B1(n_88),
.B2(n_60),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_67),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_91),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_112),
.B1(n_102),
.B2(n_113),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_101),
.B1(n_110),
.B2(n_96),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_36),
.Y(n_163)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_39),
.B(n_67),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_39),
.Y(n_139)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_149),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_120),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_142),
.B(n_144),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_99),
.B1(n_95),
.B2(n_97),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_160),
.B1(n_116),
.B2(n_136),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_129),
.B1(n_118),
.B2(n_125),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_108),
.B(n_109),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_155),
.A2(n_156),
.B(n_159),
.Y(n_174)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_98),
.A3(n_91),
.B1(n_31),
.B2(n_21),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_117),
.C(n_126),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_138),
.B(n_132),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_114),
.B1(n_78),
.B2(n_4),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_51),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_152),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_154),
.Y(n_168)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_183),
.C(n_154),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_128),
.B(n_130),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_170),
.A2(n_160),
.B1(n_151),
.B2(n_143),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_149),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_173),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_115),
.B1(n_76),
.B2(n_121),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_184),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_140),
.B1(n_146),
.B2(n_157),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_31),
.B(n_16),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_76),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_51),
.C(n_115),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_100),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_186),
.B1(n_199),
.B2(n_197),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_195),
.C(n_197),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_144),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_196),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_147),
.C(n_148),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_177),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_148),
.C(n_3),
.Y(n_197)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_201),
.B(n_202),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_164),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_170),
.C(n_173),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_212),
.C(n_2),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_182),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_205),
.B(n_209),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_190),
.A2(n_180),
.B(n_181),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_211),
.B(n_191),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_185),
.A2(n_171),
.B1(n_165),
.B2(n_176),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_210),
.B1(n_2),
.B2(n_3),
.Y(n_220)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_209),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_167),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_174),
.B(n_179),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_172),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_195),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_214),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_191),
.Y(n_214)
);

OAI321xp33_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_211),
.A3(n_207),
.B1(n_204),
.B2(n_206),
.C(n_208),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_175),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_216),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_200),
.A2(n_166),
.B(n_3),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_219),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_223),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_228),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_230),
.A2(n_217),
.B1(n_223),
.B2(n_204),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_222),
.A2(n_221),
.B(n_219),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_14),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_226),
.B(n_216),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_234),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_225),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_236),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_224),
.B(n_14),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_237),
.A2(n_229),
.B(n_227),
.Y(n_239)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_239),
.Y(n_244)
);

O2A1O1Ixp33_ASAP7_75t_R g242 ( 
.A1(n_240),
.A2(n_235),
.B(n_7),
.C(n_8),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_241),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_12),
.C2(n_6),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_238),
.A2(n_6),
.B(n_7),
.Y(n_243)
);

AO21x1_ASAP7_75t_L g246 ( 
.A1(n_243),
.A2(n_12),
.B(n_8),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_246),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_244),
.B(n_9),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_9),
.Y(n_249)
);


endmodule