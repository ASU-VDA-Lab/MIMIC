module fake_jpeg_377_n_574 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_574);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_574;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_SL g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_1),
.B(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_58),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_57),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_27),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_59),
.B(n_61),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_27),
.B(n_14),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_64),
.Y(n_167)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_65),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_71),
.B(n_76),
.Y(n_139)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_81),
.Y(n_164)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_34),
.B(n_16),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_83),
.B(n_91),
.Y(n_163)
);

BUFx4f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g132 ( 
.A(n_89),
.Y(n_132)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_31),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_34),
.B(n_14),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_16),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_16),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_100),
.B(n_105),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_29),
.B(n_11),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_41),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_107),
.B(n_19),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_58),
.B(n_40),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_113),
.B(n_40),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_19),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_115),
.B(n_129),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_124),
.B(n_171),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_63),
.B(n_19),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_81),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_130),
.B(n_136),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_32),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_53),
.A2(n_32),
.B1(n_29),
.B2(n_24),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_142),
.A2(n_146),
.B1(n_161),
.B2(n_30),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_60),
.A2(n_29),
.B1(n_32),
.B2(n_24),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_74),
.B(n_21),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_155),
.B(n_160),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_77),
.B(n_85),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_62),
.A2(n_86),
.B1(n_103),
.B2(n_69),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_67),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_170),
.B(n_101),
.Y(n_222)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_84),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_172),
.B(n_191),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_115),
.A2(n_54),
.B1(n_68),
.B2(n_90),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_173),
.A2(n_192),
.B1(n_207),
.B2(n_209),
.Y(n_247)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_132),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_177),
.B(n_187),
.Y(n_250)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_178),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g237 ( 
.A(n_179),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_180),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_55),
.C(n_95),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_181),
.B(n_186),
.C(n_35),
.Y(n_257)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_183),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_113),
.A2(n_65),
.B1(n_98),
.B2(n_99),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_184),
.B(n_217),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_185),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_SL g186 ( 
.A(n_125),
.B(n_20),
.C(n_39),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_159),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_160),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_188),
.B(n_198),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_126),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_189),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_109),
.A2(n_21),
.B(n_89),
.C(n_39),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_117),
.A2(n_84),
.B1(n_36),
.B2(n_33),
.Y(n_192)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_114),
.B(n_88),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_195),
.B(n_199),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_129),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_196),
.B(n_140),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_197),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_139),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_139),
.B(n_66),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_200),
.A2(n_228),
.B1(n_33),
.B2(n_44),
.Y(n_239)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_201),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_202),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_118),
.B(n_66),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_203),
.B(n_116),
.Y(n_276)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_153),
.Y(n_205)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_108),
.Y(n_206)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_206),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_109),
.A2(n_30),
.B1(n_44),
.B2(n_43),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_120),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_163),
.A2(n_30),
.B1(n_44),
.B2(n_43),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_28),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_210),
.B(n_213),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_122),
.Y(n_211)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_211),
.Y(n_251)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_143),
.Y(n_212)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_212),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_145),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_119),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_215),
.B(n_216),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_110),
.B(n_64),
.Y(n_216)
);

OA22x2_ASAP7_75t_L g217 ( 
.A1(n_138),
.A2(n_106),
.B1(n_152),
.B2(n_166),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_110),
.B(n_64),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_225),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_120),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_220),
.Y(n_282)
);

INVx6_ASAP7_75t_SL g221 ( 
.A(n_162),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_221),
.Y(n_273)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_222),
.Y(n_260)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_121),
.Y(n_223)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_223),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_123),
.Y(n_224)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_224),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_133),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_147),
.B(n_25),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_234),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g227 ( 
.A(n_135),
.Y(n_227)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_227),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_112),
.A2(n_94),
.B1(n_79),
.B2(n_25),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_121),
.Y(n_229)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_229),
.Y(n_272)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_154),
.Y(n_230)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_230),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_154),
.Y(n_231)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_231),
.Y(n_271)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_232),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_150),
.Y(n_233)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_148),
.B(n_11),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_239),
.A2(n_246),
.B1(n_258),
.B2(n_274),
.Y(n_320)
);

NAND3xp33_ASAP7_75t_L g314 ( 
.A(n_243),
.B(n_257),
.C(n_13),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_169),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_244),
.B(n_277),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_200),
.A2(n_210),
.B1(n_172),
.B2(n_193),
.Y(n_246)
);

OR2x2_ASAP7_75t_SL g255 ( 
.A(n_191),
.B(n_87),
.Y(n_255)
);

OR2x2_ASAP7_75t_SL g335 ( 
.A(n_255),
.B(n_22),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_217),
.A2(n_154),
.B1(n_127),
.B2(n_116),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_256),
.A2(n_221),
.B1(n_224),
.B2(n_174),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_226),
.B1(n_214),
.B2(n_190),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_164),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_259),
.B(n_261),
.C(n_206),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_181),
.B(n_167),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_217),
.A2(n_137),
.B1(n_144),
.B2(n_141),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_184),
.A2(n_166),
.B1(n_144),
.B2(n_141),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_275),
.A2(n_33),
.B1(n_28),
.B2(n_47),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_276),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_204),
.B(n_205),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_174),
.Y(n_278)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_186),
.B(n_134),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_127),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_217),
.A2(n_137),
.B1(n_134),
.B2(n_28),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_283),
.A2(n_256),
.B1(n_223),
.B2(n_247),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_290),
.Y(n_343)
);

NOR3xp33_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_203),
.C(n_194),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_292),
.B(n_310),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_250),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_293),
.B(n_307),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_260),
.A2(n_202),
.B1(n_201),
.B2(n_224),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_294),
.A2(n_324),
.B1(n_335),
.B2(n_339),
.Y(n_363)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_238),
.Y(n_295)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_295),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_203),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_296),
.B(n_309),
.Y(n_370)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_240),
.B(n_183),
.C(n_178),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_297),
.B(n_301),
.C(n_327),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_270),
.B(n_212),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_298),
.B(n_302),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_242),
.A2(n_232),
.B1(n_208),
.B2(n_229),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_299),
.A2(n_312),
.B1(n_281),
.B2(n_285),
.Y(n_346)
);

MAJx2_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_176),
.C(n_231),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_185),
.Y(n_302)
);

CKINVDCx10_ASAP7_75t_R g303 ( 
.A(n_273),
.Y(n_303)
);

BUFx5_ASAP7_75t_L g369 ( 
.A(n_303),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_267),
.B(n_231),
.Y(n_304)
);

XNOR2x1_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_315),
.Y(n_341)
);

INVx13_ASAP7_75t_L g305 ( 
.A(n_237),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_306),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_262),
.B(n_179),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_SL g308 ( 
.A1(n_242),
.A2(n_167),
.B(n_175),
.C(n_182),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_308),
.A2(n_278),
.B(n_269),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_261),
.B(n_233),
.Y(n_309)
);

AND2x6_ASAP7_75t_L g310 ( 
.A(n_255),
.B(n_167),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_266),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_311),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_274),
.A2(n_220),
.B1(n_230),
.B2(n_35),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_313),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_314),
.B(n_318),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_265),
.B(n_227),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_316),
.B(n_317),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_254),
.B(n_227),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_251),
.B(n_180),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_257),
.B(n_247),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_319),
.B(n_334),
.Y(n_342)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_245),
.Y(n_322)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_322),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_280),
.Y(n_323)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_323),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_328),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_237),
.B(n_13),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_326),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_252),
.B(n_182),
.C(n_25),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_263),
.B(n_43),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_236),
.Y(n_329)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_329),
.Y(n_368)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_245),
.Y(n_330)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_330),
.Y(n_354)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_286),
.Y(n_331)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_331),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_253),
.B(n_13),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_332),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_283),
.A2(n_127),
.B1(n_116),
.B2(n_36),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_333),
.A2(n_235),
.B1(n_249),
.B2(n_269),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_289),
.B(n_36),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_271),
.B(n_268),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_336),
.B(n_338),
.Y(n_347)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_268),
.Y(n_337)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_337),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_281),
.B(n_35),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_346),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_348),
.A2(n_312),
.B(n_305),
.Y(n_402)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_320),
.A2(n_241),
.B1(n_282),
.B2(n_285),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_360),
.A2(n_367),
.B1(n_376),
.B2(n_378),
.Y(n_389)
);

OAI32xp33_ASAP7_75t_L g364 ( 
.A1(n_319),
.A2(n_272),
.A3(n_249),
.B1(n_280),
.B2(n_287),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_364),
.B(n_308),
.Y(n_387)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_365),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_303),
.A2(n_235),
.B(n_284),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_366),
.A2(n_380),
.B(n_296),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_299),
.A2(n_282),
.B1(n_287),
.B2(n_248),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_311),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_382),
.Y(n_403)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_322),
.Y(n_373)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_309),
.A2(n_248),
.B1(n_284),
.B2(n_272),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_330),
.Y(n_377)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_377),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_309),
.A2(n_47),
.B1(n_38),
.B2(n_4),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_337),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_379),
.B(n_381),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_308),
.A2(n_38),
.B(n_3),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_300),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_327),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_341),
.B(n_315),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_384),
.B(n_386),
.C(n_421),
.Y(n_443)
);

AND2x6_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_310),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_393),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_341),
.B(n_370),
.C(n_383),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_387),
.A2(n_418),
.B1(n_360),
.B2(n_367),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_352),
.Y(n_388)
);

NOR3xp33_ASAP7_75t_L g449 ( 
.A(n_388),
.B(n_400),
.C(n_405),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_390),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_376),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_392),
.B(n_416),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_340),
.B(n_304),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_374),
.Y(n_394)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_394),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_348),
.A2(n_308),
.B(n_321),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_396),
.A2(n_401),
.B(n_402),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_291),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_397),
.B(n_398),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_349),
.B(n_300),
.Y(n_398)
);

INVx13_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_399),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_352),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_342),
.A2(n_335),
.B(n_296),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_347),
.B(n_297),
.Y(n_404)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_404),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_355),
.B(n_328),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_366),
.Y(n_406)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_406),
.Y(n_436)
);

O2A1O1Ixp33_ASAP7_75t_L g408 ( 
.A1(n_343),
.A2(n_333),
.B(n_323),
.C(n_301),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_408),
.B(n_412),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_380),
.B(n_306),
.Y(n_410)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_410),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_363),
.A2(n_38),
.B1(n_3),
.B2(n_4),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_411),
.A2(n_346),
.B1(n_356),
.B2(n_378),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_347),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_364),
.B(n_1),
.Y(n_413)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_413),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_342),
.B(n_4),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_414),
.Y(n_432)
);

NOR2x1_ASAP7_75t_L g416 ( 
.A(n_370),
.B(n_5),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_362),
.B(n_357),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_417),
.B(n_420),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_370),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_419),
.B(n_356),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_344),
.B(n_6),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_383),
.B(n_344),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_426),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_413),
.A2(n_343),
.B1(n_353),
.B2(n_354),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_427),
.A2(n_416),
.B(n_409),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_428),
.A2(n_445),
.B1(n_416),
.B2(n_359),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_398),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_430),
.B(n_435),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_384),
.B(n_368),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_431),
.B(n_444),
.C(n_450),
.Y(n_461)
);

NOR3xp33_ASAP7_75t_SL g435 ( 
.A(n_397),
.B(n_375),
.C(n_377),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_438),
.B(n_439),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_394),
.B(n_353),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_391),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_441),
.B(n_442),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_391),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_365),
.Y(n_444)
);

XNOR2x1_ASAP7_75t_L g445 ( 
.A(n_386),
.B(n_350),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_387),
.A2(n_358),
.B1(n_373),
.B2(n_354),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_448),
.A2(n_395),
.B1(n_410),
.B2(n_419),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_393),
.B(n_350),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_403),
.B(n_351),
.C(n_379),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_451),
.B(n_453),
.C(n_415),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_405),
.B(n_359),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_452),
.B(n_400),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_404),
.B(n_351),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_446),
.A2(n_406),
.B(n_390),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_455),
.A2(n_437),
.B(n_426),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_448),
.A2(n_410),
.B1(n_412),
.B2(n_392),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_457),
.A2(n_464),
.B1(n_467),
.B2(n_468),
.Y(n_492)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_458),
.Y(n_491)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_435),
.Y(n_459)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_459),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_449),
.B(n_388),
.Y(n_460)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_460),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_447),
.B(n_396),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_463),
.Y(n_498)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_423),
.Y(n_465)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_465),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_440),
.A2(n_402),
.B(n_408),
.Y(n_466)
);

OAI21xp33_ASAP7_75t_SL g506 ( 
.A1(n_466),
.A2(n_474),
.B(n_476),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_447),
.A2(n_389),
.B1(n_395),
.B2(n_411),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_454),
.A2(n_389),
.B1(n_408),
.B2(n_414),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_479),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_401),
.C(n_407),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_470),
.B(n_473),
.C(n_433),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_415),
.Y(n_471)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_471),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_437),
.A2(n_424),
.B1(n_454),
.B2(n_434),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_477),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_444),
.C(n_445),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_409),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_423),
.Y(n_475)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_475),
.Y(n_497)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_436),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_427),
.A2(n_385),
.B1(n_414),
.B2(n_407),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_478),
.A2(n_371),
.B1(n_399),
.B2(n_369),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_436),
.B(n_425),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_432),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_459),
.B(n_429),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_483),
.B(n_482),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_431),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_486),
.B(n_488),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_450),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_487),
.B(n_490),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_469),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_489),
.B(n_494),
.Y(n_524)
);

NAND3xp33_ASAP7_75t_L g490 ( 
.A(n_456),
.B(n_422),
.C(n_424),
.Y(n_490)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_493),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_461),
.B(n_446),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_422),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_502),
.C(n_505),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_501),
.A2(n_466),
.B(n_481),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_433),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_503),
.A2(n_467),
.B1(n_468),
.B2(n_463),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_471),
.B(n_371),
.C(n_399),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_488),
.B(n_480),
.C(n_460),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_508),
.B(n_510),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_489),
.B(n_455),
.C(n_477),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_465),
.Y(n_511)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_511),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_475),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_512),
.B(n_515),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_513),
.B(n_506),
.Y(n_528)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_497),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_496),
.A2(n_478),
.B(n_457),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_516),
.B(n_518),
.Y(n_534)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_500),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_517),
.B(n_520),
.Y(n_531)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_484),
.Y(n_520)
);

NOR3xp33_ASAP7_75t_SL g521 ( 
.A(n_495),
.B(n_463),
.C(n_462),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_521),
.A2(n_492),
.B1(n_504),
.B2(n_476),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_491),
.B(n_462),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_522),
.Y(n_537)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_505),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_523),
.B(n_503),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_525),
.B(n_492),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_524),
.B(n_487),
.C(n_486),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_526),
.B(n_529),
.Y(n_552)
);

BUFx24_ASAP7_75t_SL g527 ( 
.A(n_522),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_527),
.B(n_10),
.Y(n_553)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_528),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_524),
.B(n_494),
.C(n_485),
.Y(n_529)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_532),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_509),
.B(n_519),
.C(n_508),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_533),
.B(n_536),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_535),
.A2(n_540),
.B1(n_464),
.B2(n_521),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_519),
.B(n_510),
.C(n_507),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_507),
.B(n_485),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_499),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_542),
.B(n_529),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_534),
.A2(n_513),
.B(n_516),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_544),
.A2(n_551),
.B(n_528),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_530),
.B(n_511),
.C(n_515),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_545),
.B(n_546),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_526),
.B(n_538),
.C(n_535),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_537),
.A2(n_514),
.B1(n_512),
.B2(n_517),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_547),
.B(n_550),
.Y(n_557)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_539),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_551),
.B(n_553),
.Y(n_558)
);

AOI31xp33_ASAP7_75t_L g562 ( 
.A1(n_555),
.A2(n_559),
.A3(n_560),
.B(n_546),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_556),
.A2(n_542),
.B1(n_541),
.B2(n_8),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_549),
.B(n_545),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_548),
.B(n_531),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g561 ( 
.A1(n_557),
.A2(n_552),
.B(n_543),
.Y(n_561)
);

AO21x1_ASAP7_75t_L g565 ( 
.A1(n_561),
.A2(n_564),
.B(n_558),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_562),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_559),
.B(n_539),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_563),
.B(n_554),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_565),
.B(n_567),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_566),
.B(n_6),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_568),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_570),
.A2(n_569),
.B(n_7),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_571),
.A2(n_6),
.B(n_8),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_572),
.Y(n_573)
);

A2O1A1O1Ixp25_ASAP7_75t_L g574 ( 
.A1(n_573),
.A2(n_8),
.B(n_9),
.C(n_566),
.D(n_567),
.Y(n_574)
);


endmodule