module real_jpeg_26192_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_240;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_128;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_0),
.A2(n_66),
.B1(n_67),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_2),
.A2(n_66),
.B1(n_67),
.B2(n_84),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_2),
.A2(n_39),
.B1(n_41),
.B2(n_84),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

INVx8_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_6),
.A2(n_39),
.B1(n_41),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_57),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_6),
.A2(n_50),
.B1(n_51),
.B2(n_57),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_6),
.A2(n_57),
.B1(n_66),
.B2(n_67),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_7),
.A2(n_27),
.B1(n_39),
.B2(n_41),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_7),
.A2(n_27),
.B1(n_50),
.B2(n_51),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_7),
.A2(n_27),
.B1(n_66),
.B2(n_67),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_8),
.A2(n_66),
.B1(n_67),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_8),
.A2(n_50),
.B1(n_51),
.B2(n_72),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_9),
.A2(n_28),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_9),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_9),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_9),
.A2(n_43),
.B1(n_66),
.B2(n_67),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_11),
.A2(n_39),
.B1(n_41),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_11),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_11),
.A2(n_48),
.B1(n_66),
.B2(n_67),
.Y(n_165)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_13),
.B(n_30),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_13),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_13),
.B(n_38),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_13),
.B(n_51),
.C(n_53),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_13),
.A2(n_39),
.B1(n_41),
.B2(n_156),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_13),
.B(n_108),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_13),
.A2(n_50),
.B1(n_51),
.B2(n_156),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_13),
.B(n_66),
.C(n_79),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_13),
.A2(n_69),
.B(n_215),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_14),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_14),
.A2(n_50),
.B1(n_51),
.B2(n_65),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_16),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_16),
.B(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_141),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_139),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_118),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_20),
.B(n_118),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_85),
.C(n_98),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_21),
.A2(n_22),
.B1(n_85),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_61),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_45),
.B2(n_46),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_25),
.B(n_45),
.C(n_61),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_38),
.B2(n_42),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_26),
.Y(n_100)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

AOI32xp33_ASAP7_75t_L g110 ( 
.A1(n_28),
.A2(n_34),
.A3(n_41),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_31),
.B(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_31),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_31),
.A2(n_136),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_37),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_34),
.B1(n_39),
.B2(n_41),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g112 ( 
.A(n_33),
.B(n_39),
.Y(n_112)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_36),
.A2(n_156),
.B(n_157),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_37),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_37),
.B(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_41),
.B1(n_53),
.B2(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_39),
.B(n_181),
.Y(n_180)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_42),
.Y(n_133)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B(n_55),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_47),
.A2(n_49),
.B1(n_59),
.B2(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_49),
.A2(n_55),
.B(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_51),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx5_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_51),
.B(n_222),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_56),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_58),
.A2(n_106),
.B1(n_108),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_59),
.A2(n_105),
.B(n_107),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_59),
.A2(n_107),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_75),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_62),
.B(n_75),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_64),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_70),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_67),
.B1(n_79),
.B2(n_80),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_67),
.B(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_71),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_69),
.A2(n_87),
.B(n_89),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_69),
.A2(n_116),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_69),
.B(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_69),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_70),
.Y(n_242)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_74),
.A2(n_183),
.B(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_76),
.A2(n_202),
.B(n_203),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_76),
.A2(n_203),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_77),
.A2(n_94),
.B1(n_95),
.B2(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_77),
.B(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_77),
.A2(n_95),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_81),
.A2(n_82),
.B(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_81),
.A2(n_152),
.B(n_188),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_81),
.B(n_156),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_85),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_92),
.B1(n_96),
.B2(n_97),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_97),
.Y(n_127)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_95),
.B(n_153),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_98),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_104),
.C(n_109),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_99),
.B(n_104),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_109),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_110),
.B(n_113),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_114),
.A2(n_226),
.B1(n_228),
.B2(n_230),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_138),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_126),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_137),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B(n_135),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_173),
.B(n_260),
.C(n_265),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_167),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_167),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_158),
.C(n_159),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_144),
.A2(n_145),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_154),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_150),
.C(n_154),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_149),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_156),
.B(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_158),
.B(n_159),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_166),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_168),
.B(n_171),
.C(n_172),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_254),
.B(n_259),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_204),
.B(n_253),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_193),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_178),
.B(n_193),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_186),
.C(n_190),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_179),
.B(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_186),
.A2(n_190),
.B1(n_191),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_189),
.Y(n_202)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_198),
.B2(n_199),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_194),
.B(n_200),
.C(n_201),
.Y(n_258)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_247),
.B(n_252),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_223),
.B(n_246),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_217),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_217),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_221),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_233),
.B(n_245),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_231),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_231),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_229),
.B(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_238),
.B(n_244),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_236),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_243),
.Y(n_238)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_251),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_258),
.Y(n_259)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);


endmodule