module fake_ibex_1434_n_499 (n_64, n_3, n_73, n_65, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_21, n_27, n_16, n_78, n_60, n_70, n_7, n_20, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_13, n_61, n_14, n_0, n_12, n_42, n_77, n_44, n_51, n_46, n_49, n_40, n_66, n_17, n_74, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_32, n_53, n_50, n_11, n_68, n_79, n_35, n_31, n_56, n_23, n_54, n_19, n_499);

input n_64;
input n_3;
input n_73;
input n_65;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_70;
input n_7;
input n_20;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_13;
input n_61;
input n_14;
input n_0;
input n_12;
input n_42;
input n_77;
input n_44;
input n_51;
input n_46;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_32;
input n_53;
input n_50;
input n_11;
input n_68;
input n_79;
input n_35;
input n_31;
input n_56;
input n_23;
input n_54;
input n_19;

output n_499;

wire n_151;
wire n_85;
wire n_395;
wire n_84;
wire n_171;
wire n_103;
wire n_389;
wire n_204;
wire n_274;
wire n_387;
wire n_130;
wire n_177;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_124;
wire n_256;
wire n_418;
wire n_193;
wire n_446;
wire n_108;
wire n_350;
wire n_165;
wire n_452;
wire n_86;
wire n_255;
wire n_175;
wire n_398;
wire n_125;
wire n_304;
wire n_191;
wire n_153;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_478;
wire n_239;
wire n_94;
wire n_134;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_357;
wire n_88;
wire n_412;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_90;
wire n_449;
wire n_176;
wire n_216;
wire n_421;
wire n_475;
wire n_166;
wire n_163;
wire n_114;
wire n_236;
wire n_376;
wire n_377;
wire n_189;
wire n_498;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_89;
wire n_170;
wire n_144;
wire n_270;
wire n_346;
wire n_383;
wire n_113;
wire n_117;
wire n_417;
wire n_471;
wire n_265;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_91;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_228;
wire n_147;
wire n_251;
wire n_384;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_426;
wire n_323;
wire n_469;
wire n_143;
wire n_106;
wire n_386;
wire n_224;
wire n_183;
wire n_453;
wire n_333;
wire n_110;
wire n_306;
wire n_400;
wire n_169;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_109;
wire n_127;
wire n_121;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_434;
wire n_296;
wire n_120;
wire n_168;
wire n_155;
wire n_315;
wire n_441;
wire n_122;
wire n_116;
wire n_370;
wire n_431;
wire n_289;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_136;
wire n_261;
wire n_459;
wire n_367;
wire n_221;
wire n_437;
wire n_355;
wire n_474;
wire n_407;
wire n_102;
wire n_490;
wire n_448;
wire n_99;
wire n_466;
wire n_269;
wire n_156;
wire n_126;
wire n_356;
wire n_104;
wire n_420;
wire n_483;
wire n_141;
wire n_487;
wire n_222;
wire n_186;
wire n_349;
wire n_454;
wire n_295;
wire n_331;
wire n_230;
wire n_96;
wire n_185;
wire n_388;
wire n_352;
wire n_290;
wire n_174;
wire n_467;
wire n_427;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_488;
wire n_139;
wire n_429;
wire n_275;
wire n_129;
wire n_98;
wire n_267;
wire n_245;
wire n_229;
wire n_209;
wire n_472;
wire n_347;
wire n_473;
wire n_445;
wire n_335;
wire n_413;
wire n_82;
wire n_263;
wire n_353;
wire n_359;
wire n_299;
wire n_87;
wire n_262;
wire n_439;
wire n_433;
wire n_137;
wire n_338;
wire n_173;
wire n_477;
wire n_363;
wire n_402;
wire n_180;
wire n_369;
wire n_201;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_401;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_480;
wire n_416;
wire n_365;
wire n_100;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_199;
wire n_495;
wire n_410;
wire n_308;
wire n_463;
wire n_411;
wire n_135;
wire n_283;
wire n_366;
wire n_397;
wire n_111;
wire n_322;
wire n_227;
wire n_115;
wire n_248;
wire n_92;
wire n_451;
wire n_101;
wire n_190;
wire n_138;
wire n_409;
wire n_214;
wire n_238;
wire n_332;
wire n_211;
wire n_218;
wire n_314;
wire n_132;
wire n_277;
wire n_337;
wire n_479;
wire n_225;
wire n_360;
wire n_272;
wire n_468;
wire n_223;
wire n_381;
wire n_382;
wire n_95;
wire n_405;
wire n_415;
wire n_288;
wire n_285;
wire n_247;
wire n_320;
wire n_379;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_118;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_217;
wire n_324;
wire n_391;
wire n_390;
wire n_178;
wire n_303;
wire n_362;
wire n_93;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_266;
wire n_294;
wire n_112;
wire n_485;
wire n_284;
wire n_80;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_476;
wire n_461;
wire n_313;
wire n_345;
wire n_408;
wire n_119;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_212;
wire n_311;
wire n_406;
wire n_97;
wire n_197;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_252;
wire n_396;
wire n_83;
wire n_107;
wire n_149;
wire n_489;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_271;
wire n_241;
wire n_292;
wire n_394;
wire n_81;
wire n_364;
wire n_159;
wire n_231;
wire n_298;
wire n_202;
wire n_160;
wire n_184;
wire n_492;
wire n_232;
wire n_380;
wire n_281;
wire n_425;

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_31),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_13),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_9),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_6),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_18),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_51),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_4),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_39),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_59),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx10_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_26),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_77),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_10),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_49),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_14),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_21),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_24),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_12),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_5),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_12),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_42),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_23),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_15),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_28),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_25),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_32),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_37),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_33),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_8),
.Y(n_132)
);

HB1xp67_ASAP7_75t_SL g133 ( 
.A(n_48),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_52),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_3),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_71),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_80),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_135),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_0),
.Y(n_141)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_35),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_0),
.Y(n_148)
);

OAI22x1_ASAP7_75t_R g149 ( 
.A1(n_80),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_101),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_4),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

AND2x4_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_7),
.Y(n_154)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_83),
.B(n_9),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

BUFx8_ASAP7_75t_SL g165 ( 
.A(n_101),
.Y(n_165)
);

AOI22x1_ASAP7_75t_SL g166 ( 
.A1(n_110),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_89),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_120),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_133),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_91),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_93),
.B(n_27),
.Y(n_173)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_85),
.Y(n_174)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_110),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_120),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_94),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_127),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_127),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_109),
.A2(n_40),
.B(n_41),
.Y(n_183)
);

AND2x4_ASAP7_75t_L g184 ( 
.A(n_112),
.B(n_76),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

OA21x2_ASAP7_75t_L g186 ( 
.A1(n_113),
.A2(n_43),
.B(n_45),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_117),
.B(n_132),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_115),
.B(n_47),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_118),
.B(n_53),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_122),
.B(n_56),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_94),
.Y(n_192)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_94),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_125),
.B(n_61),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_128),
.B(n_63),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_129),
.B(n_64),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_95),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_141),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_142),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_134),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_146),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_158),
.B(n_131),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_145),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_185),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_171),
.A2(n_81),
.B1(n_97),
.B2(n_130),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_142),
.Y(n_218)
);

NAND2xp33_ASAP7_75t_L g219 ( 
.A(n_142),
.B(n_194),
.Y(n_219)
);

AO21x2_ASAP7_75t_L g220 ( 
.A1(n_183),
.A2(n_92),
.B(n_126),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_162),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_142),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

BUFx6f_ASAP7_75t_SL g227 ( 
.A(n_184),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_146),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

BUFx6f_ASAP7_75t_SL g233 ( 
.A(n_184),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_143),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_144),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

AND2x6_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_190),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

AND2x6_ASAP7_75t_L g239 ( 
.A(n_190),
.B(n_65),
.Y(n_239)
);

BUFx16f_ASAP7_75t_R g240 ( 
.A(n_149),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_157),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_161),
.Y(n_242)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_175),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

INVxp33_ASAP7_75t_SL g246 ( 
.A(n_138),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_178),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_178),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_189),
.B(n_98),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_160),
.A2(n_121),
.B1(n_111),
.B2(n_107),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_189),
.B(n_106),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_159),
.B(n_168),
.Y(n_252)
);

OR2x6_ASAP7_75t_L g253 ( 
.A(n_172),
.B(n_103),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_180),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_192),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_160),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_192),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_175),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_186),
.Y(n_259)
);

NAND2xp33_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_196),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_179),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_203),
.B(n_225),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_198),
.B(n_174),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_163),
.B1(n_147),
.B2(n_152),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_169),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_235),
.Y(n_266)
);

OR2x6_ASAP7_75t_L g267 ( 
.A(n_199),
.B(n_166),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_205),
.B(n_164),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_214),
.B(n_211),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_203),
.B(n_173),
.Y(n_270)
);

NAND2xp33_ASAP7_75t_L g271 ( 
.A(n_203),
.B(n_195),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_201),
.B(n_164),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_218),
.B(n_176),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_148),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_188),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_210),
.B(n_191),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_224),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_203),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_234),
.Y(n_279)
);

BUFx6f_ASAP7_75t_SL g280 ( 
.A(n_240),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_200),
.B(n_150),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_225),
.B(n_200),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_209),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_182),
.Y(n_286)
);

NOR3xp33_ASAP7_75t_L g287 ( 
.A(n_215),
.B(n_150),
.C(n_197),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_181),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_228),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_228),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_208),
.B(n_175),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_227),
.A2(n_140),
.B1(n_197),
.B2(n_193),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_140),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_208),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_212),
.B(n_197),
.Y(n_296)
);

NAND2xp33_ASAP7_75t_L g297 ( 
.A(n_239),
.B(n_186),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_253),
.B(n_165),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_L g299 ( 
.A(n_239),
.B(n_186),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_223),
.B(n_72),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_253),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_241),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_245),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_219),
.B(n_259),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_259),
.B(n_220),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_278),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_220),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_260),
.A2(n_259),
.B(n_220),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_273),
.B(n_258),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_281),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_264),
.A2(n_233),
.B1(n_242),
.B2(n_243),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_268),
.B(n_243),
.Y(n_314)
);

NOR3xp33_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_257),
.C(n_255),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_282),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_292),
.Y(n_319)
);

BUFx8_ASAP7_75t_L g320 ( 
.A(n_280),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_294),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_254),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_261),
.A2(n_229),
.B(n_204),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_265),
.A2(n_229),
.B(n_204),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_287),
.A2(n_274),
.B1(n_275),
.B2(n_288),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_262),
.A2(n_230),
.B(n_206),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_295),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_270),
.A2(n_231),
.B(n_207),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_298),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_271),
.A2(n_232),
.B(n_213),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_267),
.B(n_226),
.Y(n_331)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_284),
.A2(n_248),
.B(n_213),
.C(n_216),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_263),
.B(n_236),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_291),
.A2(n_238),
.B(n_217),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_263),
.B(n_248),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_272),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_291),
.A2(n_221),
.B(n_222),
.Y(n_337)
);

AO21x1_ASAP7_75t_L g338 ( 
.A1(n_300),
.A2(n_247),
.B(n_202),
.Y(n_338)
);

A2O1A1Ixp33_ASAP7_75t_L g339 ( 
.A1(n_289),
.A2(n_202),
.B(n_244),
.C(n_290),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_277),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_302),
.A2(n_244),
.B1(n_276),
.B2(n_279),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_278),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_305),
.A2(n_285),
.B(n_283),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_312),
.B(n_296),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_340),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_317),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_329),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_304),
.B(n_316),
.Y(n_348)
);

AO31x2_ASAP7_75t_L g349 ( 
.A1(n_339),
.A2(n_341),
.A3(n_332),
.B(n_333),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_314),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_322),
.Y(n_351)
);

AO31x2_ASAP7_75t_L g352 ( 
.A1(n_335),
.A2(n_330),
.A3(n_324),
.B(n_323),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_315),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_320),
.Y(n_354)
);

AOI21x1_ASAP7_75t_L g355 ( 
.A1(n_311),
.A2(n_328),
.B(n_337),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_320),
.Y(n_356)
);

OAI21x1_ASAP7_75t_L g357 ( 
.A1(n_334),
.A2(n_326),
.B(n_310),
.Y(n_357)
);

AOI21xp33_ASAP7_75t_L g358 ( 
.A1(n_307),
.A2(n_310),
.B(n_342),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_336),
.B(n_325),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_340),
.Y(n_360)
);

BUFx5_ASAP7_75t_L g361 ( 
.A(n_321),
.Y(n_361)
);

NAND2x1p5_ASAP7_75t_L g362 ( 
.A(n_312),
.B(n_269),
.Y(n_362)
);

AO31x2_ASAP7_75t_L g363 ( 
.A1(n_306),
.A2(n_309),
.A3(n_338),
.B(n_308),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_304),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_325),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_312),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_325),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_312),
.B(n_318),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_336),
.A2(n_325),
.B1(n_319),
.B2(n_313),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_325),
.Y(n_370)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_312),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_336),
.B(n_325),
.Y(n_372)
);

AO21x2_ASAP7_75t_L g373 ( 
.A1(n_306),
.A2(n_309),
.B(n_305),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_317),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_312),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_312),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_336),
.B(n_325),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_312),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_320),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

BUFx10_ASAP7_75t_L g381 ( 
.A(n_374),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_365),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_369),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_367),
.A2(n_372),
.B1(n_370),
.B2(n_377),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_345),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_351),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_350),
.A2(n_353),
.B(n_343),
.Y(n_387)
);

AO21x2_ASAP7_75t_L g388 ( 
.A1(n_373),
.A2(n_355),
.B(n_357),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_376),
.Y(n_389)
);

BUFx8_ASAP7_75t_L g390 ( 
.A(n_356),
.Y(n_390)
);

INVx8_ASAP7_75t_L g391 ( 
.A(n_379),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_362),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_344),
.B(n_375),
.Y(n_393)
);

NAND2x1p5_ASAP7_75t_L g394 ( 
.A(n_346),
.B(n_371),
.Y(n_394)
);

AO21x2_ASAP7_75t_L g395 ( 
.A1(n_358),
.A2(n_363),
.B(n_349),
.Y(n_395)
);

AO21x2_ASAP7_75t_L g396 ( 
.A1(n_363),
.A2(n_349),
.B(n_348),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_354),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_371),
.Y(n_399)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_363),
.A2(n_364),
.B(n_349),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_366),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_378),
.B(n_368),
.Y(n_402)
);

CKINVDCx11_ASAP7_75t_R g403 ( 
.A(n_361),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_352),
.A2(n_361),
.B(n_325),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_376),
.A2(n_181),
.B1(n_140),
.B2(n_246),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_406),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_380),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_382),
.B(n_384),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_406),
.Y(n_410)
);

BUFx4f_ASAP7_75t_SL g411 ( 
.A(n_390),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_382),
.B(n_383),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_403),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_403),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_388),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_381),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_385),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_387),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_386),
.B(n_389),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_400),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_412),
.B(n_396),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_420),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_412),
.B(n_404),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_409),
.B(n_396),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_414),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_413),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_410),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_407),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_415),
.B(n_395),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_395),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_418),
.Y(n_432)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_407),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_430),
.B(n_419),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_432),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_426),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_432),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_430),
.B(n_421),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_408),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_431),
.B(n_421),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_431),
.B(n_416),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_439),
.B(n_428),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_435),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_435),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_433),
.B(n_411),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_436),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_427),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_437),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_437),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_425),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_436),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_441),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_452),
.B(n_441),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_452),
.B(n_438),
.Y(n_454)
);

AND2x2_ASAP7_75t_SL g455 ( 
.A(n_447),
.B(n_427),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_443),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_443),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_444),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_444),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_433),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_440),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_455),
.A2(n_451),
.B(n_447),
.Y(n_462)
);

OAI322xp33_ASAP7_75t_L g463 ( 
.A1(n_460),
.A2(n_445),
.A3(n_448),
.B1(n_449),
.B2(n_450),
.C1(n_422),
.C2(n_424),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_454),
.B(n_447),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_446),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_457),
.Y(n_466)
);

OAI31xp33_ASAP7_75t_L g467 ( 
.A1(n_460),
.A2(n_414),
.A3(n_436),
.B(n_426),
.Y(n_467)
);

OAI21xp33_ASAP7_75t_L g468 ( 
.A1(n_461),
.A2(n_440),
.B(n_449),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_461),
.B(n_448),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_453),
.B(n_456),
.Y(n_470)
);

OAI21xp33_ASAP7_75t_L g471 ( 
.A1(n_468),
.A2(n_455),
.B(n_453),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_469),
.B(n_458),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_462),
.A2(n_426),
.B1(n_427),
.B2(n_414),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_465),
.B(n_456),
.Y(n_474)
);

NOR3xp33_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_463),
.C(n_405),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_473),
.A2(n_465),
.B1(n_464),
.B2(n_466),
.Y(n_476)
);

AOI222xp33_ASAP7_75t_L g477 ( 
.A1(n_472),
.A2(n_464),
.B1(n_429),
.B2(n_459),
.C1(n_402),
.C2(n_401),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_475),
.B(n_477),
.Y(n_478)
);

AOI211xp5_ASAP7_75t_L g479 ( 
.A1(n_476),
.A2(n_467),
.B(n_398),
.C(n_474),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_478),
.B(n_470),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_479),
.B(n_391),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_480),
.B(n_391),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_481),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_482),
.B(n_398),
.Y(n_484)
);

NOR2x1_ASAP7_75t_L g485 ( 
.A(n_483),
.B(n_391),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_484),
.Y(n_486)
);

NOR2xp67_ASAP7_75t_L g487 ( 
.A(n_485),
.B(n_390),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_486),
.Y(n_488)
);

NOR3xp33_ASAP7_75t_L g489 ( 
.A(n_487),
.B(n_390),
.C(n_399),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_488),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_489),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_488),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_488),
.Y(n_493)
);

AOI221xp5_ASAP7_75t_L g494 ( 
.A1(n_492),
.A2(n_399),
.B1(n_392),
.B2(n_393),
.C(n_394),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_494),
.B(n_490),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_495),
.B(n_493),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_496),
.A2(n_490),
.B(n_491),
.Y(n_497)
);

OR2x6_ASAP7_75t_L g498 ( 
.A(n_497),
.B(n_394),
.Y(n_498)
);

OAI22xp33_ASAP7_75t_L g499 ( 
.A1(n_498),
.A2(n_397),
.B1(n_417),
.B2(n_413),
.Y(n_499)
);


endmodule