module real_jpeg_9789_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_0),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_0),
.A2(n_35),
.B1(n_61),
.B2(n_62),
.Y(n_79)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_2),
.A2(n_56),
.B1(n_65),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_2),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_68),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_68),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_68),
.Y(n_194)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_4),
.A2(n_56),
.B1(n_65),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_4),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_98),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_98),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_98),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_5),
.A2(n_56),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_5),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_5),
.A2(n_61),
.B1(n_62),
.B2(n_66),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_66),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_66),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_6),
.A2(n_61),
.B1(n_62),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_6),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_77),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_77),
.Y(n_124)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_12),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_12),
.A2(n_58),
.B(n_62),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_12),
.A2(n_56),
.B1(n_65),
.B2(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_12),
.B(n_122),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_12),
.A2(n_41),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_12),
.B(n_41),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_12),
.A2(n_30),
.B1(n_106),
.B2(n_173),
.Y(n_175)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_14),
.A2(n_29),
.B1(n_41),
.B2(n_42),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_45),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_45),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_128),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_108),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_20),
.B(n_108),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_88),
.B1(n_89),
.B2(n_107),
.Y(n_20)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_81),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_24),
.B(n_36),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_33),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_25),
.A2(n_30),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_26),
.B(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_27),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_26),
.B(n_39),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_26),
.B(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_27),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_164)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_30),
.A2(n_106),
.B1(n_155),
.B2(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_30),
.A2(n_84),
.B(n_157),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_30),
.A2(n_33),
.B(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_31),
.B(n_34),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_31),
.A2(n_32),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_32),
.B(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_32),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B(n_46),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_38),
.B(n_41),
.C(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_37),
.A2(n_40),
.B1(n_50),
.B2(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_37),
.B(n_48),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_37),
.A2(n_50),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_37),
.B(n_102),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_37),
.A2(n_50),
.B1(n_163),
.B2(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_37),
.A2(n_50),
.B1(n_186),
.B2(n_194),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_37),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_38),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_41),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_42),
.B1(n_72),
.B2(n_73),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_41),
.B(n_72),
.Y(n_201)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_42),
.A2(n_74),
.B1(n_196),
.B2(n_201),
.Y(n_200)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_49),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_50),
.A2(n_194),
.B(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_51),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_69),
.B2(n_70),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_64),
.B2(n_67),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_55),
.A2(n_60),
.B1(n_64),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_55),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B(n_59),
.C(n_60),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_57),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_57),
.B(n_102),
.C(n_103),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_72),
.B(n_74),
.C(n_75),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_72),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g196 ( 
.A(n_62),
.B(n_102),
.CON(n_196),
.SN(n_196)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_76),
.B(n_78),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_71),
.A2(n_75),
.B1(n_141),
.B2(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_80),
.A2(n_92),
.B1(n_93),
.B2(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_80),
.A2(n_92),
.B1(n_117),
.B2(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_80),
.B(n_102),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_83),
.A2(n_105),
.B(n_106),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_85),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.C(n_99),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_91),
.B1(n_95),
.B2(n_96),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B(n_94),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_101),
.B1(n_104),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_102),
.B(n_106),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.C(n_113),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_123),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_116),
.B1(n_123),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_124),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_147),
.B(n_229),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_145),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_130),
.B(n_145),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.C(n_136),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_131),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_134),
.A2(n_136),
.B1(n_137),
.B2(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_134),
.Y(n_227)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.C(n_143),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_138),
.A2(n_139),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_142),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_223),
.B(n_228),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_206),
.B(n_222),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_189),
.B(n_205),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_180),
.B(n_188),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_169),
.B(n_179),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_153),
.B(n_158),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_164),
.B2(n_168),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_159),
.B(n_168),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_162),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_164),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_174),
.B(n_178),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_171),
.B(n_172),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_181),
.B(n_182),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_183),
.B(n_190),
.Y(n_205)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_185),
.CI(n_187),
.CON(n_183),
.SN(n_183)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_199),
.B2(n_204),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_193),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_195),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_198),
.C(n_204),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_199),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_202),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_208),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_214),
.B2(n_215),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_217),
.C(n_220),
.Y(n_224)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_216),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_224),
.B(n_225),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);


endmodule