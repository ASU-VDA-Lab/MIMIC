module real_jpeg_25039_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_0),
.B(n_17),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_0),
.B(n_61),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_0),
.B(n_43),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_0),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_0),
.B(n_40),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_0),
.B(n_50),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_0),
.B(n_208),
.Y(n_349)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_2),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_2),
.B(n_61),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_2),
.B(n_43),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_2),
.B(n_36),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_2),
.B(n_40),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_2),
.B(n_50),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_2),
.B(n_130),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_2),
.B(n_208),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_5),
.B(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_5),
.B(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_5),
.B(n_36),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_5),
.B(n_40),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_5),
.B(n_50),
.Y(n_192)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_5),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_5),
.B(n_228),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_6),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_6),
.B(n_61),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_6),
.B(n_43),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_6),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_6),
.B(n_50),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_6),
.B(n_130),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_6),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_7),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_7),
.B(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_7),
.B(n_61),
.Y(n_79)
);

NAND2x1_ASAP7_75t_SL g94 ( 
.A(n_7),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_7),
.B(n_40),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_7),
.B(n_50),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_7),
.B(n_130),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_7),
.B(n_228),
.Y(n_227)
);

INVx8_ASAP7_75t_SL g132 ( 
.A(n_8),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_9),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_9),
.B(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_9),
.B(n_43),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_9),
.B(n_36),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_9),
.B(n_40),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_9),
.B(n_50),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_9),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_9),
.B(n_166),
.Y(n_301)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_11),
.B(n_160),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_11),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_11),
.B(n_43),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_11),
.B(n_36),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_11),
.B(n_40),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_11),
.B(n_50),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_11),
.B(n_130),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_11),
.B(n_208),
.Y(n_364)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_12),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_13),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_13),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_13),
.B(n_36),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_13),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_13),
.B(n_61),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_13),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_14),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_14),
.B(n_43),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_14),
.B(n_40),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_14),
.B(n_50),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_14),
.B(n_330),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_16),
.B(n_43),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_16),
.B(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_16),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_16),
.B(n_50),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_16),
.B(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_16),
.B(n_208),
.Y(n_207)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_17),
.Y(n_106)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_374),
.B(n_383),
.C(n_387),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_373),
.C(n_382),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_358),
.C(n_359),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_336),
.C(n_337),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_305),
.C(n_306),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_280),
.C(n_281),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_249),
.C(n_250),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_212),
.C(n_213),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_173),
.C(n_174),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_139),
.C(n_140),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_111),
.C(n_112),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_72),
.C(n_83),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_53),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_45),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_33),
.B(n_45),
.C(n_53),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.C(n_41),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_34),
.A2(n_35),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_36),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_40),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_44),
.B(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_46),
.B(n_48),
.C(n_49),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_63),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_54),
.B(n_64),
.C(n_65),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_58),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_61),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_67),
.B(n_71),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_69),
.Y(n_233)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_70),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.C(n_82),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_77),
.B1(n_82),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_107),
.C(n_108),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_92),
.C(n_98),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_90),
.C(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.C(n_102),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_101),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_106),
.B(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_125),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_126),
.C(n_138),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_121),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_120),
.C(n_121),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_116),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_119),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx24_ASAP7_75t_SL g395 ( 
.A(n_121),
.Y(n_395)
);

FAx1_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_123),
.CI(n_124),
.CON(n_121),
.SN(n_121)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_123),
.C(n_124),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_138),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_136),
.B2(n_137),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_129),
.Y(n_135)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_131),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_131),
.B(n_257),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_131),
.B(n_219),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_131),
.B(n_234),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_135),
.C(n_137),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_155),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_144),
.C(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_151),
.C(n_154),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g392 ( 
.A(n_146),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_148),
.CI(n_149),
.CON(n_146),
.SN(n_146)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_147),
.B(n_148),
.C(n_149),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_163),
.C(n_171),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_163),
.B1(n_171),
.B2(n_172),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_158),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_161),
.B(n_162),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_161),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_162),
.B(n_199),
.C(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_169),
.C(n_170),
.Y(n_194)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_167),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_195),
.B2(n_211),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_196),
.C(n_197),
.Y(n_212)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_179),
.C(n_188),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_188),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_180),
.B(n_184),
.C(n_187),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_182),
.B(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_182),
.B(n_234),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_186),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_193),
.C(n_194),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_192),
.Y(n_193)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_202),
.B(n_205),
.C(n_207),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_204),
.B(n_234),
.Y(n_259)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_247),
.B2(n_248),
.Y(n_213)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_238),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_238),
.C(n_247),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_224),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_217),
.B(n_225),
.C(n_226),
.Y(n_268)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_217),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_220),
.CI(n_222),
.CON(n_217),
.SN(n_217)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_218),
.B(n_220),
.C(n_222),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_229),
.B1(n_230),
.B2(n_237),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_227),
.Y(n_237)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_235),
.B2(n_236),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_232),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_236),
.C(n_237),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_231),
.B(n_256),
.C(n_259),
.Y(n_303)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_241),
.C(n_242),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_245),
.C(n_246),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_253),
.C(n_279),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_267),
.B2(n_279),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_261),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_262),
.C(n_263),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_259),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_259),
.A2(n_260),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_SL g320 ( 
.A(n_259),
.B(n_285),
.C(n_288),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g391 ( 
.A(n_263),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_265),
.CI(n_266),
.CON(n_263),
.SN(n_263)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_265),
.C(n_266),
.Y(n_290)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g389 ( 
.A(n_267),
.Y(n_389)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_269),
.CI(n_270),
.CON(n_267),
.SN(n_267)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_269),
.C(n_270),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_278),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_274),
.C(n_276),
.Y(n_298)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_273),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_274),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_275),
.A2(n_276),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_276),
.B(n_302),
.C(n_303),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_304),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_295),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_295),
.C(n_304),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_289),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_284),
.B(n_290),
.C(n_291),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_287),
.A2(n_288),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_SL g347 ( 
.A(n_288),
.B(n_313),
.C(n_315),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g394 ( 
.A(n_291),
.Y(n_394)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.CI(n_294),
.CON(n_291),
.SN(n_291)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_293),
.C(n_294),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_298),
.C(n_299),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_301),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_309),
.C(n_322),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_321),
.B2(n_322),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_317),
.B2(n_318),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_319),
.C(n_320),
.Y(n_339)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_315),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_315),
.A2(n_316),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_352),
.C(n_353),
.Y(n_365)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_325),
.C(n_328),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_328),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_332),
.C(n_335),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_333),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_334),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_338),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_337)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_338),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_340),
.C(n_357),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_346),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_341),
.B(n_347),
.C(n_348),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_362),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_342),
.B(n_360),
.C(n_362),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_344),
.CI(n_345),
.CON(n_342),
.SN(n_342)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_353),
.B2(n_354),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_349),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_350),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_351),
.A2(n_352),
.B1(n_369),
.B2(n_370),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_352),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_369),
.C(n_372),
.Y(n_375)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_355),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_366),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_364),
.B(n_365),
.C(n_366),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_368),
.B1(n_371),
.B2(n_372),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_369),
.A2(n_370),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_370),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_SL g388 ( 
.A(n_370),
.B(n_377),
.C(n_380),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_371),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_374),
.Y(n_373)
);

FAx1_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_376),
.CI(n_381),
.CON(n_374),
.SN(n_374)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_379),
.A2(n_380),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_380),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_384),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_388),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_386),
.Y(n_387)
);


endmodule