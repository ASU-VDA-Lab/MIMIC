module fake_jpeg_29158_n_68 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_68);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_68;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_32),
.B(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_14),
.B1(n_23),
.B2(n_22),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_16),
.B1(n_21),
.B2(n_6),
.Y(n_46)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_39),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_2),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_27),
.C(n_15),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_43),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_27),
.B1(n_13),
.B2(n_5),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_46),
.B1(n_49),
.B2(n_3),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_2),
.B1(n_3),
.B2(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_37),
.CON(n_52),
.SN(n_52)
);

AOI211xp5_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_58),
.B(n_19),
.C(n_20),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_25),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

AO21x1_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_17),
.B(n_18),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_63),
.B(n_64),
.Y(n_65)
);

MAJx2_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_50),
.C(n_55),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_61),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_67),
.B(n_62),
.Y(n_68)
);


endmodule