module real_jpeg_12823_n_23 (n_17, n_8, n_0, n_21, n_2, n_132, n_10, n_9, n_129, n_12, n_135, n_130, n_134, n_6, n_136, n_128, n_133, n_11, n_14, n_131, n_7, n_22, n_18, n_3, n_127, n_5, n_4, n_1, n_20, n_19, n_16, n_15, n_13, n_23);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_132;
input n_10;
input n_9;
input n_129;
input n_12;
input n_135;
input n_130;
input n_134;
input n_6;
input n_136;
input n_128;
input n_133;
input n_11;
input n_14;
input n_131;
input n_7;
input n_22;
input n_18;
input n_3;
input n_127;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_23;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_0),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_1),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_1),
.B(n_88),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_3),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_3),
.B(n_59),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_4),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_4),
.B(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_5),
.B(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_6),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_6),
.B(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_7),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_7),
.B(n_99),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_8),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_10),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_11),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_11),
.B(n_55),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_12),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_12),
.B(n_49),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_13),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_13),
.B(n_82),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_14),
.B(n_36),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_16),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_16),
.B(n_72),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_17),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_19),
.B(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_20),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_21),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_22),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_47),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_27),
.B(n_116),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_27),
.B(n_120),
.Y(n_119)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_28),
.B(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_56),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_30),
.B(n_104),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B(n_125),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_117),
.B(n_121),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_113),
.Y(n_41)
);

NAND3xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_107),
.C(n_112),
.Y(n_42)
);

NAND4xp25_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_48),
.C(n_53),
.D(n_57),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_44),
.A2(n_48),
.B(n_108),
.C(n_111),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_45),
.B(n_46),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_50),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_54),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_102),
.B(n_106),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_98),
.B(n_101),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_86),
.B(n_95),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_81),
.B(n_85),
.Y(n_64)
);

OA21x2_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B(n_80),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B(n_79),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_105),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_115),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_119),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_127),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_128),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_129),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_130),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_131),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_132),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_133),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_134),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_135),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_136),
.Y(n_104)
);


endmodule