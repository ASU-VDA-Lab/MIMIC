module fake_jpeg_4963_n_65 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_65);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_65;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_44;
wire n_28;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_32;

INVx2_ASAP7_75t_SL g21 ( 
.A(n_17),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_1),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_24),
.A2(n_12),
.B1(n_14),
.B2(n_3),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_24),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_26),
.B(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_26),
.A2(n_21),
.B(n_38),
.C(n_30),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_35),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_41),
.B1(n_39),
.B2(n_50),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.Y(n_58)
);

AND2x6_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_46),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_52),
.C(n_53),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_40),
.C(n_51),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_44),
.C(n_43),
.Y(n_61)
);

A2O1A1O1Ixp25_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_62),
.B(n_54),
.C(n_36),
.D(n_49),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_60),
.A2(n_48),
.B1(n_54),
.B2(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

BUFx24_ASAP7_75t_SL g65 ( 
.A(n_64),
.Y(n_65)
);


endmodule