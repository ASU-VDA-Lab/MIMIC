module fake_jpeg_22062_n_20 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_20);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_20;

wire n_13;
wire n_14;
wire n_19;
wire n_18;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_0),
.B(n_9),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_0),
.A2(n_7),
.B1(n_2),
.B2(n_10),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_14),
.B(n_15),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_1),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_3),
.Y(n_16)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_16),
.A2(n_5),
.B(n_6),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_13),
.B(n_8),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_18),
.Y(n_20)
);


endmodule