module fake_jpeg_13120_n_661 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_661);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_661;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_3),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_63),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_8),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_64),
.B(n_127),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_69),
.Y(n_173)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_8),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_71),
.B(n_60),
.Y(n_140)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_72),
.Y(n_193)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_76),
.Y(n_192)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

BUFx24_ASAP7_75t_L g189 ( 
.A(n_77),
.Y(n_189)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_80),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_81),
.Y(n_184)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_83),
.B(n_86),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_84),
.Y(n_196)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_85),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_7),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_87),
.Y(n_212)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_88),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_92),
.Y(n_139)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_91),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_21),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_96),
.Y(n_146)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_98),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_48),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_124),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_100),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_101),
.Y(n_210)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_103),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_27),
.B(n_7),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_104),
.B(n_130),
.Y(n_155)
);

NAND2xp67_ASAP7_75t_L g105 ( 
.A(n_43),
.B(n_11),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_21),
.Y(n_145)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_28),
.Y(n_107)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_110),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_28),
.Y(n_111)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_31),
.Y(n_112)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_31),
.Y(n_113)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_114),
.Y(n_167)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_32),
.Y(n_118)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_118),
.Y(n_188)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_119),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_22),
.Y(n_120)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_25),
.Y(n_121)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_121),
.Y(n_187)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_25),
.Y(n_122)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_122),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_33),
.Y(n_123)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_48),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_40),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_129),
.Y(n_179)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_47),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_47),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_64),
.A2(n_44),
.B(n_27),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_132),
.B(n_135),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_97),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_91),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_137),
.B(n_149),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_140),
.B(n_161),
.Y(n_220)
);

BUFx12_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

BUFx4f_ASAP7_75t_SL g273 ( 
.A(n_144),
.Y(n_273)
);

NAND2xp33_ASAP7_75t_SL g221 ( 
.A(n_145),
.B(n_60),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_86),
.B(n_29),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_74),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_96),
.B(n_29),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_168),
.B(n_183),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_109),
.B(n_44),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_172),
.B(n_178),
.Y(n_269)
);

BUFx12_ASAP7_75t_L g174 ( 
.A(n_77),
.Y(n_174)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_174),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_118),
.B(n_50),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_85),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_182),
.B(n_185),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_72),
.B(n_50),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_110),
.B(n_42),
.Y(n_185)
);

HAxp5_ASAP7_75t_SL g186 ( 
.A(n_94),
.B(n_35),
.CON(n_186),
.SN(n_186)
);

AO22x1_ASAP7_75t_L g274 ( 
.A1(n_186),
.A2(n_213),
.B1(n_1),
.B2(n_2),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_102),
.A2(n_108),
.B1(n_123),
.B2(n_68),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_191),
.A2(n_201),
.B1(n_6),
.B2(n_15),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_127),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_194),
.B(n_198),
.Y(n_282)
);

BUFx12_ASAP7_75t_L g197 ( 
.A(n_106),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_121),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_122),
.B(n_36),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_205),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_69),
.A2(n_33),
.B1(n_46),
.B2(n_25),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_62),
.B(n_36),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_120),
.B(n_42),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_206),
.B(n_214),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_63),
.A2(n_35),
.B1(n_56),
.B2(n_41),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_211),
.A2(n_76),
.B1(n_87),
.B2(n_49),
.Y(n_225)
);

AO22x1_ASAP7_75t_SL g213 ( 
.A1(n_65),
.A2(n_34),
.B1(n_40),
.B2(n_22),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_79),
.B(n_59),
.Y(n_214)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

INVx3_ASAP7_75t_SL g335 ( 
.A(n_218),
.Y(n_335)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_219),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_221),
.B(n_243),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_222),
.Y(n_314)
);

INVx11_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

BUFx24_ASAP7_75t_L g315 ( 
.A(n_223),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_146),
.A2(n_56),
.B1(n_41),
.B2(n_30),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_224),
.A2(n_229),
.B1(n_236),
.B2(n_244),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_225),
.A2(n_230),
.B1(n_232),
.B2(n_156),
.Y(n_317)
);

CKINVDCx12_ASAP7_75t_R g226 ( 
.A(n_189),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_226),
.Y(n_327)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_160),
.Y(n_227)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_227),
.Y(n_297)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_228),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_146),
.A2(n_41),
.B1(n_22),
.B2(n_34),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_145),
.A2(n_67),
.B1(n_113),
.B2(n_112),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_231),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_213),
.A2(n_116),
.B1(n_111),
.B2(n_107),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_148),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_233),
.B(n_261),
.Y(n_296)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_234),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_186),
.A2(n_39),
.B1(n_59),
.B2(n_58),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_237),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_169),
.B(n_47),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_239),
.B(n_252),
.C(n_264),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_155),
.B(n_49),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_240),
.B(n_242),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_L g241 ( 
.A1(n_201),
.A2(n_100),
.B1(n_98),
.B2(n_84),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_241),
.A2(n_151),
.B1(n_152),
.B2(n_143),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_169),
.B(n_58),
.Y(n_242)
);

NAND2xp33_ASAP7_75t_SL g243 ( 
.A(n_179),
.B(n_46),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_163),
.A2(n_52),
.B1(n_39),
.B2(n_46),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_163),
.A2(n_52),
.B1(n_33),
.B2(n_101),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_246),
.A2(n_248),
.B1(n_256),
.B2(n_257),
.Y(n_308)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_164),
.Y(n_247)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_247),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_180),
.A2(n_81),
.B1(n_48),
.B2(n_3),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_249),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_159),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_250),
.Y(n_339)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_164),
.Y(n_251)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_251),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_131),
.B(n_11),
.C(n_16),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_173),
.Y(n_253)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_253),
.Y(n_325)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_142),
.Y(n_254)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_254),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_136),
.B(n_1),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_255),
.B(n_286),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_166),
.A2(n_6),
.B1(n_15),
.B2(n_3),
.Y(n_257)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_189),
.Y(n_258)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_258),
.Y(n_349)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_153),
.Y(n_259)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_259),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_173),
.Y(n_260)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_260),
.Y(n_354)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_165),
.Y(n_261)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_175),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_270),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_139),
.B(n_6),
.C(n_15),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_174),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_266),
.Y(n_305)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_141),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_179),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_267),
.B(n_289),
.Y(n_323)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_147),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_268),
.B(n_280),
.Y(n_318)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_142),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_167),
.B(n_1),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_272),
.Y(n_301)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_176),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_SL g313 ( 
.A1(n_274),
.A2(n_144),
.B(n_2),
.C(n_1),
.Y(n_313)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_202),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_279),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_157),
.A2(n_6),
.B1(n_14),
.B2(n_4),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_278),
.A2(n_158),
.B1(n_195),
.B2(n_210),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_166),
.Y(n_279)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_177),
.Y(n_280)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_177),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_281),
.B(n_283),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_184),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_176),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_284),
.B(n_285),
.Y(n_348)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_188),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_171),
.B(n_150),
.Y(n_286)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_184),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_287),
.B(n_288),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_202),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_156),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_196),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_293),
.B(n_210),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_174),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_294),
.B(n_192),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_263),
.A2(n_211),
.B1(n_200),
.B2(n_157),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_298),
.A2(n_311),
.B1(n_322),
.B2(n_279),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_235),
.B(n_193),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_302),
.B(n_303),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_235),
.B(n_138),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_263),
.A2(n_200),
.B1(n_152),
.B2(n_134),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_271),
.B(n_188),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_312),
.B(n_329),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_313),
.B(n_2),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_317),
.A2(n_331),
.B1(n_340),
.B2(n_258),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_282),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_321),
.B(n_338),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_220),
.B(n_133),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_326),
.B(n_264),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_271),
.B(n_151),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_330),
.Y(n_367)
);

AOI32xp33_ASAP7_75t_L g332 ( 
.A1(n_221),
.A2(n_212),
.A3(n_175),
.B1(n_192),
.B2(n_133),
.Y(n_332)
);

AOI32xp33_ASAP7_75t_L g379 ( 
.A1(n_332),
.A2(n_345),
.A3(n_192),
.B1(n_212),
.B2(n_238),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_240),
.B(n_143),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_334),
.B(n_337),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_286),
.B(n_134),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_277),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_241),
.A2(n_274),
.B1(n_256),
.B2(n_245),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_292),
.B(n_154),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_342),
.B(n_346),
.Y(n_398)
);

MAJx2_ASAP7_75t_L g345 ( 
.A(n_239),
.B(n_190),
.C(n_144),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_242),
.B(n_154),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_223),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_273),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_269),
.B(n_195),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_351),
.B(n_353),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_352),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_239),
.B(n_158),
.Y(n_353)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_295),
.Y(n_356)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_356),
.Y(n_404)
);

NOR2xp67_ASAP7_75t_L g357 ( 
.A(n_303),
.B(n_275),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_357),
.B(n_365),
.Y(n_427)
);

INVx11_ASAP7_75t_L g358 ( 
.A(n_315),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_358),
.Y(n_407)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_348),
.Y(n_359)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_359),
.Y(n_415)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_349),
.Y(n_360)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_360),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_361),
.A2(n_323),
.B1(n_309),
.B2(n_313),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_290),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_363),
.B(n_374),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_318),
.Y(n_365)
);

AND2x6_ASAP7_75t_L g366 ( 
.A(n_326),
.B(n_243),
.Y(n_366)
);

A2O1A1O1Ixp25_ASAP7_75t_L g434 ( 
.A1(n_366),
.A2(n_291),
.B(n_273),
.C(n_314),
.D(n_300),
.Y(n_434)
);

OA21x2_ASAP7_75t_L g432 ( 
.A1(n_368),
.A2(n_300),
.B(n_354),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_339),
.Y(n_370)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_370),
.Y(n_437)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_295),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_371),
.B(n_383),
.Y(n_406)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_299),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_372),
.B(n_380),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_373),
.B(n_310),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_255),
.Y(n_374)
);

INVx13_ASAP7_75t_L g375 ( 
.A(n_315),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_375),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_324),
.B(n_285),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_376),
.B(n_378),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_249),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_379),
.A2(n_391),
.B(n_313),
.Y(n_419)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_299),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_296),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_381),
.B(n_385),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_304),
.B(n_252),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_382),
.B(n_384),
.Y(n_442)
);

AO22x2_ASAP7_75t_L g383 ( 
.A1(n_317),
.A2(n_289),
.B1(n_272),
.B2(n_254),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_346),
.B(n_288),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_309),
.Y(n_385)
);

INVx13_ASAP7_75t_L g386 ( 
.A(n_315),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_386),
.A2(n_393),
.B1(n_399),
.B2(n_401),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_305),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_387),
.B(n_388),
.Y(n_408)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_337),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_390),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_334),
.B(n_276),
.Y(n_390)
);

BUFx5_ASAP7_75t_L g393 ( 
.A(n_327),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_343),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_394),
.B(n_396),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_308),
.A2(n_284),
.B1(n_270),
.B2(n_281),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_395),
.A2(n_335),
.B1(n_344),
.B2(n_353),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_306),
.B(n_247),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_309),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_397),
.B(n_402),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_322),
.A2(n_251),
.B1(n_262),
.B2(n_219),
.Y(n_399)
);

INVx11_ASAP7_75t_L g401 ( 
.A(n_349),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_302),
.B(n_287),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_306),
.B(n_280),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_354),
.Y(n_443)
);

OAI32xp33_ASAP7_75t_L g409 ( 
.A1(n_398),
.A2(n_304),
.A3(n_312),
.B1(n_329),
.B2(n_316),
.Y(n_409)
);

AOI32xp33_ASAP7_75t_L g458 ( 
.A1(n_409),
.A2(n_431),
.A3(n_387),
.B1(n_365),
.B2(n_383),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_389),
.A2(n_331),
.B1(n_336),
.B2(n_316),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_410),
.A2(n_413),
.B1(n_428),
.B2(n_432),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_412),
.B(n_429),
.Y(n_450)
);

FAx1_ASAP7_75t_SL g414 ( 
.A(n_362),
.B(n_310),
.CI(n_345),
.CON(n_414),
.SN(n_414)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_414),
.B(n_382),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_416),
.A2(n_406),
.B1(n_442),
.B2(n_411),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_364),
.B(n_301),
.C(n_297),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_418),
.C(n_422),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_364),
.B(n_301),
.C(n_341),
.Y(n_418)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_419),
.B(n_374),
.C(n_363),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_373),
.B(n_301),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_357),
.B(n_402),
.C(n_362),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_423),
.B(n_378),
.C(n_376),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_400),
.A2(n_313),
.B1(n_335),
.B2(n_320),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_425),
.A2(n_406),
.B1(n_384),
.B2(n_443),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_379),
.A2(n_355),
.B(n_300),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_426),
.A2(n_391),
.B(n_385),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_368),
.A2(n_203),
.B1(n_196),
.B2(n_207),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_398),
.B(n_333),
.Y(n_429)
);

OAI32xp33_ASAP7_75t_L g431 ( 
.A1(n_400),
.A2(n_343),
.A3(n_307),
.B1(n_328),
.B2(n_350),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_434),
.B(n_383),
.Y(n_444)
);

XOR2x1_ASAP7_75t_L g438 ( 
.A(n_392),
.B(n_291),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_438),
.B(n_397),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_392),
.A2(n_403),
.B1(n_396),
.B2(n_395),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_439),
.A2(n_307),
.B1(n_325),
.B2(n_370),
.Y(n_478)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_391),
.A2(n_190),
.B(n_319),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_443),
.Y(n_472)
);

AO21x1_ASAP7_75t_L g505 ( 
.A1(n_444),
.A2(n_447),
.B(n_458),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_442),
.B(n_381),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_445),
.B(n_463),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_427),
.B(n_390),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_446),
.B(n_453),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_449),
.A2(n_469),
.B1(n_477),
.B2(n_432),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_412),
.B(n_359),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_451),
.B(n_470),
.C(n_435),
.Y(n_492)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_430),
.Y(n_452)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_452),
.Y(n_484)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_434),
.B(n_366),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_454),
.A2(n_459),
.B(n_471),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_455),
.A2(n_418),
.B(n_417),
.Y(n_481)
);

INVx13_ASAP7_75t_L g456 ( 
.A(n_420),
.Y(n_456)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_456),
.Y(n_491)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_430),
.Y(n_457)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_457),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_408),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_460),
.B(n_462),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_425),
.B(n_383),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_L g493 ( 
.A1(n_461),
.A2(n_419),
.B(n_436),
.C(n_441),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_408),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_429),
.B(n_369),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_426),
.A2(n_367),
.B(n_377),
.Y(n_464)
);

AO21x1_ASAP7_75t_L g506 ( 
.A1(n_464),
.A2(n_414),
.B(n_413),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_465),
.B(n_438),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_424),
.B(n_371),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_466),
.B(n_467),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_424),
.B(n_393),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_433),
.B(n_356),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_468),
.B(n_474),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_422),
.B(n_372),
.C(n_380),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_410),
.A2(n_383),
.B1(n_360),
.B2(n_358),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_404),
.Y(n_473)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_473),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_423),
.B(n_314),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_411),
.B(n_394),
.Y(n_476)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_476),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_436),
.A2(n_325),
.B1(n_401),
.B2(n_370),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_478),
.A2(n_421),
.B1(n_415),
.B2(n_405),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_435),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_479),
.B(n_480),
.Y(n_515)
);

CKINVDCx14_ASAP7_75t_R g480 ( 
.A(n_440),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_481),
.B(n_500),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_483),
.A2(n_461),
.B1(n_475),
.B2(n_437),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_485),
.A2(n_488),
.B1(n_490),
.B2(n_510),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_486),
.B(n_448),
.C(n_450),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_469),
.A2(n_432),
.B1(n_439),
.B2(n_428),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_SL g490 ( 
.A1(n_472),
.A2(n_420),
.B1(n_415),
.B2(n_421),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_470),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_493),
.B(n_497),
.Y(n_523)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_476),
.Y(n_496)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_496),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_468),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_465),
.Y(n_498)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_498),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_477),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_499),
.B(n_503),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_451),
.B(n_409),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_452),
.Y(n_501)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_501),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_448),
.B(n_414),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_502),
.B(n_455),
.Y(n_522)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_457),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_506),
.Y(n_526)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_473),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_507),
.Y(n_533)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_466),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_509),
.B(n_511),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_449),
.A2(n_441),
.B1(n_407),
.B2(n_431),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_478),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_464),
.Y(n_512)
);

INVx13_ASAP7_75t_L g516 ( 
.A(n_512),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_517),
.B(n_519),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_492),
.B(n_450),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_520),
.B(n_522),
.Y(n_560)
);

NOR2x1_ASAP7_75t_L g524 ( 
.A(n_484),
.B(n_472),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_524),
.B(n_536),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_499),
.A2(n_462),
.B1(n_460),
.B2(n_479),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_525),
.A2(n_532),
.B1(n_537),
.B2(n_547),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_481),
.B(n_458),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_529),
.B(n_539),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_489),
.A2(n_446),
.B(n_445),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_531),
.B(n_504),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_511),
.A2(n_475),
.B1(n_461),
.B2(n_471),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_514),
.B(n_444),
.Y(n_534)
);

CKINVDCx14_ASAP7_75t_R g568 ( 
.A(n_534),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_502),
.B(n_463),
.C(n_459),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_535),
.B(n_538),
.C(n_505),
.Y(n_554)
);

CKINVDCx16_ASAP7_75t_R g536 ( 
.A(n_513),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_486),
.B(n_404),
.C(n_453),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_500),
.B(n_319),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_506),
.B(n_456),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_540),
.B(n_543),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_512),
.A2(n_456),
.B(n_386),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_541),
.B(n_491),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_483),
.A2(n_437),
.B1(n_339),
.B2(n_218),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_542),
.A2(n_491),
.B1(n_487),
.B2(n_503),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_505),
.B(n_273),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_488),
.A2(n_253),
.B1(n_250),
.B2(n_293),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_546),
.B(n_260),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_514),
.A2(n_386),
.B1(n_375),
.B2(n_283),
.Y(n_547)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_548),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_533),
.B(n_482),
.Y(n_549)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_549),
.Y(n_595)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_524),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_550),
.B(n_552),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_526),
.A2(n_489),
.B(n_510),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_551),
.A2(n_553),
.B(n_543),
.Y(n_585)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_544),
.Y(n_552)
);

OAI21xp5_ASAP7_75t_SL g553 ( 
.A1(n_526),
.A2(n_515),
.B(n_485),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_554),
.B(n_529),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_519),
.B(n_530),
.C(n_520),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_556),
.B(n_557),
.C(n_565),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_538),
.B(n_484),
.C(n_487),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_558),
.Y(n_586)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_525),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_559),
.B(n_561),
.Y(n_593)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_523),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_521),
.B(n_501),
.C(n_508),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_521),
.B(n_509),
.C(n_496),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_566),
.B(n_573),
.C(n_522),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_567),
.B(n_533),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_532),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_569),
.A2(n_570),
.B1(n_516),
.B2(n_170),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_518),
.A2(n_495),
.B1(n_507),
.B2(n_494),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_572),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_517),
.B(n_375),
.C(n_238),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_576),
.B(n_588),
.Y(n_596)
);

NOR3xp33_ASAP7_75t_SL g577 ( 
.A(n_550),
.B(n_534),
.C(n_528),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_577),
.B(n_582),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g614 ( 
.A(n_578),
.B(n_587),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_579),
.B(n_583),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_571),
.B(n_540),
.C(n_539),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_549),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_559),
.A2(n_527),
.B1(n_535),
.B2(n_545),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_584),
.A2(n_594),
.B1(n_569),
.B2(n_562),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_585),
.A2(n_548),
.B(n_553),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_563),
.B(n_541),
.Y(n_587)
);

AOI322xp5_ASAP7_75t_L g588 ( 
.A1(n_567),
.A2(n_516),
.A3(n_547),
.B1(n_197),
.B2(n_203),
.C1(n_207),
.C2(n_238),
.Y(n_588)
);

BUFx12_ASAP7_75t_L g589 ( 
.A(n_568),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_589),
.B(n_552),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_590),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_571),
.B(n_556),
.C(n_557),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_591),
.B(n_566),
.C(n_565),
.Y(n_597)
);

XNOR2x1_ASAP7_75t_L g592 ( 
.A(n_564),
.B(n_222),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_SL g604 ( 
.A(n_592),
.B(n_573),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_555),
.A2(n_212),
.B1(n_170),
.B2(n_208),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_597),
.B(n_598),
.Y(n_618)
);

INVx6_ASAP7_75t_L g598 ( 
.A(n_589),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_599),
.B(n_604),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_591),
.B(n_560),
.C(n_554),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_600),
.B(n_601),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_574),
.B(n_560),
.C(n_563),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_602),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_605),
.A2(n_607),
.B(n_611),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_574),
.B(n_562),
.C(n_564),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_606),
.B(n_608),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_593),
.A2(n_551),
.B(n_570),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_578),
.B(n_197),
.C(n_208),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_585),
.A2(n_216),
.B(n_4),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_581),
.B(n_5),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_SL g627 ( 
.A(n_612),
.B(n_5),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_584),
.B(n_2),
.C(n_17),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_613),
.B(n_595),
.C(n_575),
.Y(n_616)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_616),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_603),
.B(n_580),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_619),
.B(n_621),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_606),
.B(n_576),
.C(n_582),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_598),
.B(n_580),
.Y(n_622)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_622),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_610),
.A2(n_586),
.B1(n_575),
.B2(n_595),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_SL g635 ( 
.A1(n_623),
.A2(n_586),
.B1(n_577),
.B2(n_589),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_609),
.B(n_597),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_624),
.B(n_627),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_599),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_628),
.B(n_587),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_613),
.B(n_581),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_629),
.A2(n_605),
.B(n_590),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_620),
.B(n_614),
.C(n_601),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_630),
.A2(n_631),
.B(n_637),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_SL g631 ( 
.A1(n_618),
.A2(n_610),
.B(n_596),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_L g646 ( 
.A(n_632),
.B(n_626),
.C(n_12),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_635),
.B(n_5),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_617),
.B(n_614),
.C(n_600),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_SL g638 ( 
.A1(n_623),
.A2(n_604),
.B1(n_592),
.B2(n_608),
.Y(n_638)
);

AOI322xp5_ASAP7_75t_L g644 ( 
.A1(n_638),
.A2(n_626),
.A3(n_629),
.B1(n_625),
.B2(n_616),
.C1(n_594),
.C2(n_17),
.Y(n_644)
);

CKINVDCx14_ASAP7_75t_R g648 ( 
.A(n_640),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_SL g641 ( 
.A(n_634),
.B(n_615),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_641),
.A2(n_643),
.B(n_639),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_630),
.A2(n_621),
.B(n_625),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_644),
.A2(n_645),
.B1(n_633),
.B2(n_638),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_637),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_646),
.B(n_647),
.Y(n_651)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_649),
.A2(n_650),
.B(n_632),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_642),
.B(n_631),
.Y(n_650)
);

XNOR2xp5_ASAP7_75t_L g652 ( 
.A(n_648),
.B(n_640),
.Y(n_652)
);

XNOR2xp5_ASAP7_75t_SL g656 ( 
.A(n_652),
.B(n_653),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_654),
.B(n_655),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_651),
.A2(n_635),
.B1(n_636),
.B2(n_17),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_657),
.A2(n_656),
.B1(n_636),
.B2(n_14),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_658),
.Y(n_659)
);

BUFx24_ASAP7_75t_SL g660 ( 
.A(n_659),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_660),
.B(n_12),
.Y(n_661)
);


endmodule