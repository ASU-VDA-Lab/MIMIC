module fake_jpeg_2707_n_232 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_232);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_33),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_3),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_11),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_71),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_82),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_69),
.B1(n_57),
.B2(n_76),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_80),
.B1(n_77),
.B2(n_65),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_77),
.B1(n_60),
.B2(n_61),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_60),
.B1(n_81),
.B2(n_78),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_71),
.B1(n_56),
.B2(n_70),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_80),
.B1(n_86),
.B2(n_85),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_94),
.B1(n_93),
.B2(n_63),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_84),
.C(n_56),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_54),
.Y(n_123)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_108),
.Y(n_122)
);

FAx1_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_86),
.CI(n_68),
.CON(n_108),
.SN(n_108)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_73),
.B1(n_58),
.B2(n_55),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_68),
.B1(n_61),
.B2(n_54),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_117),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_115),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_66),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_118),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_74),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_116),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_81),
.B1(n_99),
.B2(n_57),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_99),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_66),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_125),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_9),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_105),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_109),
.A2(n_69),
.B1(n_93),
.B2(n_94),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_135),
.B1(n_4),
.B2(n_5),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_116),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_129),
.B(n_134),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_74),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_8),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_131),
.A2(n_106),
.B1(n_5),
.B2(n_6),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_70),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_2),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_67),
.B1(n_62),
.B2(n_53),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_73),
.B1(n_58),
.B2(n_55),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_139)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_155),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_151),
.B1(n_12),
.B2(n_13),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_141),
.B(n_127),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_141),
.B(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_153),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_137),
.B(n_7),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_152),
.B(n_154),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_52),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_7),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_124),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_157),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_50),
.C(n_49),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_26),
.Y(n_173)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_161),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_163),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_121),
.B(n_9),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_10),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_164),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_166),
.A2(n_175),
.B(n_179),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_141),
.B1(n_131),
.B2(n_13),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_171),
.A2(n_181),
.B1(n_167),
.B2(n_178),
.Y(n_195)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_11),
.B(n_12),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_182),
.B1(n_185),
.B2(n_157),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_32),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_20),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_151),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_145),
.B1(n_142),
.B2(n_153),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_183),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_187),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_166),
.A2(n_156),
.B(n_158),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_171),
.A3(n_168),
.B1(n_165),
.B2(n_180),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_191),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_189),
.A2(n_192),
.B1(n_195),
.B2(n_20),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_184),
.B(n_18),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_177),
.A2(n_172),
.B1(n_165),
.B2(n_175),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_183),
.Y(n_193)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_198),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_36),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_170),
.C(n_181),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_210),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_187),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_40),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_202),
.B(n_206),
.Y(n_211)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_196),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_194),
.B(n_21),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_197),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_38),
.C(n_46),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_201),
.A2(n_190),
.B(n_195),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_212),
.B(n_216),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_200),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_203),
.B(n_188),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_35),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_215),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_205),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_207),
.B(n_224),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_211),
.B(n_213),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_216),
.Y(n_228)
);

AOI321xp33_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_221),
.A3(n_214),
.B1(n_220),
.B2(n_209),
.C(n_210),
.Y(n_229)
);

AOI322xp5_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_34),
.A3(n_45),
.B1(n_44),
.B2(n_29),
.C1(n_48),
.C2(n_43),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_230),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_24),
.Y(n_232)
);


endmodule