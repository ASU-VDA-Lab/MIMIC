module fake_aes_1010_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_SL g10 ( .A(n_0), .Y(n_10) );
HB1xp67_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_7), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_4), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_3), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_2), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_11), .B(n_0), .Y(n_17) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_13), .B(n_1), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_16), .B(n_3), .Y(n_21) );
AOI21xp5_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_14), .B(n_15), .Y(n_22) );
AOI22xp33_ASAP7_75t_L g23 ( .A1(n_19), .A2(n_12), .B1(n_10), .B2(n_6), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_19), .Y(n_24) );
OR2x6_ASAP7_75t_L g25 ( .A(n_21), .B(n_4), .Y(n_25) );
AOI33xp33_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_20), .A3(n_17), .B1(n_18), .B2(n_5), .B3(n_7), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_23), .B1(n_22), .B2(n_18), .Y(n_27) );
AOI21xp5_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_18), .B(n_8), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_27), .B(n_25), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_18), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
NOR2xp33_ASAP7_75t_L g32 ( .A(n_30), .B(n_5), .Y(n_32) );
XNOR2xp5_ASAP7_75t_L g33 ( .A(n_31), .B(n_6), .Y(n_33) );
OAI211xp5_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_18), .B(n_26), .C(n_9), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_31), .Y(n_35) );
NAND3xp33_ASAP7_75t_SL g36 ( .A(n_34), .B(n_35), .C(n_23), .Y(n_36) );
NAND2xp5_ASAP7_75t_L g37 ( .A(n_36), .B(n_33), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_37), .Y(n_38) );
endmodule