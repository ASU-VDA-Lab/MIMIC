module fake_jpeg_29248_n_395 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_395);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_395;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_48),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_61),
.Y(n_99)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_26),
.B(n_36),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_53),
.B(n_79),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_59),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_63),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_72),
.Y(n_145)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_23),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_76),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_31),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_31),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_78),
.Y(n_129)
);

BUFx16f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_29),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_83),
.Y(n_131)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_1),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_25),
.C(n_29),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_40),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_84),
.B(n_85),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_28),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_36),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_28),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_87),
.B(n_93),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_16),
.B1(n_33),
.B2(n_21),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_25),
.B(n_14),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_96),
.B(n_111),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_44),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_132),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_55),
.A2(n_38),
.B1(n_46),
.B2(n_41),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_107),
.A2(n_116),
.B1(n_133),
.B2(n_136),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_109),
.A2(n_47),
.B1(n_78),
.B2(n_68),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_46),
.B1(n_38),
.B2(n_41),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_113),
.A2(n_115),
.B1(n_121),
.B2(n_124),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_69),
.A2(n_46),
.B1(n_38),
.B2(n_16),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_65),
.B1(n_54),
.B2(n_57),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_58),
.A2(n_44),
.B1(n_42),
.B2(n_35),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_117),
.A2(n_118),
.B1(n_127),
.B2(n_137),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_60),
.A2(n_42),
.B1(n_30),
.B2(n_35),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_64),
.A2(n_33),
.B1(n_21),
.B2(n_16),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_33),
.B1(n_21),
.B2(n_30),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_66),
.A2(n_29),
.B1(n_33),
.B2(n_21),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_33),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_50),
.A2(n_21),
.B1(n_29),
.B2(n_4),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_67),
.A2(n_37),
.B1(n_3),
.B2(n_4),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_134),
.A2(n_135),
.B1(n_140),
.B2(n_84),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_71),
.A2(n_37),
.B1(n_4),
.B2(n_5),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_56),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_59),
.A2(n_37),
.B1(n_6),
.B2(n_7),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_70),
.A2(n_37),
.B1(n_7),
.B2(n_8),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_72),
.A2(n_74),
.B1(n_86),
.B2(n_62),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_52),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_142),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_150),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_99),
.B(n_76),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_49),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_156),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_96),
.Y(n_156)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_63),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_166),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_162),
.A2(n_184),
.B1(n_94),
.B2(n_122),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_105),
.B(n_83),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_167),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_179),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_101),
.B(n_100),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_126),
.B(n_132),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_48),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_171),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_170),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_48),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_80),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_172),
.B(n_173),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_81),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_73),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_174),
.B(n_178),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_177),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_90),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_89),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_131),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_182),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_89),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_111),
.B(n_88),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_186),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_138),
.A2(n_78),
.B1(n_47),
.B2(n_91),
.Y(n_184)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_188),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_98),
.B(n_118),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_127),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_106),
.B(n_2),
.Y(n_188)
);

AO21x1_ASAP7_75t_L g238 ( 
.A1(n_200),
.A2(n_204),
.B(n_208),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_117),
.B1(n_146),
.B2(n_125),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_212),
.B1(n_186),
.B2(n_163),
.Y(n_224)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_157),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_206),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_180),
.A2(n_119),
.B1(n_122),
.B2(n_94),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_207),
.A2(n_209),
.B1(n_221),
.B2(n_104),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_116),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_154),
.A2(n_119),
.B1(n_130),
.B2(n_103),
.Y(n_209)
);

BUFx24_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_174),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_181),
.A2(n_107),
.B1(n_146),
.B2(n_103),
.Y(n_212)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_158),
.B(n_95),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_214),
.B(n_158),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_106),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_222),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_153),
.A2(n_130),
.B1(n_144),
.B2(n_123),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_156),
.B(n_104),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_224),
.A2(n_233),
.B1(n_245),
.B2(n_193),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_SL g267 ( 
.A1(n_226),
.A2(n_210),
.B(n_217),
.Y(n_267)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_235),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_173),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_231),
.Y(n_261)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_170),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_212),
.A2(n_181),
.B1(n_176),
.B2(n_160),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_197),
.A2(n_183),
.B(n_172),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_234),
.A2(n_237),
.B(n_249),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_210),
.A2(n_187),
.B1(n_185),
.B2(n_104),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_247),
.B1(n_250),
.B2(n_108),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_189),
.A2(n_165),
.B(n_158),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_192),
.B(n_149),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_239),
.B(n_240),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_192),
.B(n_179),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_202),
.B(n_160),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_242),
.B(n_248),
.Y(n_268)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_244),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_197),
.A2(n_176),
.B1(n_167),
.B2(n_165),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_200),
.A2(n_152),
.B1(n_114),
.B2(n_139),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_191),
.B(n_123),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_189),
.A2(n_187),
.B(n_95),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_200),
.A2(n_139),
.B1(n_144),
.B2(n_159),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_191),
.B(n_112),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_252),
.B(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_205),
.Y(n_253)
);

XNOR2x2_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_214),
.Y(n_254)
);

AOI21xp33_ASAP7_75t_L g295 ( 
.A1(n_254),
.A2(n_248),
.B(n_252),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_262),
.A2(n_267),
.B1(n_274),
.B2(n_245),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_216),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_264),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_202),
.C(n_215),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_231),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_273),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_225),
.A2(n_189),
.B(n_210),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_276),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_240),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_225),
.A2(n_193),
.B1(n_208),
.B2(n_201),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_249),
.A2(n_216),
.B(n_208),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_244),
.B(n_228),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_235),
.A2(n_249),
.B(n_246),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_277),
.A2(n_279),
.B1(n_250),
.B2(n_247),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_237),
.B(n_213),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_220),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_233),
.A2(n_201),
.B1(n_218),
.B2(n_220),
.Y(n_279)
);

AOI21xp33_ASAP7_75t_L g281 ( 
.A1(n_254),
.A2(n_239),
.B(n_213),
.Y(n_281)
);

OAI322xp33_ASAP7_75t_L g312 ( 
.A1(n_281),
.A2(n_284),
.A3(n_295),
.B1(n_286),
.B2(n_293),
.C1(n_288),
.C2(n_280),
.Y(n_312)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_265),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_291),
.Y(n_304)
);

OA21x2_ASAP7_75t_SL g284 ( 
.A1(n_261),
.A2(n_246),
.B(n_237),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_293),
.B1(n_299),
.B2(n_300),
.Y(n_303)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_287),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_297),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_256),
.A2(n_236),
.B(n_226),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_290),
.Y(n_321)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_256),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_292),
.B(n_296),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_262),
.A2(n_224),
.B1(n_238),
.B2(n_218),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_298),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_270),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_257),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_238),
.B1(n_227),
.B2(n_230),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_279),
.A2(n_238),
.B1(n_219),
.B2(n_243),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_269),
.B1(n_275),
.B2(n_276),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_261),
.B(n_219),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_258),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_307),
.A2(n_198),
.B1(n_199),
.B2(n_159),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_278),
.C(n_259),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_313),
.C(n_315),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_263),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_311),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_264),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_SL g326 ( 
.A1(n_312),
.A2(n_295),
.A3(n_284),
.B1(n_300),
.B2(n_290),
.C1(n_298),
.C2(n_291),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_274),
.C(n_268),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_282),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_271),
.C(n_215),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_280),
.A2(n_257),
.B1(n_260),
.B2(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_296),
.A2(n_272),
.B1(n_260),
.B2(n_243),
.Y(n_317)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_317),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_241),
.C(n_232),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_320),
.C(n_299),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_251),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_223),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_253),
.C(n_95),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_302),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_324),
.B(n_325),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_287),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_326),
.A2(n_338),
.B1(n_313),
.B2(n_309),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_333),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_329),
.B(n_330),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_304),
.B(n_294),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_291),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_334),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_314),
.B(n_195),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_223),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_206),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_323),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_336),
.A2(n_206),
.B(n_112),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_315),
.B(n_195),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_217),
.C(n_198),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_306),
.C(n_305),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_340),
.A2(n_323),
.B1(n_320),
.B2(n_318),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_341),
.A2(n_303),
.B1(n_321),
.B2(n_319),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_344),
.A2(n_340),
.B1(n_324),
.B2(n_336),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_346),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_306),
.C(n_311),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_347),
.B(n_355),
.C(n_331),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_325),
.A2(n_199),
.B(n_198),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_348),
.B(n_351),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_349),
.B(n_353),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_337),
.A2(n_169),
.B1(n_164),
.B2(n_151),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_169),
.C(n_164),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_365),
.Y(n_369)
);

MAJx2_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_327),
.C(n_339),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_357),
.A2(n_343),
.B(n_346),
.Y(n_367)
);

OR2x6_ASAP7_75t_L g358 ( 
.A(n_354),
.B(n_333),
.Y(n_358)
);

NOR2x1_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_349),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_361),
.B(n_343),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g362 ( 
.A(n_355),
.B(n_335),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_362),
.A2(n_364),
.B(n_97),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_350),
.A2(n_332),
.B(n_331),
.Y(n_364)
);

O2A1O1Ixp33_ASAP7_75t_L g365 ( 
.A1(n_342),
.A2(n_151),
.B(n_148),
.C(n_120),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_370),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_359),
.B(n_344),
.Y(n_370)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_371),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_352),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_372),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_356),
.B(n_348),
.C(n_351),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_373),
.A2(n_375),
.B(n_376),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_358),
.B(n_353),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_374),
.B(n_363),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_148),
.C(n_139),
.Y(n_375)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_377),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_373),
.B(n_358),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_378),
.A2(n_383),
.B(n_381),
.Y(n_386)
);

AOI322xp5_ASAP7_75t_L g384 ( 
.A1(n_380),
.A2(n_363),
.A3(n_371),
.B1(n_369),
.B2(n_375),
.C1(n_97),
.C2(n_51),
.Y(n_384)
);

AOI322xp5_ASAP7_75t_L g390 ( 
.A1(n_384),
.A2(n_385),
.A3(n_387),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_390)
);

AOI322xp5_ASAP7_75t_L g385 ( 
.A1(n_382),
.A2(n_97),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_2),
.C2(n_11),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_386),
.B(n_378),
.C(n_388),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_9),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_389),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_390),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_386),
.B(n_10),
.C(n_13),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_391),
.C(n_13),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_392),
.C(n_13),
.Y(n_395)
);


endmodule