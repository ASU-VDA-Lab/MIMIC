module fake_netlist_1_12209_n_24 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_24);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_24;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
wire n_7;
INVx2_ASAP7_75t_L g7 ( .A(n_1), .Y(n_7) );
NAND2xp5_ASAP7_75t_SL g8 ( .A(n_1), .B(n_4), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_2), .Y(n_9) );
AOI22xp33_ASAP7_75t_L g10 ( .A1(n_6), .A2(n_3), .B1(n_0), .B2(n_2), .Y(n_10) );
AND2x4_ASAP7_75t_L g11 ( .A(n_5), .B(n_0), .Y(n_11) );
INVx3_ASAP7_75t_L g12 ( .A(n_3), .Y(n_12) );
OAI21x1_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_8), .B(n_7), .Y(n_13) );
AND2x4_ASAP7_75t_L g14 ( .A(n_12), .B(n_9), .Y(n_14) );
NAND2xp5_ASAP7_75t_SL g15 ( .A(n_12), .B(n_11), .Y(n_15) );
O2A1O1Ixp33_ASAP7_75t_L g16 ( .A1(n_9), .A2(n_7), .B(n_11), .C(n_10), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
OR2x2_ASAP7_75t_L g18 ( .A(n_14), .B(n_11), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_18), .B(n_15), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_17), .B(n_16), .Y(n_20) );
OAI22xp33_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_13), .B1(n_16), .B2(n_19), .Y(n_21) );
NOR3xp33_ASAP7_75t_L g22 ( .A(n_21), .B(n_20), .C(n_19), .Y(n_22) );
AOI21xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_20), .B(n_19), .Y(n_23) );
OA21x2_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_19), .B(n_22), .Y(n_24) );
endmodule