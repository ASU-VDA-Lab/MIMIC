module fake_jpeg_25781_n_96 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_45),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_10),
.B1(n_24),
.B2(n_22),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_46),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_57),
.B1(n_3),
.B2(n_4),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_38),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_33),
.B1(n_12),
.B2(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_2),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_3),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_68),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_48),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_9),
.B1(n_21),
.B2(n_19),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_4),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_5),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_5),
.Y(n_71)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_25),
.B1(n_8),
.B2(n_7),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_17),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_6),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_6),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_61),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_89),
.A2(n_64),
.B(n_81),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_90),
.A2(n_91),
.B1(n_83),
.B2(n_66),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_87),
.C(n_62),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_79),
.B(n_81),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_84),
.C(n_72),
.Y(n_94)
);

OAI21x1_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_75),
.B(n_80),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_66),
.B1(n_76),
.B2(n_77),
.Y(n_96)
);


endmodule