module fake_jpeg_10044_n_337 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_37),
.Y(n_48)
);

NAND2x1p5_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_28),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_17),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_60),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_35),
.B1(n_30),
.B2(n_17),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_40),
.B1(n_23),
.B2(n_26),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_35),
.B1(n_30),
.B2(n_17),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_58),
.B1(n_18),
.B2(n_21),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_35),
.B1(n_30),
.B2(n_23),
.Y(n_58)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_35),
.B1(n_30),
.B2(n_23),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_18),
.B1(n_21),
.B2(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_37),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_82),
.Y(n_99)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_40),
.B1(n_38),
.B2(n_41),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_71),
.A2(n_57),
.B1(n_38),
.B2(n_18),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_41),
.B1(n_45),
.B2(n_44),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_73),
.A2(n_60),
.B1(n_59),
.B2(n_54),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_40),
.B1(n_45),
.B2(n_44),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_74),
.A2(n_81),
.B1(n_86),
.B2(n_88),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_45),
.C(n_44),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_85),
.Y(n_103)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_78),
.A2(n_69),
.B1(n_60),
.B2(n_59),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_93),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_23),
.B1(n_20),
.B2(n_33),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_20),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_36),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_29),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_64),
.B1(n_54),
.B2(n_69),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_61),
.A2(n_20),
.B1(n_33),
.B2(n_36),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_98),
.B1(n_49),
.B2(n_57),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_49),
.A2(n_33),
.B1(n_24),
.B2(n_26),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_34),
.B1(n_59),
.B2(n_54),
.Y(n_118)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_95),
.Y(n_122)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_27),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_49),
.A2(n_36),
.B1(n_43),
.B2(n_24),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_97),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_100),
.B(n_101),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_102),
.A2(n_118),
.B1(n_76),
.B2(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_87),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_107),
.B1(n_84),
.B2(n_80),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_43),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_119),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_116),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_110),
.Y(n_156)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_113),
.A2(n_84),
.B(n_80),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_79),
.A2(n_21),
.B1(n_26),
.B2(n_34),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_91),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_46),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_71),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_76),
.B1(n_94),
.B2(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_75),
.C(n_83),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_132),
.C(n_143),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_131),
.A2(n_135),
.B(n_139),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_99),
.C(n_105),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_134),
.A2(n_138),
.B1(n_38),
.B2(n_47),
.Y(n_172)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_136),
.B(n_142),
.Y(n_158)
);

XNOR2x1_ASAP7_75t_SL g139 ( 
.A(n_99),
.B(n_70),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_122),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_83),
.C(n_70),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_144),
.B(n_149),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_71),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_148),
.C(n_119),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_124),
.B1(n_115),
.B2(n_105),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_147),
.A2(n_155),
.B1(n_46),
.B2(n_47),
.Y(n_173)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_71),
.C(n_47),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_153),
.Y(n_174)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_152),
.A2(n_120),
.B1(n_104),
.B2(n_91),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_110),
.B(n_71),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_154),
.B(n_29),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_115),
.A2(n_78),
.B1(n_93),
.B2(n_46),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_100),
.B1(n_107),
.B2(n_113),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_157),
.A2(n_161),
.B1(n_162),
.B2(n_171),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_113),
.B1(n_112),
.B2(n_118),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_109),
.B1(n_117),
.B2(n_114),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_163),
.A2(n_168),
.B1(n_180),
.B2(n_181),
.Y(n_209)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_136),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_127),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_120),
.B1(n_104),
.B2(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_169),
.B(n_179),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_128),
.A2(n_120),
.B1(n_104),
.B2(n_34),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_170),
.A2(n_31),
.B(n_16),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_130),
.A2(n_47),
.B1(n_46),
.B2(n_90),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_31),
.B1(n_27),
.B2(n_16),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_173),
.A2(n_175),
.B1(n_185),
.B2(n_146),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_147),
.A2(n_90),
.B1(n_72),
.B2(n_22),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_72),
.B1(n_22),
.B2(n_32),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_176),
.A2(n_177),
.B1(n_182),
.B2(n_183),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_32),
.B1(n_25),
.B2(n_38),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_144),
.A2(n_32),
.B1(n_25),
.B2(n_2),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_32),
.B1(n_25),
.B2(n_29),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_129),
.B(n_32),
.Y(n_184)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_139),
.A2(n_25),
.B1(n_29),
.B2(n_27),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_131),
.A2(n_29),
.B(n_25),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_186),
.A2(n_189),
.B(n_133),
.Y(n_199)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_142),
.A2(n_31),
.B(n_27),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_169),
.B(n_154),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_191),
.B(n_200),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_132),
.C(n_143),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_196),
.C(n_205),
.Y(n_219)
);

INVx3_ASAP7_75t_SL g194 ( 
.A(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_187),
.A2(n_180),
.B1(n_179),
.B2(n_157),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_201),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g242 ( 
.A1(n_199),
.A2(n_218),
.B(n_167),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_158),
.Y(n_200)
);

A2O1A1O1Ixp25_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_148),
.B(n_135),
.C(n_145),
.D(n_127),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_159),
.B(n_133),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_207),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_203),
.A2(n_168),
.B1(n_161),
.B2(n_162),
.Y(n_223)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_211),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_31),
.C(n_27),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_184),
.B(n_16),
.Y(n_207)
);

OAI22x1_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_182),
.B1(n_218),
.B2(n_194),
.Y(n_234)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_160),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_174),
.A2(n_27),
.B(n_31),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_213),
.A2(n_163),
.B(n_2),
.Y(n_243)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_166),
.B(n_31),
.C(n_1),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_216),
.C(n_189),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_174),
.Y(n_216)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_197),
.A2(n_173),
.B1(n_170),
.B2(n_172),
.Y(n_224)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_237),
.C(n_240),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_178),
.Y(n_226)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_226),
.Y(n_262)
);

XOR2x2_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_186),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_233),
.B(n_245),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_210),
.B1(n_208),
.B2(n_198),
.Y(n_250)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_236),
.Y(n_258)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_175),
.C(n_177),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_238),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_195),
.B(n_188),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_241),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_176),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_213),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_217),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_15),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_207),
.Y(n_259)
);

XOR2x2_ASAP7_75t_SL g245 ( 
.A(n_201),
.B(n_199),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_234),
.A2(n_211),
.B1(n_198),
.B2(n_206),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_246),
.A2(n_233),
.B1(n_238),
.B2(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_232),
.A2(n_195),
.B1(n_206),
.B2(n_217),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_230),
.B1(n_222),
.B2(n_3),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_267),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_226),
.Y(n_255)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_259),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_205),
.C(n_225),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_261),
.C(n_266),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_215),
.C(n_208),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_14),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_265),
.Y(n_270)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_208),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_269),
.A2(n_248),
.B(n_253),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_229),
.Y(n_272)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_251),
.A2(n_227),
.B1(n_243),
.B2(n_237),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_269),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_240),
.C(n_244),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_279),
.C(n_281),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_249),
.A2(n_231),
.B(n_224),
.C(n_223),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_278),
.A2(n_280),
.B1(n_276),
.B2(n_277),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_231),
.C(n_221),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_0),
.C(n_2),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_247),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_256),
.B1(n_246),
.B2(n_260),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_4),
.C(n_5),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_264),
.C(n_259),
.Y(n_290)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_286),
.Y(n_310)
);

AO21x1_ASAP7_75t_L g304 ( 
.A1(n_287),
.A2(n_292),
.B(n_295),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_262),
.B(n_258),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_296),
.Y(n_303)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_290),
.B(n_293),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_260),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_279),
.C(n_274),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_266),
.B1(n_267),
.B2(n_6),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_294),
.A2(n_297),
.B1(n_284),
.B2(n_8),
.Y(n_302)
);

OA22x2_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_267),
.B1(n_5),
.B2(n_7),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_14),
.B(n_13),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_282),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_12),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_299),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_12),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_309),
.C(n_311),
.Y(n_314)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_302),
.A2(n_295),
.B(n_296),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_271),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_294),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_274),
.C(n_271),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_308),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_12),
.Y(n_307)
);

NOR2x1_ASAP7_75t_SL g319 ( 
.A(n_307),
.B(n_13),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_4),
.C(n_8),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_4),
.C(n_8),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_318),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_292),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_319),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_287),
.B(n_295),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_321),
.B1(n_304),
.B2(n_302),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_SL g317 ( 
.A(n_304),
.B(n_295),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_303),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_310),
.A2(n_289),
.B(n_13),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_324),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_300),
.Y(n_324)
);

NOR3xp33_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_327),
.C(n_328),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_301),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_308),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_325),
.A2(n_303),
.B1(n_309),
.B2(n_10),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_325),
.B(n_322),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_329),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_330),
.C(n_9),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_8),
.B(n_9),
.Y(n_335)
);

A2O1A1Ixp33_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_9),
.B(n_11),
.C(n_319),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_9),
.B(n_11),
.Y(n_337)
);


endmodule