module fake_jpeg_26039_n_278 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_22),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_33),
.Y(n_54)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_30),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_19),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_28),
.C(n_17),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_47),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_17),
.B1(n_28),
.B2(n_33),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_42),
.B1(n_41),
.B2(n_40),
.Y(n_73)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_31),
.B(n_28),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_89)
);

NAND2x1_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_36),
.B(n_32),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_61),
.B(n_25),
.Y(n_67)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_64),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_75),
.Y(n_100)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_67),
.B(n_80),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_53),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_41),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_43),
.C(n_53),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_89),
.Y(n_108)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_33),
.B1(n_27),
.B2(n_21),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_76),
.A2(n_79),
.B1(n_90),
.B2(n_36),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_77),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_27),
.B1(n_23),
.B2(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_20),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_83),
.Y(n_110)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_24),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_87),
.B(n_92),
.Y(n_103)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_43),
.A2(n_27),
.B1(n_41),
.B2(n_40),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_88),
.A2(n_36),
.B1(n_40),
.B2(n_45),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_56),
.A2(n_41),
.B1(n_40),
.B2(n_19),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_96),
.B(n_97),
.Y(n_142)
);

OAI211xp5_ASAP7_75t_L g97 ( 
.A1(n_71),
.A2(n_51),
.B(n_46),
.C(n_31),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_35),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_88),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_72),
.B(n_51),
.C(n_34),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_122),
.B(n_69),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_41),
.C(n_45),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_111),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_45),
.C(n_35),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_18),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_113),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_18),
.Y(n_113)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_78),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_93),
.B1(n_94),
.B2(n_91),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_35),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_126),
.A2(n_129),
.B(n_131),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_63),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_127),
.B(n_136),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_78),
.B(n_68),
.Y(n_128)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_114),
.B(n_103),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_62),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_115),
.B1(n_102),
.B2(n_106),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_133),
.Y(n_158)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_68),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_105),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_137),
.Y(n_166)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_116),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_69),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_122),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_64),
.B(n_82),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_102),
.B(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_148),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_82),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_146),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_SL g147 ( 
.A1(n_107),
.A2(n_15),
.A3(n_24),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g177 ( 
.A(n_147),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_113),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_83),
.B1(n_86),
.B2(n_81),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_59),
.B1(n_36),
.B2(n_37),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_66),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_150),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_25),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_75),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_165),
.B1(n_170),
.B2(n_140),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_159),
.A2(n_172),
.B1(n_179),
.B2(n_129),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_167),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_145),
.A2(n_124),
.B1(n_141),
.B2(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_108),
.B(n_122),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_168),
.A2(n_4),
.B(n_6),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_133),
.A2(n_108),
.B1(n_114),
.B2(n_115),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_36),
.B1(n_23),
.B2(n_29),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_35),
.C(n_37),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_123),
.C(n_131),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_129),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_178),
.Y(n_198)
);

AO21x1_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_23),
.B(n_29),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_175),
.B(n_176),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_34),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_35),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_182),
.B(n_184),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_188),
.C(n_199),
.Y(n_211)
);

AOI22x1_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_140),
.B1(n_123),
.B2(n_125),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_189),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_140),
.B1(n_146),
.B2(n_134),
.Y(n_186)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_SL g187 ( 
.A1(n_177),
.A2(n_134),
.A3(n_146),
.B1(n_2),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_187)
);

OA21x2_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_153),
.B(n_175),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_138),
.C(n_35),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_59),
.B1(n_26),
.B2(n_19),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_26),
.B1(n_35),
.B2(n_37),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_161),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_192),
.B(n_194),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_170),
.A2(n_34),
.B1(n_25),
.B2(n_26),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_193),
.Y(n_205)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_26),
.B1(n_35),
.B2(n_2),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_0),
.C(n_1),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_167),
.A2(n_163),
.B1(n_161),
.B2(n_153),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_1),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_203),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_202),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_197),
.B(n_186),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_208),
.B(n_212),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_154),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_156),
.C(n_154),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_215),
.C(n_218),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_156),
.C(n_169),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_171),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_181),
.B(n_157),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_220),
.B(n_221),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_180),
.C(n_166),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_189),
.Y(n_224)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_216),
.A2(n_192),
.B1(n_195),
.B2(n_193),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_226),
.Y(n_238)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_217),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_230),
.Y(n_239)
);

AOI22x1_ASAP7_75t_L g229 ( 
.A1(n_206),
.A2(n_198),
.B1(n_196),
.B2(n_179),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_233),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_213),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_232),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_190),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_162),
.B1(n_199),
.B2(n_9),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_222),
.A2(n_162),
.B1(n_8),
.B2(n_9),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_236),
.B(n_237),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_205),
.A2(n_7),
.B(n_8),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_211),
.C(n_222),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_246),
.Y(n_254)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_223),
.B(n_215),
.CI(n_214),
.CON(n_241),
.SN(n_241)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_218),
.B(n_208),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_225),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_211),
.C(n_212),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_207),
.C(n_219),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_232),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_236),
.A2(n_207),
.B(n_9),
.Y(n_249)
);

OAI21x1_ASAP7_75t_SL g259 ( 
.A1(n_249),
.A2(n_8),
.B(n_10),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_253),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_239),
.B(n_235),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_258),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_234),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_233),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_256),
.C(n_247),
.Y(n_266)
);

AOI31xp33_ASAP7_75t_L g257 ( 
.A1(n_249),
.A2(n_241),
.A3(n_244),
.B(n_245),
.Y(n_257)
);

AOI21xp33_ASAP7_75t_L g261 ( 
.A1(n_257),
.A2(n_250),
.B(n_242),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_248),
.B(n_244),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_259),
.A2(n_231),
.B1(n_243),
.B2(n_13),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_13),
.B(n_10),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_238),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_263),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_265),
.B(n_266),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_263),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_269),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_254),
.C(n_253),
.Y(n_270)
);

FAx1_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_271),
.CI(n_12),
.CON(n_274),
.SN(n_274)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_267),
.A2(n_264),
.B1(n_10),
.B2(n_12),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_268),
.C(n_12),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_274),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_272),
.B(n_274),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_275),
.Y(n_278)
);


endmodule