module fake_jpeg_10810_n_111 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_18),
.Y(n_48)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_46),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_52),
.Y(n_67)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_56),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_48),
.B1(n_41),
.B2(n_44),
.Y(n_55)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_1),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_55),
.B(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_43),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_42),
.B1(n_40),
.B2(n_37),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_65),
.B1(n_36),
.B2(n_4),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_5),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_42),
.B1(n_48),
.B2(n_47),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_59),
.B1(n_67),
.B2(n_60),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_27),
.B1(n_12),
.B2(n_14),
.Y(n_90)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_78),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_2),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_73),
.Y(n_86)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_81),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_21),
.B(n_35),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_80),
.B(n_26),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_47),
.B1(n_36),
.B2(n_5),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_11),
.B1(n_16),
.B2(n_17),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_3),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_3),
.B(n_4),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_7),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_36),
.B(n_6),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_34),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_8),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_92),
.B(n_94),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_74),
.B1(n_80),
.B2(n_32),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_93),
.B1(n_76),
.B2(n_75),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_28),
.C(n_15),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_97),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_29),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_92),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.C(n_90),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_85),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_105),
.A2(n_106),
.B(n_83),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_82),
.C(n_86),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_96),
.B(n_100),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_108),
.Y(n_109)
);

AO221x1_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_102),
.B1(n_94),
.B2(n_33),
.C(n_31),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_30),
.Y(n_111)
);


endmodule