module fake_jpeg_31317_n_540 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_540);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_540;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_18;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

INVx8_ASAP7_75t_SL g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_57),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_59),
.Y(n_163)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g168 ( 
.A(n_65),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_66),
.Y(n_174)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_68),
.Y(n_160)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_69),
.Y(n_156)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_70),
.Y(n_172)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_74),
.Y(n_159)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_80),
.Y(n_176)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_82),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_88),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_22),
.B(n_9),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_92),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_17),
.Y(n_90)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_91),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_22),
.B(n_9),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_93),
.Y(n_166)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_27),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_96),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_39),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_17),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_97),
.Y(n_153)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_98),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_16),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_106),
.Y(n_126)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

BUFx4f_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_109),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_55),
.A2(n_78),
.B1(n_61),
.B2(n_82),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_118),
.A2(n_134),
.B1(n_144),
.B2(n_149),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_24),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_122),
.B(n_123),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_24),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_59),
.B(n_53),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_131),
.B(n_141),
.Y(n_186)
);

BUFx12f_ASAP7_75t_SL g133 ( 
.A(n_65),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_133),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_62),
.A2(n_26),
.B1(n_50),
.B2(n_16),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_60),
.B(n_41),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_87),
.A2(n_53),
.B1(n_46),
.B2(n_41),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_142),
.A2(n_157),
.B1(n_161),
.B2(n_164),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_90),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_63),
.A2(n_50),
.B1(n_16),
.B2(n_28),
.Y(n_149)
);

INVx6_ASAP7_75t_SL g152 ( 
.A(n_65),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_152),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_64),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_68),
.A2(n_50),
.B1(n_28),
.B2(n_48),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_88),
.A2(n_50),
.B1(n_44),
.B2(n_52),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_106),
.B(n_46),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_45),
.Y(n_210)
);

NAND2xp33_ASAP7_75t_SL g177 ( 
.A(n_112),
.B(n_54),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_177),
.B(n_183),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_121),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_178),
.B(n_192),
.Y(n_250)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_179),
.Y(n_244)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_116),
.Y(n_180)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_145),
.A2(n_94),
.B1(n_93),
.B2(n_70),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_181),
.A2(n_197),
.B1(n_206),
.B2(n_209),
.Y(n_260)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_126),
.B(n_66),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_185),
.Y(n_247)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_126),
.B(n_57),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_188),
.B(n_201),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_115),
.B(n_18),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_189),
.B(n_191),
.Y(n_240)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_190),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_115),
.B(n_121),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_171),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_193),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_18),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_194),
.B(n_212),
.Y(n_241)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_124),
.Y(n_195)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_195),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_145),
.A2(n_105),
.B1(n_97),
.B2(n_76),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_196),
.A2(n_217),
.B1(n_226),
.B2(n_158),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_120),
.A2(n_28),
.B1(n_77),
.B2(n_83),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_198),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_125),
.B(n_101),
.C(n_99),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_202),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_171),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_203),
.B(n_207),
.Y(n_251)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_204),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_127),
.Y(n_205)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_205),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_120),
.A2(n_72),
.B1(n_44),
.B2(n_52),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_208),
.B(n_210),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_175),
.A2(n_52),
.B1(n_20),
.B2(n_45),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_150),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_211),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_136),
.B(n_21),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_136),
.B(n_43),
.C(n_21),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_213),
.B(n_27),
.Y(n_236)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_114),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_214),
.B(n_215),
.Y(n_261)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_223),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_137),
.A2(n_102),
.B1(n_75),
.B2(n_27),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_138),
.B(n_47),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_222),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_175),
.A2(n_48),
.B1(n_47),
.B2(n_43),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_220),
.A2(n_168),
.B1(n_143),
.B2(n_153),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_135),
.B(n_38),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_159),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_163),
.B(n_27),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_224),
.B(n_227),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_38),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_225),
.B(n_228),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_146),
.A2(n_169),
.B1(n_162),
.B2(n_155),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_154),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_111),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_132),
.A2(n_20),
.B1(n_27),
.B2(n_10),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_230),
.A2(n_161),
.B1(n_149),
.B2(n_134),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_232),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_189),
.B(n_140),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_234),
.B(n_221),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_198),
.A2(n_172),
.B1(n_151),
.B2(n_147),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_235),
.A2(n_263),
.B1(n_228),
.B2(n_192),
.Y(n_290)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_236),
.A2(n_259),
.B(n_265),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_239),
.A2(n_242),
.B1(n_271),
.B2(n_224),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_166),
.B1(n_147),
.B2(n_160),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_200),
.B(n_194),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_257),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_191),
.B(n_113),
.Y(n_257)
);

OR2x4_ASAP7_75t_L g259 ( 
.A(n_177),
.B(n_188),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_199),
.A2(n_118),
.B1(n_160),
.B2(n_151),
.Y(n_263)
);

OA22x2_ASAP7_75t_L g266 ( 
.A1(n_199),
.A2(n_119),
.B1(n_156),
.B2(n_130),
.Y(n_266)
);

AO22x1_ASAP7_75t_SL g298 ( 
.A1(n_266),
.A2(n_211),
.B1(n_204),
.B2(n_195),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_229),
.A2(n_168),
.B1(n_153),
.B2(n_119),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_222),
.A2(n_143),
.B1(n_27),
.B2(n_10),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_272),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_250),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_274),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_250),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_276),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_240),
.B(n_186),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_281),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_260),
.A2(n_219),
.B(n_212),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_280),
.A2(n_234),
.B(n_227),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_240),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_188),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_282),
.B(n_252),
.Y(n_327)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_261),
.Y(n_283)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_183),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_284),
.B(n_286),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_231),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_285),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_257),
.B(n_183),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_287),
.A2(n_299),
.B1(n_267),
.B2(n_228),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_253),
.B(n_215),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_288),
.B(n_289),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_201),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_290),
.A2(n_294),
.B1(n_298),
.B2(n_239),
.Y(n_307)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_291),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_241),
.B(n_213),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_292),
.B(n_295),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_263),
.A2(n_255),
.B1(n_266),
.B2(n_232),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_245),
.Y(n_296)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_296),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_247),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_297),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_255),
.A2(n_224),
.B1(n_182),
.B2(n_187),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_300),
.Y(n_328)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_254),
.Y(n_301)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_301),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_221),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_302),
.B(n_269),
.Y(n_316)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_243),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_307),
.A2(n_276),
.B1(n_294),
.B2(n_284),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_280),
.A2(n_231),
.B(n_259),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_309),
.A2(n_280),
.B(n_273),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_310),
.A2(n_321),
.B1(n_323),
.B2(n_282),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_311),
.B(n_329),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_316),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_303),
.A2(n_231),
.B1(n_266),
.B2(n_236),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_319),
.A2(n_307),
.B1(n_309),
.B2(n_286),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_303),
.A2(n_266),
.B1(n_241),
.B2(n_267),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_287),
.A2(n_289),
.B1(n_281),
.B2(n_274),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_293),
.A2(n_267),
.B(n_233),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_324),
.A2(n_333),
.B(n_293),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_282),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_295),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_272),
.A2(n_262),
.B1(n_237),
.B2(n_190),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_330),
.Y(n_344)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_296),
.Y(n_334)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_334),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_335),
.B(n_359),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_323),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_358),
.C(n_331),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_329),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_337),
.B(n_363),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_308),
.B(n_278),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_338),
.B(n_346),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_340),
.A2(n_341),
.B1(n_347),
.B2(n_350),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_342),
.A2(n_355),
.B1(n_312),
.B2(n_326),
.Y(n_364)
);

INVx5_ASAP7_75t_SL g343 ( 
.A(n_313),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_343),
.B(n_352),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_345),
.B(n_353),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_278),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_319),
.A2(n_305),
.B1(n_315),
.B2(n_317),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_324),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_238),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_326),
.A2(n_288),
.B1(n_293),
.B2(n_292),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_331),
.B(n_279),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_325),
.B(n_283),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_354),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_310),
.A2(n_290),
.B1(n_277),
.B2(n_291),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_317),
.Y(n_356)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_356),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_237),
.Y(n_357)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_357),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_312),
.B(n_301),
.C(n_300),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_305),
.A2(n_299),
.B(n_298),
.Y(n_359)
);

AOI22x1_ASAP7_75t_L g360 ( 
.A1(n_315),
.A2(n_298),
.B1(n_275),
.B2(n_304),
.Y(n_360)
);

AO22x2_ASAP7_75t_L g377 ( 
.A1(n_360),
.A2(n_332),
.B1(n_328),
.B2(n_320),
.Y(n_377)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_318),
.Y(n_361)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_361),
.Y(n_391)
);

BUFx12f_ASAP7_75t_L g362 ( 
.A(n_314),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_362),
.Y(n_381)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_364),
.A2(n_383),
.B1(n_360),
.B2(n_238),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_365),
.B(n_193),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_344),
.A2(n_321),
.B1(n_306),
.B2(n_333),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_366),
.A2(n_374),
.B1(n_379),
.B2(n_384),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_337),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_372),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_306),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_382),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_337),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_347),
.A2(n_313),
.B1(n_298),
.B2(n_328),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_336),
.B(n_334),
.C(n_332),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_375),
.B(n_256),
.C(n_180),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_377),
.Y(n_415)
);

AO22x1_ASAP7_75t_L g378 ( 
.A1(n_349),
.A2(n_320),
.B1(n_322),
.B2(n_297),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_378),
.A2(n_393),
.B(n_363),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_341),
.A2(n_314),
.B1(n_275),
.B2(n_262),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_248),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_342),
.A2(n_355),
.B1(n_359),
.B2(n_335),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_339),
.A2(n_314),
.B1(n_304),
.B2(n_270),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_344),
.A2(n_270),
.B1(n_243),
.B2(n_207),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_386),
.A2(n_387),
.B1(n_390),
.B2(n_246),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_345),
.A2(n_258),
.B1(n_248),
.B2(n_184),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_356),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_351),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_348),
.A2(n_205),
.B1(n_254),
.B2(n_256),
.Y(n_390)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_392),
.Y(n_394)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_394),
.Y(n_425)
);

NAND3xp33_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_352),
.C(n_338),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_409),
.Y(n_427)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_392),
.Y(n_398)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_398),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_399),
.Y(n_428)
);

A2O1A1Ixp33_ASAP7_75t_SL g400 ( 
.A1(n_378),
.A2(n_360),
.B(n_343),
.C(n_361),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_400),
.A2(n_411),
.B(n_376),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_385),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_406),
.Y(n_434)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_370),
.Y(n_402)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_402),
.Y(n_435)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_391),
.Y(n_403)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_403),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_371),
.B(n_358),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_405),
.B(n_422),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_377),
.B(n_346),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_407),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_377),
.B(n_351),
.Y(n_408)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_408),
.Y(n_426)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_377),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_410),
.A2(n_379),
.B1(n_387),
.B2(n_369),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_376),
.A2(n_362),
.B(n_247),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_393),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_413),
.Y(n_432)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_390),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_374),
.Y(n_414)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_414),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_373),
.B(n_223),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_416),
.A2(n_419),
.B1(n_420),
.B2(n_421),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_417),
.A2(n_404),
.B1(n_413),
.B2(n_414),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_365),
.C(n_383),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_381),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_388),
.B(n_362),
.Y(n_420)
);

INVx13_ASAP7_75t_L g421 ( 
.A(n_381),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_423),
.A2(n_424),
.B(n_445),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_395),
.A2(n_376),
.B(n_366),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_429),
.A2(n_415),
.B1(n_409),
.B2(n_411),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_405),
.B(n_375),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_430),
.B(n_436),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_396),
.B(n_367),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_437),
.B(n_441),
.C(n_444),
.Y(n_447)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_439),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_422),
.B(n_367),
.C(n_382),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_364),
.C(n_369),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_399),
.A2(n_386),
.B(n_362),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_410),
.A2(n_216),
.B1(n_244),
.B2(n_246),
.Y(n_446)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_446),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_SL g449 ( 
.A1(n_425),
.A2(n_398),
.B1(n_394),
.B2(n_412),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_449),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_407),
.Y(n_450)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_450),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_438),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_452),
.B(n_453),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_433),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_208),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_408),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_458),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_423),
.Y(n_457)
);

NOR3xp33_ASAP7_75t_L g483 ( 
.A(n_457),
.B(n_462),
.C(n_179),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_415),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_435),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_460),
.A2(n_463),
.B1(n_426),
.B2(n_442),
.Y(n_473)
);

XNOR2x1_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_396),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_461),
.B(n_464),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_432),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_443),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_428),
.A2(n_400),
.B(n_403),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_437),
.B(n_402),
.C(n_400),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_465),
.B(n_445),
.C(n_428),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_440),
.B(n_400),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_466),
.B(n_464),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_467),
.B(n_473),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_447),
.B(n_430),
.C(n_431),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_469),
.B(n_472),
.Y(n_491)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_471),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_431),
.C(n_441),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_424),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_477),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_439),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_451),
.B(n_442),
.C(n_429),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_479),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_451),
.B(n_426),
.C(n_446),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_452),
.A2(n_421),
.B1(n_244),
.B2(n_246),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_480),
.A2(n_459),
.B1(n_463),
.B2(n_460),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_448),
.B(n_202),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_482),
.B(n_484),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_185),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_477),
.B(n_454),
.C(n_457),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_485),
.B(n_488),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_454),
.C(n_455),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_453),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_489),
.B(n_490),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_466),
.C(n_462),
.Y(n_490)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_493),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_481),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_494),
.B(n_495),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_468),
.A2(n_448),
.B(n_456),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_496),
.A2(n_499),
.B1(n_8),
.B2(n_14),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_450),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_498),
.A2(n_214),
.B1(n_8),
.B2(n_11),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_471),
.A2(n_459),
.B1(n_484),
.B2(n_482),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_496),
.B(n_475),
.Y(n_501)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_501),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_475),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_502),
.B(n_504),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_506),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_6),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_507),
.A2(n_508),
.B(n_509),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_11),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_11),
.C(n_14),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_R g512 ( 
.A(n_498),
.B(n_15),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_512),
.A2(n_514),
.B(n_13),
.Y(n_520)
);

MAJx2_ASAP7_75t_L g513 ( 
.A(n_486),
.B(n_15),
.C(n_13),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_513),
.B(n_511),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_12),
.C(n_13),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_510),
.B(n_490),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_519),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_522),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_507),
.B(n_505),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_501),
.B(n_485),
.Y(n_523)
);

MAJx2_ASAP7_75t_L g525 ( 
.A(n_523),
.B(n_488),
.C(n_500),
.Y(n_525)
);

NOR3xp33_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_511),
.C(n_503),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_524),
.B(n_526),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_525),
.B(n_529),
.C(n_518),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_521),
.A2(n_500),
.B(n_1),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_523),
.A2(n_0),
.B(n_1),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_528),
.A2(n_519),
.B(n_515),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g535 ( 
.A1(n_530),
.A2(n_532),
.B(n_533),
.Y(n_535)
);

OAI21xp33_ASAP7_75t_SL g533 ( 
.A1(n_527),
.A2(n_0),
.B(n_2),
.Y(n_533)
);

OAI311xp33_ASAP7_75t_L g534 ( 
.A1(n_531),
.A2(n_0),
.A3(n_2),
.B1(n_3),
.C1(n_5),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_534),
.B(n_2),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_536),
.B(n_2),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_535),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_538),
.B(n_3),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_3),
.B(n_5),
.Y(n_540)
);


endmodule