module fake_jpeg_1203_n_202 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_202);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_SL g54 ( 
.A(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_0),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_36),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_5),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_46),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_75),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

CKINVDCx6p67_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_80),
.B(n_91),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_54),
.B1(n_50),
.B2(n_47),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_85),
.B1(n_88),
.B2(n_72),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_54),
.B1(n_47),
.B2(n_51),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_56),
.B(n_48),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_61),
.C(n_60),
.Y(n_96)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_62),
.B1(n_64),
.B2(n_51),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_96),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_64),
.B1(n_59),
.B2(n_51),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_101),
.B1(n_104),
.B2(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_99),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_63),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_105),
.Y(n_123)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_49),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_107),
.Y(n_119)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_58),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_67),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_76),
.B1(n_85),
.B2(n_65),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_114),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_59),
.B1(n_87),
.B2(n_53),
.Y(n_114)
);

XOR2x2_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_53),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_44),
.C(n_43),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_35),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_122),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_37),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_128),
.Y(n_147)
);

AO22x1_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_78),
.B1(n_53),
.B2(n_45),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_127),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_33),
.Y(n_128)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_102),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_148),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_95),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_144),
.C(n_149),
.Y(n_159)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_134),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_0),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_1),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_136),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_123),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_30),
.Y(n_160)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_1),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_143),
.Y(n_162)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_95),
.C(n_78),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_2),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_78),
.C(n_42),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_117),
.B1(n_110),
.B2(n_127),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_155),
.B1(n_156),
.B2(n_165),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_128),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_153),
.B(n_160),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_133),
.B(n_130),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_154),
.A2(n_9),
.B(n_10),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_127),
.B1(n_114),
.B2(n_4),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_41),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_12),
.C(n_13),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_169),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_178)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_167),
.Y(n_176)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_39),
.B(n_32),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_172),
.B(n_174),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_152),
.A2(n_31),
.B(n_29),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_175),
.B(n_178),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_21),
.B(n_20),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_179),
.A2(n_163),
.B1(n_160),
.B2(n_162),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_158),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_180),
.B(n_157),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_151),
.C(n_155),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_168),
.B1(n_164),
.B2(n_159),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_182),
.A2(n_185),
.B1(n_170),
.B2(n_174),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_159),
.C(n_173),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_184),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_181),
.Y(n_194)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_191),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_171),
.B(n_177),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_194),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_193),
.A2(n_183),
.B1(n_186),
.B2(n_189),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_195),
.B(n_197),
.Y(n_198)
);

AOI322xp5_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_17),
.A3(n_18),
.B1(n_19),
.B2(n_190),
.C1(n_192),
.C2(n_195),
.Y(n_199)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_17),
.B(n_19),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g201 ( 
.A(n_200),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_198),
.Y(n_202)
);


endmodule