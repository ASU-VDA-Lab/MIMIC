module fake_jpeg_18266_n_88 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_51),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_0),
.CON(n_51),
.SN(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

AO22x1_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_34),
.B1(n_38),
.B2(n_26),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_50),
.B(n_3),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_42),
.B1(n_40),
.B2(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_60),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_44),
.B1(n_37),
.B2(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_1),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_1),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_53),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_71),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_78),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_74),
.B(n_71),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_70),
.C(n_23),
.Y(n_79)
);

AOI322xp5_ASAP7_75t_SL g80 ( 
.A1(n_79),
.A2(n_25),
.A3(n_33),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_11),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_28),
.B(n_32),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_82),
.A2(n_76),
.B1(n_27),
.B2(n_14),
.Y(n_83)
);

AOI322xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_29),
.A3(n_31),
.B1(n_17),
.B2(n_18),
.C1(n_19),
.C2(n_20),
.Y(n_84)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_30),
.CI(n_24),
.CON(n_85),
.SN(n_85)
);

AOI322xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_61),
.A3(n_72),
.B1(n_2),
.B2(n_4),
.C1(n_73),
.C2(n_81),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_85),
.B(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_87),
.B(n_4),
.Y(n_88)
);


endmodule