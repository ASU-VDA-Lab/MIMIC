module fake_jpeg_20216_n_174 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_44),
.Y(n_49)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_24),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_0),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_23),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_62),
.B1(n_63),
.B2(n_33),
.Y(n_78)
);

AO22x1_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_27),
.B1(n_23),
.B2(n_26),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_38),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_29),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_27),
.B(n_22),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_18),
.B1(n_32),
.B2(n_30),
.Y(n_85)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_28),
.B1(n_31),
.B2(n_22),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_34),
.A2(n_29),
.B1(n_28),
.B2(n_32),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_0),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_1),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_70),
.B(n_73),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_85),
.B1(n_47),
.B2(n_69),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_52),
.B(n_20),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_67),
.A3(n_55),
.B1(n_68),
.B2(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_53),
.B1(n_43),
.B2(n_39),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_86),
.B1(n_50),
.B2(n_35),
.Y(n_99)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_41),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_87),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_65),
.A2(n_44),
.B1(n_43),
.B2(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_91),
.Y(n_103)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_90),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_54),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_54),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_48),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_92),
.A2(n_102),
.B1(n_109),
.B2(n_87),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_65),
.B1(n_48),
.B2(n_59),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_99),
.B1(n_79),
.B2(n_89),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_90),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_84),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_39),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_106),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_53),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_80),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_82),
.C(n_85),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_98),
.C(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_120),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_18),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_119),
.Y(n_132)
);

AND2x4_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_116),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_117),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_118),
.A2(n_121),
.B1(n_99),
.B2(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_76),
.B1(n_72),
.B2(n_30),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_76),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_122),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_106),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_15),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_20),
.B1(n_15),
.B2(n_107),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_127),
.B(n_107),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_118),
.Y(n_140)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_109),
.B(n_105),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_116),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_110),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_141),
.B(n_134),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_144),
.A3(n_129),
.B1(n_130),
.B2(n_136),
.C1(n_128),
.C2(n_126),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_120),
.B(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_111),
.B1(n_110),
.B2(n_112),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_145),
.A2(n_148),
.B1(n_138),
.B2(n_133),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_147),
.C(n_134),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_94),
.C(n_93),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_93),
.B1(n_6),
.B2(n_10),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_137),
.C(n_2),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_132),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_151),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_135),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_152),
.A2(n_156),
.B1(n_141),
.B2(n_139),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_142),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_155),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_157),
.B(n_162),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_154),
.A2(n_148),
.B1(n_133),
.B2(n_137),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_155),
.B1(n_153),
.B2(n_151),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_3),
.C(n_4),
.Y(n_166)
);

AOI31xp67_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_1),
.A3(n_2),
.B(n_3),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_165),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_149),
.B(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_162),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_168),
.C(n_158),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_158),
.B(n_161),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_12),
.C(n_13),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_171),
.B(n_3),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_5),
.Y(n_174)
);


endmodule