module fake_aes_10898_n_21 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_21);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_21;
wire n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
CKINVDCx20_ASAP7_75t_R g8 ( .A(n_2), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_5), .Y(n_9) );
BUFx3_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
BUFx2_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
BUFx3_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_13), .B(n_12), .Y(n_14) );
XNOR2xp5_ASAP7_75t_L g15 ( .A(n_14), .B(n_8), .Y(n_15) );
INVx4_ASAP7_75t_R g16 ( .A(n_15), .Y(n_16) );
OR2x2_ASAP7_75t_L g17 ( .A(n_15), .B(n_13), .Y(n_17) );
NAND2xp5_ASAP7_75t_SL g18 ( .A(n_17), .B(n_10), .Y(n_18) );
AOI22xp33_ASAP7_75t_SL g19 ( .A1(n_16), .A2(n_11), .B1(n_0), .B2(n_1), .Y(n_19) );
OAI221xp5_ASAP7_75t_SL g20 ( .A1(n_19), .A2(n_2), .B1(n_3), .B2(n_4), .C(n_6), .Y(n_20) );
OAI22xp5_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_18), .B1(n_3), .B2(n_7), .Y(n_21) );
endmodule