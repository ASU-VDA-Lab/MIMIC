module fake_jpeg_4764_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_21),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_17),
.B1(n_29),
.B2(n_28),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_54),
.B1(n_62),
.B2(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_47),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_18),
.B1(n_25),
.B2(n_20),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_18),
.B1(n_25),
.B2(n_20),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_60),
.Y(n_67)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

CKINVDCx6p67_ASAP7_75t_R g58 ( 
.A(n_31),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_23),
.B(n_29),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_18),
.B1(n_25),
.B2(n_27),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_64),
.B(n_50),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_30),
.B1(n_26),
.B2(n_22),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_62),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_48),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_81),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_30),
.B1(n_26),
.B2(n_22),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_26),
.B1(n_41),
.B2(n_16),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_53),
.B(n_39),
.C(n_46),
.Y(n_88)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_57),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_42),
.A2(n_37),
.B1(n_36),
.B2(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_72),
.B1(n_65),
.B2(n_45),
.Y(n_103)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_94),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_91),
.B1(n_73),
.B2(n_51),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_43),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_58),
.B(n_46),
.C(n_16),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_59),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_58),
.C(n_59),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_77),
.C(n_66),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_16),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_100),
.A2(n_102),
.B(n_70),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_16),
.B(n_23),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_104),
.B1(n_110),
.B2(n_118),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_119),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_113),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_82),
.B1(n_97),
.B2(n_88),
.Y(n_110)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_70),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_86),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_77),
.C(n_66),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_65),
.B(n_2),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_115),
.A2(n_96),
.B1(n_85),
.B2(n_88),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_123),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_61),
.B1(n_73),
.B2(n_51),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_87),
.C(n_100),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_51),
.B1(n_23),
.B2(n_29),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_102),
.B1(n_84),
.B2(n_101),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_71),
.C(n_16),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_109),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_83),
.A2(n_0),
.B(n_29),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_121),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_125),
.B(n_126),
.Y(n_162)
);

INVxp67_ASAP7_75t_SL g126 ( 
.A(n_112),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_111),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_135),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_R g133 ( 
.A(n_117),
.B(n_93),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_136),
.B(n_0),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_92),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_R g136 ( 
.A(n_117),
.B(n_90),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_104),
.C(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_90),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_139),
.Y(n_148)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_105),
.Y(n_140)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_141),
.A2(n_122),
.B1(n_113),
.B2(n_119),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_103),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_142),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_108),
.B(n_101),
.Y(n_143)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_108),
.B(n_143),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_160),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_134),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_110),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_151),
.C(n_132),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_SL g154 ( 
.A1(n_133),
.A2(n_114),
.A3(n_104),
.B1(n_107),
.B2(n_123),
.C1(n_95),
.C2(n_106),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g176 ( 
.A(n_154),
.Y(n_176)
);

AOI32xp33_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_107),
.A3(n_95),
.B1(n_71),
.B2(n_28),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_137),
.B(n_124),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_141),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_142),
.B1(n_131),
.B2(n_125),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_161),
.B1(n_132),
.B2(n_128),
.Y(n_175)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_28),
.B1(n_23),
.B2(n_19),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_165),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_127),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_172),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_159),
.B(n_160),
.Y(n_166)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_178),
.C(n_19),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_171),
.A2(n_146),
.B(n_157),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_134),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_129),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_174),
.Y(n_185)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_175),
.A2(n_157),
.B1(n_146),
.B2(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_0),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_186),
.Y(n_196)
);

OA21x2_ASAP7_75t_SL g182 ( 
.A1(n_165),
.A2(n_155),
.B(n_148),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_183),
.B(n_189),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_169),
.A2(n_153),
.B1(n_152),
.B2(n_159),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_161),
.B1(n_130),
.B2(n_19),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_163),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_19),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_190),
.C(n_178),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_195),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_164),
.C(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_17),
.C(n_3),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_198),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_2),
.C(n_4),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_4),
.B(n_5),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_200),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_184),
.A2(n_4),
.B(n_5),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_5),
.Y(n_201)
);

NOR2xp67_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_189),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_6),
.Y(n_202)
);

AOI21x1_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_191),
.B(n_9),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_193),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_204),
.A2(n_207),
.B(n_208),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_196),
.A2(n_181),
.B1(n_184),
.B2(n_179),
.Y(n_208)
);

OAI221xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_185),
.B1(n_202),
.B2(n_10),
.C(n_11),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_196),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_214),
.C(n_6),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_206),
.B(n_191),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_213),
.B(n_216),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_194),
.C(n_185),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_204),
.A2(n_208),
.B(n_186),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_215),
.A2(n_203),
.B(n_9),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_218),
.A2(n_219),
.B(n_220),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_203),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_217),
.A2(n_6),
.B(n_10),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_12),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_11),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_223),
.A2(n_12),
.B(n_13),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_225),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_221),
.Y(n_227)
);


endmodule