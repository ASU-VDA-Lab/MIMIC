module fake_ibex_905_n_1917 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_124, n_37, n_256, n_193, n_108, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_88, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_15, n_24, n_189, n_280, n_317, n_340, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_235, n_22, n_136, n_261, n_30, n_221, n_102, n_52, n_99, n_269, n_156, n_126, n_25, n_104, n_45, n_141, n_222, n_186, n_295, n_331, n_230, n_96, n_185, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_335, n_82, n_263, n_27, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_180, n_201, n_14, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_4, n_6, n_100, n_179, n_206, n_329, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_272, n_23, n_223, n_95, n_285, n_288, n_247, n_320, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_118, n_164, n_38, n_198, n_264, n_217, n_324, n_78, n_20, n_69, n_39, n_178, n_303, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_119, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_281, n_1917);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_88;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_221;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_335;
input n_82;
input n_263;
input n_27;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_180;
input n_201;
input n_14;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_4;
input n_6;
input n_100;
input n_179;
input n_206;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_272;
input n_23;
input n_223;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_118;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_119;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_281;

output n_1917;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_1802;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1883;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_369;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_745;
wire n_447;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_579;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_379;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1717;
wire n_1609;
wire n_391;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_395;
wire n_1786;
wire n_1319;
wire n_389;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_1831;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_388;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_363;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_351;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_1470;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_650;
wire n_409;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_1857;
wire n_545;
wire n_887;
wire n_1162;
wire n_1894;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_1830;
wire n_1629;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_1340;
wire n_348;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_370;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_1899;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_1538;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_1889;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_1057;
wire n_354;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_1779;
wire n_360;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_362;
wire n_505;
wire n_1621;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1893;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_387;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_1872;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_1767;
wire n_1768;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1584;
wire n_1481;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1892;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1635;
wire n_1572;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_714;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1397;
wire n_1211;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_1868;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1757;
wire n_699;
wire n_368;
wire n_918;
wire n_1913;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_548;
wire n_1158;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_405;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_414;
wire n_378;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1900;
wire n_519;
wire n_1843;
wire n_408;
wire n_361;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_1902;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

BUFx5_ASAP7_75t_L g345 ( 
.A(n_241),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_35),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_250),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_270),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_293),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_323),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_96),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_60),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_225),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_L g354 ( 
.A(n_55),
.B(n_245),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_185),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_246),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_292),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_117),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_251),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_168),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_202),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_271),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_213),
.Y(n_363)
);

BUFx5_ASAP7_75t_L g364 ( 
.A(n_318),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_222),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_266),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_184),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_199),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_71),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_90),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_215),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_272),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_102),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_306),
.Y(n_374)
);

BUFx8_ASAP7_75t_SL g375 ( 
.A(n_175),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_248),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_163),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_147),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_9),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_55),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_255),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_141),
.Y(n_382)
);

INVxp33_ASAP7_75t_L g383 ( 
.A(n_85),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_329),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_313),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_122),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_321),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_38),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_300),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_104),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_279),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_218),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_274),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_233),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_13),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_334),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_63),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_310),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_217),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_106),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_122),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_295),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_73),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_31),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_1),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_204),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_261),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_332),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_105),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_70),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_31),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_94),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_286),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_98),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_210),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_214),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_11),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_269),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_309),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_198),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_171),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_74),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_312),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_21),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_227),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_208),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_97),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_224),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_264),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_111),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_117),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_13),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_284),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_71),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_307),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_229),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_324),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_83),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_340),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_108),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_326),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_287),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_253),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_120),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_308),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_235),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_190),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_30),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_265),
.Y(n_449)
);

CKINVDCx14_ASAP7_75t_R g450 ( 
.A(n_128),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_180),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_113),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_216),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g454 ( 
.A(n_109),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_110),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_136),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_194),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_41),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_177),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_76),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_260),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_231),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_333),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_296),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_77),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_151),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_302),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_90),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_63),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_277),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_100),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_311),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_341),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_136),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_317),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_124),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_337),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_280),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_130),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_148),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_59),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_339),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_6),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_316),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_61),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_335),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_196),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_189),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_100),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_178),
.Y(n_490)
);

BUFx8_ASAP7_75t_SL g491 ( 
.A(n_273),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_195),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_155),
.Y(n_493)
);

BUFx5_ASAP7_75t_L g494 ( 
.A(n_283),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_249),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_143),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_219),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_30),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_85),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_110),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_197),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_282),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_325),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_221),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_232),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_7),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_181),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_108),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_38),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_303),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_205),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_259),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_182),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_342),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_226),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_29),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_240),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_228),
.Y(n_518)
);

BUFx8_ASAP7_75t_SL g519 ( 
.A(n_234),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_220),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_16),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_344),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_297),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_87),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_58),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_80),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_247),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_68),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_65),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_243),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_14),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_57),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_285),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_238),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_254),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_105),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_111),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_191),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_73),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_294),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_252),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_212),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_244),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_5),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_104),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_130),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_32),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_49),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_20),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_338),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_87),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_169),
.Y(n_552)
);

INVx1_ASAP7_75t_SL g553 ( 
.A(n_47),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_298),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_134),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_157),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_4),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_288),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_201),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_176),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_120),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_67),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_159),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_343),
.Y(n_564)
);

CKINVDCx14_ASAP7_75t_R g565 ( 
.A(n_44),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_18),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_91),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_29),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_47),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_19),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_236),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_33),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_262),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_92),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_19),
.Y(n_575)
);

BUFx5_ASAP7_75t_L g576 ( 
.A(n_50),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_51),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_45),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_86),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_304),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_148),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_268),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_242),
.Y(n_583)
);

BUFx10_ASAP7_75t_L g584 ( 
.A(n_128),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_336),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_211),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_51),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_267),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_152),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_43),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_124),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_558),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_450),
.Y(n_593)
);

AOI22x1_ASAP7_75t_SL g594 ( 
.A1(n_465),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_450),
.Y(n_595)
);

BUFx8_ASAP7_75t_SL g596 ( 
.A(n_465),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_376),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_431),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_454),
.A2(n_565),
.B1(n_392),
.B2(n_406),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_454),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_376),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_565),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_558),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_383),
.B(n_3),
.Y(n_604)
);

BUFx8_ASAP7_75t_SL g605 ( 
.A(n_521),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_431),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_376),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_572),
.Y(n_608)
);

NOR2x1_ASAP7_75t_L g609 ( 
.A(n_555),
.B(n_153),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_376),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_576),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_SL g612 ( 
.A1(n_521),
.A2(n_575),
.B1(n_378),
.B2(n_388),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_576),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_555),
.Y(n_614)
);

OAI22x1_ASAP7_75t_R g615 ( 
.A1(n_575),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_414),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_363),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_420),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_383),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_394),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_420),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_501),
.Y(n_622)
);

OA21x2_ASAP7_75t_L g623 ( 
.A1(n_413),
.A2(n_156),
.B(n_154),
.Y(n_623)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_420),
.Y(n_624)
);

NOR2x1_ASAP7_75t_L g625 ( 
.A(n_495),
.B(n_158),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_518),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_556),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_576),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_572),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_438),
.Y(n_630)
);

OA21x2_ASAP7_75t_L g631 ( 
.A1(n_413),
.A2(n_161),
.B(n_160),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_438),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_466),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_515),
.B(n_10),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_349),
.Y(n_635)
);

AND2x6_ASAP7_75t_L g636 ( 
.A(n_433),
.B(n_162),
.Y(n_636)
);

CKINVDCx16_ASAP7_75t_R g637 ( 
.A(n_365),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_468),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g639 ( 
.A(n_468),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_576),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_425),
.B(n_10),
.Y(n_641)
);

OAI22x1_ASAP7_75t_R g642 ( 
.A1(n_380),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_397),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_397),
.B(n_12),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_422),
.Y(n_645)
);

OAI22x1_ASAP7_75t_SL g646 ( 
.A1(n_496),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_422),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_369),
.Y(n_648)
);

OA21x2_ASAP7_75t_L g649 ( 
.A1(n_425),
.A2(n_165),
.B(n_164),
.Y(n_649)
);

OAI21x1_ASAP7_75t_L g650 ( 
.A1(n_436),
.A2(n_167),
.B(n_166),
.Y(n_650)
);

BUFx12f_ASAP7_75t_L g651 ( 
.A(n_572),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_576),
.B(n_17),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_369),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_369),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_346),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_375),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_584),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_369),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_440),
.Y(n_659)
);

BUFx8_ASAP7_75t_SL g660 ( 
.A(n_375),
.Y(n_660)
);

BUFx8_ASAP7_75t_SL g661 ( 
.A(n_491),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_504),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_491),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_506),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_351),
.B(n_18),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_506),
.Y(n_666)
);

INVx5_ASAP7_75t_L g667 ( 
.A(n_504),
.Y(n_667)
);

BUFx12f_ASAP7_75t_L g668 ( 
.A(n_352),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_506),
.Y(n_669)
);

INVx5_ASAP7_75t_L g670 ( 
.A(n_520),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_506),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_520),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_SL g673 ( 
.A1(n_499),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_673)
);

BUFx12f_ASAP7_75t_L g674 ( 
.A(n_358),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_480),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_350),
.Y(n_676)
);

AO22x2_ASAP7_75t_L g677 ( 
.A1(n_590),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_382),
.B(n_25),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_436),
.A2(n_172),
.B(n_170),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_562),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_534),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_562),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_353),
.Y(n_683)
);

NOR2x1_ASAP7_75t_L g684 ( 
.A(n_386),
.B(n_173),
.Y(n_684)
);

BUFx8_ASAP7_75t_SL g685 ( 
.A(n_519),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_395),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_562),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_373),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_345),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_562),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_619),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_651),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_597),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_644),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_660),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_619),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_600),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_614),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_637),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_R g700 ( 
.A(n_656),
.B(n_663),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_597),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_661),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_661),
.Y(n_703)
);

AND2x6_ASAP7_75t_L g704 ( 
.A(n_609),
.B(n_534),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_593),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_685),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_685),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_596),
.Y(n_708)
);

AOI21x1_ASAP7_75t_L g709 ( 
.A1(n_611),
.A2(n_457),
.B(n_445),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_643),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_643),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_647),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_R g713 ( 
.A(n_629),
.B(n_356),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_605),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_668),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_674),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_R g717 ( 
.A(n_595),
.B(n_356),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_R g718 ( 
.A(n_629),
.B(n_402),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_655),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_599),
.A2(n_512),
.B1(n_517),
.B2(n_467),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_R g721 ( 
.A(n_657),
.B(n_402),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_612),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_688),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_604),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_630),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_R g726 ( 
.A(n_657),
.B(n_473),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_635),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_R g728 ( 
.A(n_608),
.B(n_473),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_676),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_676),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_598),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_R g732 ( 
.A(n_620),
.B(n_622),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_683),
.Y(n_733)
);

AND3x2_ASAP7_75t_L g734 ( 
.A(n_617),
.B(n_370),
.C(n_387),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_688),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_617),
.B(n_443),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_626),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_616),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_606),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_662),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_672),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_615),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_627),
.B(n_445),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_632),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_632),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_R g746 ( 
.A(n_636),
.B(n_467),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_633),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_633),
.B(n_638),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_638),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_639),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_642),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_681),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_594),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_646),
.Y(n_754)
);

XOR2xp5_ASAP7_75t_L g755 ( 
.A(n_602),
.B(n_512),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_673),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_SL g757 ( 
.A(n_634),
.B(n_517),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_686),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_659),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_659),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_678),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_592),
.B(n_457),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_665),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_597),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_652),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_625),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_592),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_675),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_675),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_641),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_613),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_645),
.B(n_379),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_603),
.B(n_390),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_641),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_628),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_640),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_603),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_636),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_636),
.Y(n_779)
);

AND3x2_ASAP7_75t_L g780 ( 
.A(n_677),
.B(n_410),
.C(n_403),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_677),
.A2(n_589),
.B1(n_573),
.B2(n_401),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_677),
.A2(n_589),
.B1(n_573),
.B2(n_404),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_684),
.B(n_412),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_689),
.Y(n_784)
);

NOR2xp67_ASAP7_75t_L g785 ( 
.A(n_667),
.B(n_348),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_667),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_667),
.Y(n_787)
);

INVx1_ASAP7_75t_SL g788 ( 
.A(n_667),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_690),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_670),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_670),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_670),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_690),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_618),
.B(n_400),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_618),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_618),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_650),
.Y(n_797)
);

AND2x6_ASAP7_75t_L g798 ( 
.A(n_597),
.B(n_464),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_679),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_648),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_624),
.Y(n_801)
);

NOR2xp67_ASAP7_75t_L g802 ( 
.A(n_624),
.B(n_355),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_648),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_623),
.Y(n_804)
);

INVxp33_ASAP7_75t_SL g805 ( 
.A(n_623),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_648),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_653),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_653),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_653),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_654),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_654),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_687),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_658),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_687),
.B(n_516),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_687),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_658),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_658),
.Y(n_817)
);

NAND2xp33_ASAP7_75t_R g818 ( 
.A(n_631),
.B(n_405),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_682),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_664),
.B(n_417),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_664),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_666),
.B(n_464),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_666),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_631),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_631),
.Y(n_825)
);

INVxp67_ASAP7_75t_SL g826 ( 
.A(n_649),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_601),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_669),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_669),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_601),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_669),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_671),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_671),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_649),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_671),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_680),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_R g837 ( 
.A(n_680),
.B(n_511),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_698),
.B(n_347),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_758),
.B(n_359),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_789),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_814),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_691),
.B(n_409),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_731),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_724),
.B(n_649),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_694),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_691),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_696),
.B(n_411),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_694),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_763),
.B(n_360),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_R g850 ( 
.A(n_715),
.B(n_585),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_724),
.B(n_357),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_727),
.B(n_362),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_747),
.B(n_361),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_729),
.B(n_366),
.Y(n_854)
);

OA21x2_ASAP7_75t_L g855 ( 
.A1(n_797),
.A2(n_482),
.B(n_475),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_759),
.B(n_367),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_692),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_760),
.B(n_748),
.Y(n_858)
);

INVx8_ASAP7_75t_L g859 ( 
.A(n_767),
.Y(n_859)
);

NOR3xp33_ASAP7_75t_L g860 ( 
.A(n_720),
.B(n_553),
.C(n_537),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_696),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_697),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_770),
.B(n_368),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_774),
.B(n_371),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_697),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_752),
.B(n_372),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_730),
.B(n_374),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_750),
.B(n_424),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_733),
.B(n_377),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_735),
.B(n_427),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_732),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_L g872 ( 
.A(n_818),
.B(n_384),
.C(n_381),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_735),
.B(n_430),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_820),
.Y(n_874)
);

NOR2xp67_ASAP7_75t_L g875 ( 
.A(n_716),
.B(n_26),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_732),
.Y(n_876)
);

AOI221xp5_ASAP7_75t_L g877 ( 
.A1(n_710),
.A2(n_455),
.B1(n_458),
.B2(n_452),
.C(n_432),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_711),
.B(n_712),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_736),
.B(n_434),
.Y(n_879)
);

INVxp67_ASAP7_75t_SL g880 ( 
.A(n_737),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_705),
.Y(n_881)
);

NAND3xp33_ASAP7_75t_L g882 ( 
.A(n_818),
.B(n_391),
.C(n_385),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_738),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_783),
.B(n_393),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_713),
.B(n_389),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_779),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_784),
.B(n_398),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_725),
.B(n_407),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_699),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_740),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_741),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_762),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_768),
.B(n_416),
.Y(n_893)
);

BUFx5_ASAP7_75t_L g894 ( 
.A(n_798),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_744),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_769),
.B(n_766),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_709),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_739),
.B(n_419),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_745),
.B(n_444),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_761),
.B(n_426),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_762),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_822),
.Y(n_902)
);

OR2x2_ASAP7_75t_L g903 ( 
.A(n_719),
.B(n_448),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_749),
.B(n_428),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_822),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_793),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_772),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_743),
.B(n_429),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_704),
.B(n_805),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_704),
.B(n_396),
.Y(n_910)
);

NAND2xp33_ASAP7_75t_SL g911 ( 
.A(n_713),
.B(n_456),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_704),
.B(n_399),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_773),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_785),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_802),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_708),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_717),
.B(n_460),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_780),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_L g919 ( 
.A(n_746),
.B(n_345),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_704),
.B(n_408),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_804),
.B(n_415),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_794),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_806),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_807),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_808),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_804),
.B(n_824),
.Y(n_926)
);

INVx8_ASAP7_75t_L g927 ( 
.A(n_777),
.Y(n_927)
);

AND3x2_ASAP7_75t_L g928 ( 
.A(n_751),
.B(n_476),
.C(n_471),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_824),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_826),
.B(n_418),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_811),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_721),
.B(n_441),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_726),
.B(n_718),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_728),
.B(n_447),
.Y(n_934)
);

INVx8_ASAP7_75t_L g935 ( 
.A(n_825),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_798),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_771),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_786),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_734),
.B(n_451),
.Y(n_939)
);

AO21x2_ASAP7_75t_L g940 ( 
.A1(n_834),
.A2(n_423),
.B(n_421),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_781),
.B(n_453),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_757),
.B(n_459),
.Y(n_942)
);

BUFx6f_ASAP7_75t_SL g943 ( 
.A(n_695),
.Y(n_943)
);

BUFx6f_ASAP7_75t_SL g944 ( 
.A(n_702),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_782),
.B(n_470),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_775),
.B(n_478),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_755),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_813),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_816),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_776),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_SL g951 ( 
.A(n_798),
.B(n_484),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_788),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_817),
.Y(n_953)
);

NOR3xp33_ASAP7_75t_L g954 ( 
.A(n_753),
.B(n_474),
.C(n_469),
.Y(n_954)
);

NOR2xp67_ASAP7_75t_L g955 ( 
.A(n_703),
.B(n_27),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_837),
.B(n_486),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_787),
.B(n_487),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_790),
.B(n_488),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_791),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_792),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_700),
.B(n_481),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_821),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_700),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_829),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_832),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_795),
.B(n_490),
.Y(n_966)
);

INVx8_ASAP7_75t_L g967 ( 
.A(n_798),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_833),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_796),
.B(n_492),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_801),
.B(n_435),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_835),
.B(n_497),
.Y(n_971)
);

NAND2xp33_ASAP7_75t_L g972 ( 
.A(n_798),
.B(n_345),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_836),
.B(n_503),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_714),
.B(n_513),
.Y(n_974)
);

OR2x6_ASAP7_75t_L g975 ( 
.A(n_706),
.B(n_479),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_800),
.B(n_514),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_810),
.B(n_522),
.Y(n_977)
);

INVx8_ASAP7_75t_L g978 ( 
.A(n_707),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_812),
.B(n_523),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_815),
.B(n_527),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_819),
.B(n_530),
.Y(n_981)
);

NAND3xp33_ASAP7_75t_L g982 ( 
.A(n_823),
.B(n_439),
.C(n_437),
.Y(n_982)
);

AO221x1_ASAP7_75t_L g983 ( 
.A1(n_742),
.A2(n_508),
.B1(n_524),
.B2(n_498),
.C(n_485),
.Y(n_983)
);

AO221x1_ASAP7_75t_L g984 ( 
.A1(n_722),
.A2(n_544),
.B1(n_547),
.B2(n_531),
.C(n_526),
.Y(n_984)
);

NAND3xp33_ASAP7_75t_L g985 ( 
.A(n_828),
.B(n_446),
.C(n_442),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_756),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_754),
.B(n_483),
.Y(n_987)
);

OR2x6_ASAP7_75t_L g988 ( 
.A(n_803),
.B(n_548),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_693),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_693),
.B(n_533),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_831),
.B(n_489),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_693),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_809),
.B(n_540),
.Y(n_993)
);

BUFx6f_ASAP7_75t_SL g994 ( 
.A(n_701),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_701),
.B(n_541),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_701),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_701),
.B(n_500),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_764),
.B(n_542),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_764),
.B(n_550),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_764),
.B(n_509),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_827),
.B(n_559),
.Y(n_1001)
);

NOR2xp67_ASAP7_75t_L g1002 ( 
.A(n_830),
.B(n_28),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_R g1003 ( 
.A(n_715),
.B(n_525),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_758),
.B(n_563),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_778),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_765),
.B(n_449),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_814),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_765),
.B(n_461),
.Y(n_1008)
);

OR2x6_ASAP7_75t_L g1009 ( 
.A(n_692),
.B(n_549),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_814),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_789),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_814),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_789),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_846),
.B(n_528),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_861),
.B(n_529),
.Y(n_1015)
);

AO22x1_ASAP7_75t_L g1016 ( 
.A1(n_880),
.A2(n_536),
.B1(n_539),
.B2(n_532),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_862),
.B(n_569),
.Y(n_1017)
);

NOR3xp33_ASAP7_75t_SL g1018 ( 
.A(n_941),
.B(n_546),
.C(n_545),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_865),
.B(n_551),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_845),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_927),
.Y(n_1021)
);

OR2x6_ASAP7_75t_L g1022 ( 
.A(n_978),
.B(n_578),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_848),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_879),
.A2(n_907),
.B1(n_858),
.B2(n_878),
.Y(n_1024)
);

BUFx12f_ASAP7_75t_SL g1025 ( 
.A(n_1009),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_881),
.B(n_557),
.Y(n_1026)
);

INVx5_ASAP7_75t_L g1027 ( 
.A(n_967),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_850),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_895),
.B(n_561),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1006),
.B(n_566),
.Y(n_1030)
);

INVx1_ASAP7_75t_SL g1031 ( 
.A(n_903),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_967),
.Y(n_1032)
);

INVxp67_ASAP7_75t_SL g1033 ( 
.A(n_926),
.Y(n_1033)
);

NAND2x1p5_ASAP7_75t_L g1034 ( 
.A(n_857),
.B(n_579),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_870),
.A2(n_568),
.B1(n_570),
.B2(n_567),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_1009),
.Y(n_1036)
);

NAND2x1p5_ASAP7_75t_L g1037 ( 
.A(n_871),
.B(n_354),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_927),
.Y(n_1038)
);

NAND2xp33_ASAP7_75t_L g1039 ( 
.A(n_926),
.B(n_345),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_967),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1006),
.B(n_1008),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_841),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_876),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_873),
.A2(n_577),
.B1(n_581),
.B2(n_574),
.Y(n_1044)
);

INVx5_ASAP7_75t_L g1045 ( 
.A(n_936),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1007),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_883),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1010),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_842),
.A2(n_591),
.B1(n_587),
.B2(n_462),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_927),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_847),
.A2(n_463),
.B1(n_477),
.B2(n_472),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_868),
.B(n_28),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_936),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1012),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_936),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_906),
.B(n_493),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_874),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_899),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_844),
.A2(n_505),
.B(n_507),
.C(n_502),
.Y(n_1059)
);

BUFx2_ASAP7_75t_SL g1060 ( 
.A(n_943),
.Y(n_1060)
);

BUFx4f_ASAP7_75t_L g1061 ( 
.A(n_978),
.Y(n_1061)
);

INVx8_ASAP7_75t_L g1062 ( 
.A(n_978),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_963),
.B(n_510),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_886),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_843),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_991),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_853),
.B(n_571),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_889),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_890),
.Y(n_1069)
);

AND2x2_ASAP7_75t_SL g1070 ( 
.A(n_860),
.B(n_535),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_859),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_945),
.A2(n_543),
.B1(n_552),
.B2(n_538),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_1003),
.Y(n_1073)
);

OAI21xp33_ASAP7_75t_L g1074 ( 
.A1(n_838),
.A2(n_582),
.B(n_580),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_859),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_884),
.B(n_586),
.Y(n_1076)
);

AND2x6_ASAP7_75t_L g1077 ( 
.A(n_929),
.B(n_554),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_884),
.B(n_588),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_961),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_859),
.Y(n_1080)
);

INVxp67_ASAP7_75t_SL g1081 ( 
.A(n_930),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_997),
.Y(n_1082)
);

NOR3xp33_ASAP7_75t_L g1083 ( 
.A(n_947),
.B(n_564),
.C(n_560),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_959),
.B(n_960),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1000),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_891),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_916),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_886),
.Y(n_1088)
);

OR2x2_ASAP7_75t_L g1089 ( 
.A(n_986),
.B(n_34),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_851),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_937),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_918),
.B(n_583),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_938),
.Y(n_1093)
);

INVx5_ASAP7_75t_L g1094 ( 
.A(n_938),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_950),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_917),
.Y(n_1096)
);

INVx8_ASAP7_75t_L g1097 ( 
.A(n_975),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_975),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_975),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_892),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_901),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_952),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_844),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_900),
.B(n_34),
.Y(n_1104)
);

CKINVDCx8_ASAP7_75t_R g1105 ( 
.A(n_935),
.Y(n_1105)
);

AND2x6_ASAP7_75t_SL g1106 ( 
.A(n_987),
.B(n_36),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_1005),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_922),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_943),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_913),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_863),
.B(n_364),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_872),
.A2(n_494),
.B1(n_364),
.B2(n_680),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_840),
.Y(n_1113)
);

AND3x1_ASAP7_75t_L g1114 ( 
.A(n_954),
.B(n_36),
.C(n_37),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_872),
.A2(n_494),
.B1(n_682),
.B2(n_607),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_864),
.B(n_494),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_904),
.B(n_37),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_882),
.A2(n_494),
.B1(n_607),
.B2(n_601),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_1005),
.Y(n_1119)
);

BUFx8_ASAP7_75t_L g1120 ( 
.A(n_944),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1011),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_908),
.B(n_494),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_962),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_935),
.Y(n_1124)
);

OR2x6_ASAP7_75t_L g1125 ( 
.A(n_935),
.B(n_39),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_964),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1013),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_921),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_921),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_930),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_902),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_905),
.Y(n_1132)
);

OR2x2_ASAP7_75t_SL g1133 ( 
.A(n_944),
.B(n_39),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_914),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_989),
.Y(n_1135)
);

INVx8_ASAP7_75t_L g1136 ( 
.A(n_988),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_942),
.B(n_40),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_855),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_994),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_915),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_965),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_897),
.A2(n_621),
.B(n_610),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_910),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_898),
.B(n_42),
.Y(n_1144)
);

BUFx4f_ASAP7_75t_L g1145 ( 
.A(n_988),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_910),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_928),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_896),
.B(n_44),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_R g1149 ( 
.A(n_911),
.B(n_45),
.Y(n_1149)
);

OAI22xp33_ASAP7_75t_SL g1150 ( 
.A1(n_933),
.A2(n_50),
.B1(n_46),
.B2(n_48),
.Y(n_1150)
);

INVx2_ASAP7_75t_SL g1151 ( 
.A(n_856),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_888),
.B(n_46),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_887),
.B(n_877),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_912),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_994),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_989),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_912),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_988),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_893),
.Y(n_1159)
);

OR2x6_ASAP7_75t_L g1160 ( 
.A(n_875),
.B(n_52),
.Y(n_1160)
);

BUFx10_ASAP7_75t_L g1161 ( 
.A(n_974),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_855),
.A2(n_999),
.B(n_998),
.Y(n_1162)
);

OR2x6_ASAP7_75t_L g1163 ( 
.A(n_955),
.B(n_52),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_849),
.B(n_53),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_923),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_970),
.B(n_54),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_909),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_839),
.B(n_62),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_970),
.B(n_62),
.Y(n_1169)
);

OR2x6_ASAP7_75t_L g1170 ( 
.A(n_1004),
.B(n_64),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_920),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_866),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_924),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_940),
.B(n_65),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_925),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_940),
.B(n_934),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_946),
.B(n_66),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_951),
.B(n_66),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_931),
.Y(n_1179)
);

OR2x6_ASAP7_75t_L g1180 ( 
.A(n_939),
.B(n_67),
.Y(n_1180)
);

OR2x2_ASAP7_75t_SL g1181 ( 
.A(n_983),
.B(n_984),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_948),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_949),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_957),
.B(n_69),
.Y(n_1184)
);

AND2x2_ASAP7_75t_SL g1185 ( 
.A(n_919),
.B(n_70),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_958),
.B(n_72),
.Y(n_1186)
);

INVx2_ASAP7_75t_SL g1187 ( 
.A(n_953),
.Y(n_1187)
);

OR2x6_ASAP7_75t_L g1188 ( 
.A(n_852),
.B(n_72),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_854),
.B(n_74),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_R g1190 ( 
.A(n_951),
.B(n_75),
.Y(n_1190)
);

OAI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_966),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_968),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1002),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_894),
.Y(n_1194)
);

INVxp67_ASAP7_75t_L g1195 ( 
.A(n_969),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_982),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_867),
.B(n_78),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_869),
.B(n_79),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1062),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1145),
.B(n_971),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1108),
.Y(n_1201)
);

AND2x4_ASAP7_75t_SL g1202 ( 
.A(n_1021),
.B(n_989),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_R g1203 ( 
.A(n_1025),
.B(n_972),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1090),
.B(n_885),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1031),
.B(n_956),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_1036),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1081),
.A2(n_973),
.B1(n_932),
.B2(n_982),
.Y(n_1207)
);

NOR2xp67_ASAP7_75t_L g1208 ( 
.A(n_1021),
.B(n_1038),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1110),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1103),
.A2(n_977),
.B(n_976),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1058),
.B(n_979),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1128),
.A2(n_985),
.B(n_980),
.C(n_981),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_1062),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1079),
.B(n_990),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1070),
.A2(n_995),
.B1(n_993),
.B2(n_1001),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1061),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_SL g1217 ( 
.A1(n_1133),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1042),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1130),
.B(n_84),
.Y(n_1219)
);

BUFx12f_ASAP7_75t_L g1220 ( 
.A(n_1120),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_R g1221 ( 
.A(n_1087),
.B(n_84),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1181),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_1222)
);

NAND2xp33_ASAP7_75t_L g1223 ( 
.A(n_1077),
.B(n_1128),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1136),
.Y(n_1224)
);

INVxp33_ASAP7_75t_SL g1225 ( 
.A(n_1073),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1096),
.B(n_91),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1061),
.Y(n_1227)
);

CKINVDCx11_ASAP7_75t_R g1228 ( 
.A(n_1097),
.Y(n_1228)
);

AO21x1_ASAP7_75t_L g1229 ( 
.A1(n_1174),
.A2(n_1178),
.B(n_1039),
.Y(n_1229)
);

OAI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1196),
.A2(n_996),
.B(n_992),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1117),
.A2(n_1132),
.B(n_1131),
.C(n_1172),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_SL g1232 ( 
.A1(n_1125),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_1232)
);

NOR2xp67_ASAP7_75t_SL g1233 ( 
.A(n_1060),
.B(n_996),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1155),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1046),
.Y(n_1235)
);

CKINVDCx16_ASAP7_75t_R g1236 ( 
.A(n_1022),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1122),
.A2(n_179),
.B(n_174),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1136),
.Y(n_1238)
);

NOR3xp33_ASAP7_75t_SL g1239 ( 
.A(n_1109),
.B(n_93),
.C(n_97),
.Y(n_1239)
);

BUFx4f_ASAP7_75t_L g1240 ( 
.A(n_1097),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1048),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1054),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1022),
.Y(n_1243)
);

INVx5_ASAP7_75t_L g1244 ( 
.A(n_1155),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1131),
.A2(n_1132),
.B(n_1100),
.C(n_1101),
.Y(n_1245)
);

INVxp67_ASAP7_75t_L g1246 ( 
.A(n_1098),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1111),
.A2(n_186),
.B(n_183),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1099),
.B(n_98),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1059),
.A2(n_99),
.B(n_101),
.C(n_103),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1158),
.B(n_99),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1158),
.B(n_101),
.Y(n_1251)
);

O2A1O1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1166),
.A2(n_103),
.B(n_107),
.C(n_112),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1027),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1125),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1116),
.A2(n_188),
.B(n_187),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1148),
.A2(n_107),
.B(n_112),
.C(n_113),
.Y(n_1256)
);

O2A1O1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1169),
.A2(n_114),
.B(n_115),
.C(n_116),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1024),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1185),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1135),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1066),
.B(n_1017),
.Y(n_1261)
);

AOI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1162),
.A2(n_1193),
.B(n_1142),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1019),
.B(n_118),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1034),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1050),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1017),
.B(n_119),
.Y(n_1266)
);

NOR2xp67_ASAP7_75t_SL g1267 ( 
.A(n_1105),
.B(n_121),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1030),
.B(n_123),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1159),
.B(n_123),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1196),
.A2(n_193),
.B(n_192),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_1068),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1102),
.B(n_125),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1035),
.B(n_125),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1044),
.B(n_1052),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1195),
.B(n_126),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1152),
.A2(n_1146),
.B(n_1154),
.C(n_1143),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1157),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1026),
.B(n_129),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1120),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1028),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1083),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_1281)
);

OA22x2_ASAP7_75t_L g1282 ( 
.A1(n_1170),
.A2(n_1188),
.B1(n_1180),
.B2(n_1147),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1077),
.Y(n_1283)
);

INVx5_ASAP7_75t_L g1284 ( 
.A(n_1139),
.Y(n_1284)
);

BUFx12f_ASAP7_75t_L g1285 ( 
.A(n_1106),
.Y(n_1285)
);

INVx4_ASAP7_75t_L g1286 ( 
.A(n_1027),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1082),
.A2(n_132),
.B(n_133),
.C(n_134),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1171),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1091),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1085),
.A2(n_135),
.B(n_137),
.C(n_138),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1164),
.A2(n_1168),
.B1(n_1197),
.B2(n_1189),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1137),
.A2(n_139),
.B(n_140),
.C(n_141),
.Y(n_1292)
);

OAI22x1_ASAP7_75t_L g1293 ( 
.A1(n_1164),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.Y(n_1293)
);

BUFx8_ASAP7_75t_L g1294 ( 
.A(n_1071),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1095),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1191),
.A2(n_142),
.B(n_143),
.C(n_144),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1168),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1150),
.A2(n_145),
.B(n_146),
.C(n_147),
.Y(n_1298)
);

INVx4_ASAP7_75t_L g1299 ( 
.A(n_1027),
.Y(n_1299)
);

AND2x6_ASAP7_75t_SL g1300 ( 
.A(n_1170),
.B(n_149),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1047),
.B(n_149),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1151),
.B(n_150),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1188),
.Y(n_1303)
);

NAND2x1_ASAP7_75t_L g1304 ( 
.A(n_1156),
.B(n_1040),
.Y(n_1304)
);

OAI21xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1160),
.A2(n_200),
.B(n_203),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1040),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1189),
.A2(n_206),
.B1(n_207),
.B2(n_209),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1029),
.B(n_223),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1065),
.Y(n_1309)
);

BUFx12f_ASAP7_75t_L g1310 ( 
.A(n_1075),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1069),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1057),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1020),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_R g1314 ( 
.A(n_1080),
.B(n_230),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1016),
.B(n_237),
.Y(n_1315)
);

OR2x6_ASAP7_75t_L g1316 ( 
.A(n_1124),
.B(n_239),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_SL g1317 ( 
.A1(n_1114),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.Y(n_1317)
);

NOR2x1_ASAP7_75t_L g1318 ( 
.A(n_1160),
.B(n_263),
.Y(n_1318)
);

INVx2_ASAP7_75t_SL g1319 ( 
.A(n_1094),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_1149),
.B(n_275),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1093),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1051),
.B(n_276),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1112),
.A2(n_278),
.B(n_281),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1077),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1156),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1023),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1053),
.Y(n_1327)
);

INVx6_ASAP7_75t_L g1328 ( 
.A(n_1084),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1084),
.B(n_289),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1018),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1049),
.B(n_290),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1064),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1067),
.A2(n_1078),
.B(n_1076),
.Y(n_1333)
);

NAND2xp33_ASAP7_75t_L g1334 ( 
.A(n_1077),
.B(n_291),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1179),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1014),
.B(n_299),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1056),
.B(n_301),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1015),
.B(n_305),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1056),
.B(n_1180),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1173),
.B(n_1175),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1053),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1063),
.B(n_314),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1123),
.B(n_315),
.Y(n_1343)
);

INVx1_ASAP7_75t_SL g1344 ( 
.A(n_1184),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1184),
.A2(n_319),
.B1(n_320),
.B2(n_322),
.Y(n_1345)
);

A2O1A1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1177),
.A2(n_327),
.B(n_328),
.C(n_330),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1063),
.B(n_331),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1190),
.Y(n_1348)
);

AOI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1186),
.A2(n_1092),
.B1(n_1104),
.B2(n_1144),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1183),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1053),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1089),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1086),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1126),
.B(n_1141),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1163),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_SL g1356 ( 
.A(n_1045),
.B(n_1161),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1182),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_R g1358 ( 
.A(n_1161),
.B(n_1043),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1192),
.B(n_1187),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1113),
.A2(n_1127),
.B(n_1121),
.Y(n_1360)
);

BUFx2_ASAP7_75t_SL g1361 ( 
.A(n_1045),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1092),
.B(n_1072),
.Y(n_1362)
);

INVxp33_ASAP7_75t_L g1363 ( 
.A(n_1037),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1165),
.B(n_1140),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1074),
.A2(n_1198),
.B1(n_1165),
.B2(n_1167),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_R g1366 ( 
.A(n_1088),
.B(n_1107),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1134),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1088),
.A2(n_1119),
.B1(n_1032),
.B2(n_1045),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1115),
.A2(n_1118),
.B1(n_1194),
.B2(n_1055),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1055),
.B(n_1194),
.Y(n_1370)
);

AOI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1176),
.A2(n_1138),
.B(n_799),
.Y(n_1371)
);

A2O1A1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1041),
.A2(n_1128),
.B(n_1129),
.C(n_1130),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1108),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1031),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1041),
.A2(n_805),
.B(n_826),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1108),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1031),
.B(n_1058),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1081),
.A2(n_1033),
.B1(n_1130),
.B2(n_1041),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1090),
.B(n_1041),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1062),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1041),
.A2(n_805),
.B(n_826),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1031),
.B(n_1058),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1041),
.A2(n_1128),
.B(n_1129),
.C(n_1130),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1041),
.A2(n_805),
.B(n_826),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1041),
.A2(n_926),
.B(n_929),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1041),
.A2(n_805),
.B(n_826),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1041),
.A2(n_805),
.B(n_826),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1090),
.B(n_1041),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1041),
.A2(n_805),
.B(n_826),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1041),
.A2(n_805),
.B(n_826),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1062),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1031),
.B(n_1058),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1108),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1041),
.A2(n_805),
.B(n_826),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1025),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1090),
.B(n_1041),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1155),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1041),
.A2(n_805),
.B(n_826),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1041),
.A2(n_805),
.B(n_826),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1145),
.B(n_862),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1062),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1041),
.A2(n_1128),
.B(n_1129),
.C(n_1130),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1135),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1145),
.B(n_862),
.Y(n_1404)
);

O2A1O1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1041),
.A2(n_1153),
.B(n_1059),
.C(n_858),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1041),
.A2(n_926),
.B(n_929),
.Y(n_1406)
);

OR2x6_ASAP7_75t_L g1407 ( 
.A(n_1136),
.B(n_1062),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1031),
.B(n_691),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1033),
.A2(n_723),
.B1(n_865),
.B2(n_862),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1408),
.B(n_1374),
.Y(n_1410)
);

INVx5_ASAP7_75t_L g1411 ( 
.A(n_1407),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1379),
.B(n_1388),
.Y(n_1412)
);

BUFx4f_ASAP7_75t_L g1413 ( 
.A(n_1220),
.Y(n_1413)
);

INVx6_ASAP7_75t_L g1414 ( 
.A(n_1294),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1372),
.A2(n_1402),
.B(n_1383),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1201),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1228),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1270),
.A2(n_1323),
.B(n_1229),
.Y(n_1418)
);

BUFx5_ASAP7_75t_L g1419 ( 
.A(n_1353),
.Y(n_1419)
);

NAND2x1p5_ASAP7_75t_L g1420 ( 
.A(n_1240),
.B(n_1253),
.Y(n_1420)
);

AO21x2_ASAP7_75t_L g1421 ( 
.A1(n_1231),
.A2(n_1276),
.B(n_1212),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1373),
.Y(n_1422)
);

INVx5_ASAP7_75t_L g1423 ( 
.A(n_1407),
.Y(n_1423)
);

OAI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1375),
.A2(n_1384),
.B(n_1381),
.Y(n_1424)
);

BUFx8_ASAP7_75t_L g1425 ( 
.A(n_1279),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1253),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1396),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1208),
.B(n_1407),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1391),
.B(n_1401),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1376),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1393),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1370),
.A2(n_1304),
.B(n_1210),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1378),
.A2(n_1223),
.B(n_1333),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1218),
.Y(n_1434)
);

INVx5_ASAP7_75t_L g1435 ( 
.A(n_1236),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1286),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1286),
.Y(n_1437)
);

BUFx12f_ASAP7_75t_L g1438 ( 
.A(n_1199),
.Y(n_1438)
);

CKINVDCx20_ASAP7_75t_R g1439 ( 
.A(n_1213),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1332),
.A2(n_1255),
.B(n_1247),
.Y(n_1440)
);

INVxp67_ASAP7_75t_SL g1441 ( 
.A(n_1260),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_1240),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1244),
.B(n_1216),
.Y(n_1443)
);

BUFx2_ASAP7_75t_SL g1444 ( 
.A(n_1227),
.Y(n_1444)
);

NAND2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1299),
.B(n_1283),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1244),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_1221),
.Y(n_1447)
);

INVx4_ASAP7_75t_L g1448 ( 
.A(n_1244),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1299),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1409),
.B(n_1377),
.Y(n_1450)
);

CKINVDCx16_ASAP7_75t_R g1451 ( 
.A(n_1314),
.Y(n_1451)
);

OR2x6_ASAP7_75t_L g1452 ( 
.A(n_1316),
.B(n_1361),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1245),
.B(n_1405),
.Y(n_1453)
);

INVx4_ASAP7_75t_L g1454 ( 
.A(n_1316),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1235),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1382),
.B(n_1392),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1264),
.B(n_1339),
.Y(n_1457)
);

INVx4_ASAP7_75t_L g1458 ( 
.A(n_1316),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1332),
.A2(n_1237),
.B(n_1368),
.Y(n_1459)
);

NAND2x1p5_ASAP7_75t_L g1460 ( 
.A(n_1324),
.B(n_1380),
.Y(n_1460)
);

AO21x2_ASAP7_75t_L g1461 ( 
.A1(n_1386),
.A2(n_1389),
.B(n_1387),
.Y(n_1461)
);

INVx4_ASAP7_75t_L g1462 ( 
.A(n_1224),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1366),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1285),
.Y(n_1464)
);

BUFx12f_ASAP7_75t_L g1465 ( 
.A(n_1310),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1202),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_SL g1467 ( 
.A1(n_1318),
.A2(n_1291),
.B(n_1385),
.Y(n_1467)
);

INVx4_ASAP7_75t_L g1468 ( 
.A(n_1238),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1241),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1390),
.A2(n_1398),
.B(n_1394),
.Y(n_1470)
);

OAI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1399),
.A2(n_1406),
.B(n_1219),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1306),
.Y(n_1472)
);

CKINVDCx6p67_ASAP7_75t_R g1473 ( 
.A(n_1395),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1242),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1294),
.Y(n_1475)
);

BUFx6f_ASAP7_75t_SL g1476 ( 
.A(n_1269),
.Y(n_1476)
);

NAND2x1p5_ASAP7_75t_L g1477 ( 
.A(n_1233),
.B(n_1284),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1328),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1268),
.A2(n_1360),
.B(n_1369),
.Y(n_1479)
);

BUFx2_ASAP7_75t_SL g1480 ( 
.A(n_1282),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1306),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1284),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1289),
.Y(n_1483)
);

INVx5_ASAP7_75t_L g1484 ( 
.A(n_1300),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1274),
.B(n_1328),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1295),
.Y(n_1486)
);

BUFx2_ASAP7_75t_L g1487 ( 
.A(n_1243),
.Y(n_1487)
);

BUFx4f_ASAP7_75t_L g1488 ( 
.A(n_1254),
.Y(n_1488)
);

BUFx12f_ASAP7_75t_L g1489 ( 
.A(n_1300),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1335),
.B(n_1273),
.Y(n_1490)
);

INVx5_ASAP7_75t_L g1491 ( 
.A(n_1325),
.Y(n_1491)
);

BUFx12f_ASAP7_75t_L g1492 ( 
.A(n_1280),
.Y(n_1492)
);

AO21x2_ASAP7_75t_L g1493 ( 
.A1(n_1346),
.A2(n_1365),
.B(n_1272),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1234),
.Y(n_1494)
);

BUFx8_ASAP7_75t_L g1495 ( 
.A(n_1348),
.Y(n_1495)
);

INVx5_ASAP7_75t_L g1496 ( 
.A(n_1403),
.Y(n_1496)
);

BUFx2_ASAP7_75t_R g1497 ( 
.A(n_1330),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1261),
.B(n_1344),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1309),
.B(n_1311),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1340),
.Y(n_1500)
);

OAI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1249),
.A2(n_1207),
.B(n_1204),
.Y(n_1501)
);

OA21x2_ASAP7_75t_L g1502 ( 
.A1(n_1292),
.A2(n_1256),
.B(n_1345),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1313),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1321),
.B(n_1352),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1312),
.B(n_1326),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1358),
.Y(n_1506)
);

INVx4_ASAP7_75t_L g1507 ( 
.A(n_1397),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1225),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1303),
.B(n_1271),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1397),
.Y(n_1510)
);

CKINVDCx6p67_ASAP7_75t_R g1511 ( 
.A(n_1355),
.Y(n_1511)
);

AO21x2_ASAP7_75t_L g1512 ( 
.A1(n_1334),
.A2(n_1250),
.B(n_1251),
.Y(n_1512)
);

AO21x2_ASAP7_75t_L g1513 ( 
.A1(n_1322),
.A2(n_1349),
.B(n_1266),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1350),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1206),
.Y(n_1515)
);

INVx4_ASAP7_75t_L g1516 ( 
.A(n_1327),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1362),
.B(n_1205),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1211),
.B(n_1331),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1364),
.Y(n_1519)
);

NOR2xp67_ASAP7_75t_L g1520 ( 
.A(n_1305),
.B(n_1315),
.Y(n_1520)
);

OR2x6_ASAP7_75t_L g1521 ( 
.A(n_1232),
.B(n_1404),
.Y(n_1521)
);

AO21x1_ASAP7_75t_L g1522 ( 
.A1(n_1259),
.A2(n_1252),
.B(n_1257),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1307),
.A2(n_1298),
.B(n_1290),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1265),
.Y(n_1524)
);

OR2x6_ASAP7_75t_L g1525 ( 
.A(n_1232),
.B(n_1400),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1200),
.B(n_1337),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1357),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_SL g1528 ( 
.A1(n_1296),
.A2(n_1319),
.B(n_1297),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1287),
.A2(n_1215),
.B(n_1338),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1293),
.Y(n_1530)
);

AO21x2_ASAP7_75t_L g1531 ( 
.A1(n_1263),
.A2(n_1275),
.B(n_1336),
.Y(n_1531)
);

INVx4_ASAP7_75t_L g1532 ( 
.A(n_1341),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_1342),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1308),
.A2(n_1278),
.B(n_1320),
.Y(n_1534)
);

NAND3xp33_ASAP7_75t_L g1535 ( 
.A(n_1239),
.B(n_1258),
.C(n_1281),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1277),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1288),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1354),
.Y(n_1538)
);

AOI22x1_ASAP7_75t_L g1539 ( 
.A1(n_1347),
.A2(n_1351),
.B1(n_1367),
.B2(n_1246),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1214),
.B(n_1302),
.Y(n_1540)
);

BUFx4f_ASAP7_75t_L g1541 ( 
.A(n_1351),
.Y(n_1541)
);

CKINVDCx8_ASAP7_75t_R g1542 ( 
.A(n_1359),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1226),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1329),
.A2(n_1343),
.B(n_1301),
.Y(n_1544)
);

INVx4_ASAP7_75t_L g1545 ( 
.A(n_1356),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_SL g1546 ( 
.A1(n_1217),
.A2(n_1222),
.B1(n_1363),
.B2(n_1317),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_SL g1547 ( 
.A1(n_1317),
.A2(n_1222),
.B(n_1217),
.Y(n_1547)
);

INVx4_ASAP7_75t_L g1548 ( 
.A(n_1203),
.Y(n_1548)
);

AND2x2_ASAP7_75t_SL g1549 ( 
.A(n_1267),
.B(n_1248),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1391),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1379),
.B(n_1388),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1209),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1209),
.Y(n_1553)
);

AO21x2_ASAP7_75t_L g1554 ( 
.A1(n_1371),
.A2(n_1262),
.B(n_1230),
.Y(n_1554)
);

BUFx2_ASAP7_75t_SL g1555 ( 
.A(n_1391),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1391),
.Y(n_1556)
);

BUFx4f_ASAP7_75t_SL g1557 ( 
.A(n_1220),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1379),
.B(n_1388),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1409),
.B(n_846),
.Y(n_1559)
);

BUFx4f_ASAP7_75t_SL g1560 ( 
.A(n_1220),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1409),
.B(n_846),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1412),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1452),
.B(n_1412),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1551),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1427),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1551),
.B(n_1558),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1558),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1427),
.Y(n_1568)
);

OAI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1501),
.A2(n_1453),
.B(n_1433),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1414),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1452),
.A2(n_1454),
.B1(n_1458),
.B2(n_1546),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_SL g1572 ( 
.A(n_1454),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1452),
.Y(n_1573)
);

INVx6_ASAP7_75t_L g1574 ( 
.A(n_1425),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1450),
.B(n_1559),
.Y(n_1575)
);

BUFx6f_ASAP7_75t_L g1576 ( 
.A(n_1541),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1547),
.A2(n_1480),
.B1(n_1458),
.B2(n_1530),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1535),
.A2(n_1518),
.B1(n_1525),
.B2(n_1521),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1417),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1499),
.Y(n_1580)
);

OAI21xp33_ASAP7_75t_L g1581 ( 
.A1(n_1540),
.A2(n_1561),
.B(n_1518),
.Y(n_1581)
);

OR2x6_ASAP7_75t_L g1582 ( 
.A(n_1414),
.B(n_1545),
.Y(n_1582)
);

OAI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1501),
.A2(n_1453),
.B(n_1471),
.Y(n_1583)
);

BUFx4f_ASAP7_75t_L g1584 ( 
.A(n_1465),
.Y(n_1584)
);

OAI21xp5_ASAP7_75t_SL g1585 ( 
.A1(n_1420),
.A2(n_1428),
.B(n_1475),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1546),
.A2(n_1476),
.B1(n_1484),
.B2(n_1521),
.Y(n_1586)
);

INVx6_ASAP7_75t_L g1587 ( 
.A(n_1425),
.Y(n_1587)
);

CKINVDCx20_ASAP7_75t_R g1588 ( 
.A(n_1557),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1535),
.A2(n_1521),
.B1(n_1525),
.B2(n_1536),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1525),
.A2(n_1540),
.B1(n_1476),
.B2(n_1537),
.Y(n_1590)
);

BUFx2_ASAP7_75t_R g1591 ( 
.A(n_1464),
.Y(n_1591)
);

BUFx10_ASAP7_75t_L g1592 ( 
.A(n_1429),
.Y(n_1592)
);

BUFx2_ASAP7_75t_R g1593 ( 
.A(n_1555),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1471),
.A2(n_1415),
.B(n_1523),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1499),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1505),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1484),
.A2(n_1517),
.B1(n_1489),
.B2(n_1467),
.Y(n_1597)
);

OAI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1451),
.A2(n_1484),
.B1(n_1533),
.B2(n_1520),
.Y(n_1598)
);

NAND2x1p5_ASAP7_75t_L g1599 ( 
.A(n_1411),
.B(n_1423),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1416),
.Y(n_1600)
);

BUFx12f_ASAP7_75t_L g1601 ( 
.A(n_1438),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1517),
.A2(n_1490),
.B1(n_1522),
.B2(n_1543),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1485),
.B(n_1456),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1451),
.A2(n_1533),
.B1(n_1506),
.B2(n_1447),
.Y(n_1604)
);

CKINVDCx11_ASAP7_75t_R g1605 ( 
.A(n_1439),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1520),
.A2(n_1513),
.B1(n_1549),
.B2(n_1528),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1422),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1504),
.B(n_1410),
.Y(n_1608)
);

OAI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1459),
.A2(n_1440),
.B(n_1432),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1430),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1486),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1435),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_1557),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1415),
.A2(n_1470),
.B(n_1424),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1431),
.Y(n_1615)
);

OAI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1545),
.A2(n_1411),
.B1(n_1423),
.B2(n_1500),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1550),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1434),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1455),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1513),
.A2(n_1538),
.B1(n_1526),
.B2(n_1498),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1469),
.Y(n_1621)
);

NAND2x1p5_ASAP7_75t_L g1622 ( 
.A(n_1411),
.B(n_1423),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1474),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1552),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1483),
.Y(n_1625)
);

BUFx4f_ASAP7_75t_L g1626 ( 
.A(n_1420),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1503),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_SL g1628 ( 
.A1(n_1435),
.A2(n_1560),
.B1(n_1508),
.B2(n_1442),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1553),
.Y(n_1629)
);

INVx6_ASAP7_75t_L g1630 ( 
.A(n_1442),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1514),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1526),
.A2(n_1502),
.B1(n_1544),
.B2(n_1519),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1441),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1539),
.A2(n_1544),
.B1(n_1445),
.B2(n_1435),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_1560),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1524),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1448),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1448),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1446),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1494),
.Y(n_1640)
);

BUFx2_ASAP7_75t_SL g1641 ( 
.A(n_1428),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1510),
.Y(n_1642)
);

BUFx10_ASAP7_75t_L g1643 ( 
.A(n_1429),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1421),
.A2(n_1531),
.B1(n_1461),
.B2(n_1479),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1515),
.B(n_1487),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1527),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_1541),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1441),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1457),
.B(n_1515),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1426),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1509),
.A2(n_1495),
.B1(n_1548),
.B2(n_1488),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1426),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1603),
.B(n_1462),
.Y(n_1653)
);

CKINVDCx8_ASAP7_75t_R g1654 ( 
.A(n_1635),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1633),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1617),
.B(n_1542),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1588),
.Y(n_1657)
);

BUFx8_ASAP7_75t_SL g1658 ( 
.A(n_1584),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1565),
.B(n_1462),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_R g1660 ( 
.A(n_1584),
.B(n_1413),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1600),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1566),
.B(n_1468),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1607),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1605),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1574),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1579),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1608),
.B(n_1468),
.Y(n_1667)
);

NOR2x1_ASAP7_75t_L g1668 ( 
.A(n_1585),
.B(n_1482),
.Y(n_1668)
);

BUFx3_ASAP7_75t_L g1669 ( 
.A(n_1574),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1626),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1610),
.Y(n_1671)
);

NAND2xp33_ASAP7_75t_R g1672 ( 
.A(n_1582),
.B(n_1443),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1565),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_R g1674 ( 
.A(n_1626),
.B(n_1413),
.Y(n_1674)
);

INVx4_ASAP7_75t_L g1675 ( 
.A(n_1574),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1601),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1580),
.B(n_1419),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1595),
.B(n_1479),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_R g1679 ( 
.A(n_1587),
.B(n_1548),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1575),
.B(n_1437),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1586),
.A2(n_1445),
.B1(n_1488),
.B2(n_1460),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1649),
.B(n_1449),
.Y(n_1682)
);

CKINVDCx5p33_ASAP7_75t_R g1683 ( 
.A(n_1587),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1596),
.B(n_1493),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1587),
.Y(n_1685)
);

O2A1O1Ixp33_ASAP7_75t_SL g1686 ( 
.A1(n_1571),
.A2(n_1463),
.B(n_1449),
.C(n_1437),
.Y(n_1686)
);

CKINVDCx20_ASAP7_75t_R g1687 ( 
.A(n_1613),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_R g1688 ( 
.A(n_1613),
.B(n_1556),
.Y(n_1688)
);

O2A1O1Ixp33_ASAP7_75t_SL g1689 ( 
.A1(n_1571),
.A2(n_1463),
.B(n_1436),
.C(n_1466),
.Y(n_1689)
);

CKINVDCx16_ASAP7_75t_R g1690 ( 
.A(n_1628),
.Y(n_1690)
);

NAND2x1p5_ASAP7_75t_L g1691 ( 
.A(n_1576),
.B(n_1491),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1568),
.B(n_1436),
.Y(n_1692)
);

INVx1_ASAP7_75t_SL g1693 ( 
.A(n_1572),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1568),
.B(n_1562),
.Y(n_1694)
);

NAND2xp33_ASAP7_75t_R g1695 ( 
.A(n_1582),
.B(n_1443),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1615),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1599),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1563),
.B(n_1507),
.Y(n_1698)
);

BUFx6f_ASAP7_75t_L g1699 ( 
.A(n_1592),
.Y(n_1699)
);

OAI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1582),
.A2(n_1482),
.B1(n_1511),
.B2(n_1460),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1618),
.Y(n_1701)
);

AND2x4_ASAP7_75t_SL g1702 ( 
.A(n_1592),
.B(n_1473),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_SL g1703 ( 
.A1(n_1573),
.A2(n_1534),
.B1(n_1495),
.B2(n_1512),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1564),
.B(n_1478),
.Y(n_1704)
);

CKINVDCx16_ASAP7_75t_R g1705 ( 
.A(n_1572),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_R g1706 ( 
.A(n_1643),
.B(n_1492),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1602),
.B(n_1534),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1611),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1602),
.B(n_1583),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1573),
.B(n_1491),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_R g1711 ( 
.A(n_1643),
.B(n_1466),
.Y(n_1711)
);

NOR3xp33_ASAP7_75t_SL g1712 ( 
.A(n_1598),
.B(n_1497),
.C(n_1470),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1591),
.Y(n_1713)
);

CKINVDCx16_ASAP7_75t_R g1714 ( 
.A(n_1570),
.Y(n_1714)
);

AO32x2_ASAP7_75t_L g1715 ( 
.A1(n_1634),
.A2(n_1532),
.A3(n_1516),
.B1(n_1554),
.B2(n_1418),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1591),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1645),
.B(n_1444),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1619),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1567),
.B(n_1589),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1581),
.A2(n_1529),
.B1(n_1512),
.B2(n_1461),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1621),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1589),
.B(n_1472),
.Y(n_1722)
);

OAI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1709),
.A2(n_1583),
.B(n_1614),
.Y(n_1723)
);

INVxp67_ASAP7_75t_L g1724 ( 
.A(n_1655),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1705),
.A2(n_1578),
.B1(n_1586),
.B2(n_1577),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1693),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1684),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1655),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1673),
.B(n_1614),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1719),
.B(n_1644),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1659),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1693),
.B(n_1598),
.Y(n_1732)
);

INVx4_ASAP7_75t_L g1733 ( 
.A(n_1699),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1678),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1709),
.B(n_1633),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1694),
.B(n_1594),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1707),
.B(n_1648),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1707),
.B(n_1594),
.Y(n_1738)
);

BUFx3_ASAP7_75t_L g1739 ( 
.A(n_1699),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1661),
.B(n_1569),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1667),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1712),
.B(n_1569),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1653),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1663),
.B(n_1632),
.Y(n_1744)
);

INVx2_ASAP7_75t_SL g1745 ( 
.A(n_1668),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1714),
.B(n_1604),
.Y(n_1746)
);

BUFx3_ASAP7_75t_L g1747 ( 
.A(n_1699),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1671),
.Y(n_1748)
);

NOR2x1_ASAP7_75t_L g1749 ( 
.A(n_1681),
.B(n_1616),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1722),
.A2(n_1578),
.B1(n_1590),
.B2(n_1577),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1696),
.B(n_1632),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1692),
.Y(n_1752)
);

OR2x6_ASAP7_75t_L g1753 ( 
.A(n_1681),
.B(n_1634),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1701),
.B(n_1620),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1718),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1721),
.B(n_1620),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_1662),
.Y(n_1757)
);

CKINVDCx16_ASAP7_75t_R g1758 ( 
.A(n_1679),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1682),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1741),
.B(n_1743),
.Y(n_1760)
);

NAND2x1_ASAP7_75t_SL g1761 ( 
.A(n_1749),
.B(n_1675),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1740),
.B(n_1720),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1748),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1727),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1748),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1746),
.B(n_1665),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1758),
.B(n_1669),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1730),
.B(n_1715),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1731),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1757),
.B(n_1708),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1740),
.B(n_1609),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1758),
.B(n_1690),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1730),
.B(n_1715),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1755),
.Y(n_1774)
);

OAI221xp5_ASAP7_75t_SL g1775 ( 
.A1(n_1750),
.A2(n_1597),
.B1(n_1606),
.B2(n_1700),
.C(n_1717),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1744),
.B(n_1751),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1738),
.B(n_1715),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1738),
.B(n_1703),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1755),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1735),
.B(n_1677),
.Y(n_1780)
);

INVx2_ASAP7_75t_SL g1781 ( 
.A(n_1739),
.Y(n_1781)
);

NAND2x1_ASAP7_75t_SL g1782 ( 
.A(n_1749),
.B(n_1675),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1736),
.B(n_1703),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1781),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1763),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1776),
.B(n_1729),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1769),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1771),
.B(n_1745),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1783),
.B(n_1778),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1783),
.B(n_1729),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1763),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1764),
.Y(n_1792)
);

OAI31xp33_ASAP7_75t_SL g1793 ( 
.A1(n_1772),
.A2(n_1725),
.A3(n_1726),
.B(n_1732),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1760),
.B(n_1752),
.Y(n_1794)
);

INVx3_ASAP7_75t_L g1795 ( 
.A(n_1781),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1765),
.Y(n_1796)
);

OR2x6_ASAP7_75t_L g1797 ( 
.A(n_1761),
.B(n_1753),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1765),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1780),
.B(n_1735),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1774),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1780),
.B(n_1737),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1774),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1768),
.B(n_1756),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1770),
.B(n_1759),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1779),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1779),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1768),
.B(n_1756),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1764),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1787),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1787),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1801),
.Y(n_1811)
);

AOI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1789),
.A2(n_1725),
.B1(n_1742),
.B2(n_1778),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1801),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1789),
.B(n_1773),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1794),
.B(n_1775),
.Y(n_1815)
);

INVx1_ASAP7_75t_SL g1816 ( 
.A(n_1784),
.Y(n_1816)
);

NAND2xp33_ASAP7_75t_L g1817 ( 
.A(n_1795),
.B(n_1660),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1790),
.B(n_1773),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1799),
.B(n_1804),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1790),
.B(n_1762),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1799),
.Y(n_1821)
);

A2O1A1Ixp33_ASAP7_75t_L g1822 ( 
.A1(n_1793),
.A2(n_1767),
.B(n_1782),
.C(n_1761),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1795),
.B(n_1762),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1785),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1791),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1796),
.Y(n_1826)
);

BUFx2_ASAP7_75t_L g1827 ( 
.A(n_1795),
.Y(n_1827)
);

NAND3xp33_ASAP7_75t_L g1828 ( 
.A(n_1798),
.B(n_1742),
.C(n_1712),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1800),
.Y(n_1829)
);

OAI22xp33_ASAP7_75t_SL g1830 ( 
.A1(n_1797),
.A2(n_1753),
.B1(n_1745),
.B2(n_1726),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1792),
.Y(n_1831)
);

NOR3xp33_ASAP7_75t_L g1832 ( 
.A(n_1828),
.B(n_1656),
.C(n_1616),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1810),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_SL g1834 ( 
.A1(n_1830),
.A2(n_1742),
.B1(n_1797),
.B2(n_1788),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1810),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1831),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1815),
.A2(n_1742),
.B1(n_1753),
.B2(n_1797),
.Y(n_1837)
);

XNOR2x1_ASAP7_75t_L g1838 ( 
.A(n_1812),
.B(n_1666),
.Y(n_1838)
);

AOI21xp33_ASAP7_75t_L g1839 ( 
.A1(n_1815),
.A2(n_1766),
.B(n_1745),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1817),
.A2(n_1753),
.B1(n_1687),
.B2(n_1797),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1819),
.Y(n_1841)
);

AO21x1_ASAP7_75t_L g1842 ( 
.A1(n_1817),
.A2(n_1733),
.B(n_1788),
.Y(n_1842)
);

NOR3xp33_ASAP7_75t_L g1843 ( 
.A(n_1822),
.B(n_1646),
.C(n_1636),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1836),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1841),
.B(n_1818),
.Y(n_1845)
);

AOI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1843),
.A2(n_1809),
.B1(n_1816),
.B2(n_1822),
.C(n_1813),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1832),
.A2(n_1823),
.B1(n_1811),
.B2(n_1821),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1833),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1838),
.B(n_1664),
.Y(n_1849)
);

AOI322xp5_ASAP7_75t_L g1850 ( 
.A1(n_1834),
.A2(n_1814),
.A3(n_1786),
.B1(n_1807),
.B2(n_1803),
.C1(n_1820),
.C2(n_1713),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1835),
.Y(n_1851)
);

NAND2x1_ASAP7_75t_L g1852 ( 
.A(n_1840),
.B(n_1827),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1837),
.B(n_1814),
.Y(n_1853)
);

AOI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1839),
.A2(n_1829),
.B1(n_1826),
.B2(n_1825),
.C(n_1824),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1840),
.B(n_1788),
.Y(n_1855)
);

OAI221xp5_ASAP7_75t_SL g1856 ( 
.A1(n_1842),
.A2(n_1597),
.B1(n_1753),
.B2(n_1606),
.C(n_1651),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1841),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1834),
.B(n_1762),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1857),
.B(n_1831),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1848),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1846),
.A2(n_1716),
.B(n_1685),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1846),
.B(n_1683),
.Y(n_1862)
);

AO22x1_ASAP7_75t_L g1863 ( 
.A1(n_1849),
.A2(n_1676),
.B1(n_1733),
.B2(n_1697),
.Y(n_1863)
);

OAI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1850),
.A2(n_1782),
.B(n_1689),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1854),
.B(n_1777),
.Y(n_1865)
);

OAI21xp5_ASAP7_75t_SL g1866 ( 
.A1(n_1850),
.A2(n_1702),
.B(n_1593),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1851),
.B(n_1777),
.Y(n_1867)
);

NAND3xp33_ASAP7_75t_L g1868 ( 
.A(n_1856),
.B(n_1639),
.C(n_1638),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_SL g1869 ( 
.A(n_1855),
.B(n_1593),
.Y(n_1869)
);

NOR2x1_ASAP7_75t_L g1870 ( 
.A(n_1852),
.B(n_1657),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_SL g1871 ( 
.A(n_1870),
.B(n_1858),
.Y(n_1871)
);

NOR3x1_ASAP7_75t_L g1872 ( 
.A(n_1866),
.B(n_1853),
.C(n_1658),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1869),
.A2(n_1862),
.B1(n_1868),
.B2(n_1864),
.Y(n_1873)
);

AOI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1863),
.A2(n_1847),
.B(n_1844),
.Y(n_1874)
);

OAI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1861),
.A2(n_1865),
.B(n_1860),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1859),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1867),
.Y(n_1877)
);

AOI211x1_ASAP7_75t_L g1878 ( 
.A1(n_1862),
.A2(n_1723),
.B(n_1802),
.C(n_1805),
.Y(n_1878)
);

AO22x1_ASAP7_75t_L g1879 ( 
.A1(n_1870),
.A2(n_1670),
.B1(n_1697),
.B2(n_1612),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1866),
.A2(n_1845),
.B(n_1686),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1860),
.Y(n_1881)
);

OAI221xp5_ASAP7_75t_L g1882 ( 
.A1(n_1873),
.A2(n_1654),
.B1(n_1672),
.B2(n_1695),
.C(n_1622),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1878),
.B(n_1806),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1876),
.Y(n_1884)
);

OAI322xp33_ASAP7_75t_L g1885 ( 
.A1(n_1881),
.A2(n_1724),
.A3(n_1642),
.B1(n_1640),
.B2(n_1625),
.C1(n_1623),
.C2(n_1631),
.Y(n_1885)
);

AOI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1871),
.A2(n_1670),
.B(n_1637),
.Y(n_1886)
);

NAND4xp25_ASAP7_75t_L g1887 ( 
.A(n_1872),
.B(n_1674),
.C(n_1733),
.D(n_1497),
.Y(n_1887)
);

AOI221xp5_ASAP7_75t_L g1888 ( 
.A1(n_1875),
.A2(n_1688),
.B1(n_1706),
.B2(n_1680),
.C(n_1723),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1880),
.B(n_1874),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1877),
.B(n_1762),
.Y(n_1890)
);

NOR3x1_ASAP7_75t_L g1891 ( 
.A(n_1879),
.B(n_1711),
.C(n_1728),
.Y(n_1891)
);

AOI222xp33_ASAP7_75t_L g1892 ( 
.A1(n_1875),
.A2(n_1627),
.B1(n_1724),
.B2(n_1728),
.C1(n_1704),
.C2(n_1771),
.Y(n_1892)
);

AOI222xp33_ASAP7_75t_L g1893 ( 
.A1(n_1875),
.A2(n_1771),
.B1(n_1754),
.B2(n_1734),
.C1(n_1630),
.C2(n_1751),
.Y(n_1893)
);

NAND3xp33_ASAP7_75t_L g1894 ( 
.A(n_1889),
.B(n_1491),
.C(n_1496),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_1884),
.Y(n_1895)
);

INVxp33_ASAP7_75t_SL g1896 ( 
.A(n_1888),
.Y(n_1896)
);

NOR4xp25_ASAP7_75t_L g1897 ( 
.A(n_1882),
.B(n_1652),
.C(n_1650),
.D(n_1481),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1890),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1885),
.Y(n_1899)
);

AOI221xp5_ASAP7_75t_L g1900 ( 
.A1(n_1899),
.A2(n_1883),
.B1(n_1886),
.B2(n_1887),
.C(n_1891),
.Y(n_1900)
);

OAI211xp5_ASAP7_75t_SL g1901 ( 
.A1(n_1895),
.A2(n_1893),
.B(n_1892),
.C(n_1630),
.Y(n_1901)
);

OAI31xp33_ASAP7_75t_L g1902 ( 
.A1(n_1896),
.A2(n_1622),
.A3(n_1599),
.B(n_1477),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1898),
.B(n_1808),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1894),
.A2(n_1641),
.B1(n_1733),
.B2(n_1698),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1903),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1904),
.Y(n_1906)
);

OAI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1906),
.A2(n_1900),
.B1(n_1901),
.B2(n_1902),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1905),
.B(n_1897),
.Y(n_1908)
);

HB1xp67_ASAP7_75t_L g1909 ( 
.A(n_1907),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1908),
.B(n_1624),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1909),
.B(n_1629),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_1910),
.Y(n_1912)
);

CKINVDCx20_ASAP7_75t_R g1913 ( 
.A(n_1912),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1913),
.B(n_1911),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1914),
.A2(n_1747),
.B1(n_1739),
.B2(n_1710),
.Y(n_1915)
);

OR2x6_ASAP7_75t_L g1916 ( 
.A(n_1915),
.B(n_1691),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1916),
.A2(n_1739),
.B1(n_1747),
.B2(n_1647),
.Y(n_1917)
);


endmodule