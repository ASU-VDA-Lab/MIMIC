module fake_netlist_5_558_n_1970 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1970);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1970;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_174;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_192;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1928;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_990;
wire n_836;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_86),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_42),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_63),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_63),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_58),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_68),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_47),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_98),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_104),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_164),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_159),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_82),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_94),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_46),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_148),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_2),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_48),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_31),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_91),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_81),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_75),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_13),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_32),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_51),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_95),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_53),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_61),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_158),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_83),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_143),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_33),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_40),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_156),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_31),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_49),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_137),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_116),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_53),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_20),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_9),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_73),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_36),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_141),
.Y(n_228)
);

INVxp33_ASAP7_75t_R g229 ( 
.A(n_17),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_147),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_15),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_46),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_121),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_4),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_10),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_17),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_35),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_28),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_32),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_119),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_85),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_19),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_57),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_96),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_27),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_170),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_69),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_56),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_92),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_146),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_100),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_108),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_117),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_101),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_69),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_49),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_13),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_110),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_162),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_6),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_2),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_88),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_58),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_70),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_87),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_60),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_130),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_134),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_65),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_103),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_71),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_21),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_12),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_93),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_64),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_155),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_136),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_68),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_50),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_56),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_72),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_42),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_66),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_26),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_26),
.Y(n_285)
);

BUFx2_ASAP7_75t_SL g286 ( 
.A(n_45),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_79),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_23),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_27),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_90),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_23),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_61),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_97),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_65),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_80),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_102),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_99),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_37),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_76),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_70),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_25),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_60),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_138),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_118),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_30),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_48),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_52),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_150),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_33),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_145),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_4),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_62),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_19),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_171),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_109),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_160),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_5),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_59),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_16),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_28),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_41),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_140),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_29),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_8),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_3),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_37),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_45),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_8),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_51),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_78),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_127),
.Y(n_331)
);

BUFx5_ASAP7_75t_L g332 ( 
.A(n_47),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_131),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_52),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_57),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_3),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_62),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_10),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_151),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_7),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_113),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_133),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_38),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_40),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_332),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_194),
.B(n_0),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_227),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_173),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_192),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_184),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_332),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_332),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_185),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_R g354 ( 
.A(n_219),
.B(n_122),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_191),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_194),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_212),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_206),
.B(n_0),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_186),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_332),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_332),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_188),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_332),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_240),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_332),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_332),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_198),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_257),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_257),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_257),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_270),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_200),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_202),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_257),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_256),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_211),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_257),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_213),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_257),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_288),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_225),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_241),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_288),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_288),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_183),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_288),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_288),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_288),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_191),
.B(n_1),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_303),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_256),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_216),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_221),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_230),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_231),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_244),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_231),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_206),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_249),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g400 ( 
.A(n_272),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_270),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_231),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_250),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_231),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_251),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_231),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_189),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_189),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_R g409 ( 
.A(n_252),
.B(n_123),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_326),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_326),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_253),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_232),
.B(n_1),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_225),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_254),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_232),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_338),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_338),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_196),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_174),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_174),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_259),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_175),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_175),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_268),
.Y(n_425)
);

NOR2xp67_ASAP7_75t_L g426 ( 
.A(n_236),
.B(n_5),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_178),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_178),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_179),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_176),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_356),
.B(n_274),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_371),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_371),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_395),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_395),
.B(n_274),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_397),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_397),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_347),
.B(n_346),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_349),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_348),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_402),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_350),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_353),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_401),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_404),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_359),
.Y(n_448)
);

AND2x6_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_207),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_362),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_367),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_372),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_404),
.B(n_277),
.Y(n_453)
);

BUFx12f_ASAP7_75t_L g454 ( 
.A(n_373),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_406),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_401),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_376),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_347),
.B(n_225),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_401),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_406),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_368),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_378),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_357),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_345),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_368),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_345),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_358),
.B(n_222),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_369),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_369),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_364),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_370),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_370),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_374),
.Y(n_473)
);

BUFx8_ASAP7_75t_L g474 ( 
.A(n_375),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_R g475 ( 
.A(n_375),
.B(n_181),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_351),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_374),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_377),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_392),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_389),
.B(n_246),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_377),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_R g482 ( 
.A(n_393),
.B(n_296),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_379),
.Y(n_483)
);

NOR2xp67_ASAP7_75t_L g484 ( 
.A(n_351),
.B(n_180),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_379),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_394),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_352),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_396),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_380),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_380),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_403),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_383),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_405),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_383),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_426),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_384),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_355),
.B(n_297),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_384),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_415),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_422),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_426),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_386),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_352),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_382),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_386),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_360),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_413),
.B(n_243),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_440),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_466),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_464),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_464),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_L g512 ( 
.A(n_449),
.B(n_207),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_495),
.B(n_419),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_467),
.B(n_399),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_497),
.B(n_355),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_507),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_464),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_495),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_474),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_464),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_466),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_464),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_507),
.B(n_416),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_472),
.Y(n_524)
);

INVx6_ASAP7_75t_L g525 ( 
.A(n_466),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_497),
.B(n_387),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_480),
.B(n_453),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_480),
.B(n_207),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_467),
.B(n_412),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_476),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_472),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_466),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_476),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_507),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_476),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_453),
.B(n_387),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_435),
.B(n_177),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_476),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_466),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_431),
.B(n_388),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_476),
.Y(n_541)
);

INVx6_ASAP7_75t_L g542 ( 
.A(n_466),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_431),
.B(n_425),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_503),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_474),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_503),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_458),
.B(n_381),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_474),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_503),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_501),
.B(n_388),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_466),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_503),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_501),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_503),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_458),
.B(n_381),
.Y(n_555)
);

AND2x2_ASAP7_75t_SL g556 ( 
.A(n_436),
.B(n_389),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_461),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_487),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_SL g559 ( 
.A(n_475),
.B(n_400),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_461),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_472),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_487),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_487),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_487),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_435),
.B(n_398),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_463),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_441),
.B(n_443),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_487),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_470),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_449),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_465),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_449),
.B(n_385),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_449),
.B(n_360),
.Y(n_573)
);

BUFx4f_ASAP7_75t_L g574 ( 
.A(n_487),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_504),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_437),
.B(n_407),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_439),
.A2(n_414),
.B1(n_430),
.B2(n_391),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_482),
.B(n_414),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_449),
.A2(n_245),
.B1(n_236),
.B2(n_243),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_449),
.B(n_361),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_437),
.B(n_407),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_465),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_468),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_487),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_449),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_439),
.A2(n_328),
.B1(n_203),
.B2(n_204),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_506),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_449),
.B(n_361),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_506),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_475),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_482),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_449),
.B(n_363),
.Y(n_592)
);

OR2x6_ASAP7_75t_L g593 ( 
.A(n_454),
.B(n_286),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_506),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_468),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_506),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_438),
.B(n_177),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_444),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_448),
.B(n_419),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_506),
.B(n_363),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_506),
.B(n_365),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_469),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_506),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_469),
.B(n_365),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_438),
.B(n_408),
.Y(n_605)
);

INVxp33_ASAP7_75t_L g606 ( 
.A(n_436),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_471),
.B(n_366),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_471),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_473),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_433),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_474),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_433),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_450),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_473),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_451),
.B(n_390),
.Y(n_615)
);

INVx6_ASAP7_75t_L g616 ( 
.A(n_433),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_484),
.A2(n_245),
.B1(n_279),
.B2(n_199),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_474),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_477),
.Y(n_619)
);

INVxp67_ASAP7_75t_SL g620 ( 
.A(n_484),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_454),
.B(n_286),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_433),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_452),
.B(n_354),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_477),
.Y(n_624)
);

INVx5_ASAP7_75t_L g625 ( 
.A(n_433),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_478),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_433),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_433),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_454),
.B(n_457),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_481),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_442),
.B(n_408),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_481),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_445),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_485),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_445),
.Y(n_635)
);

NAND2x1p5_ASAP7_75t_L g636 ( 
.A(n_485),
.B(n_182),
.Y(n_636)
);

OR2x6_ASAP7_75t_L g637 ( 
.A(n_442),
.B(n_279),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_462),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_489),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_489),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_494),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_479),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_494),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_486),
.B(n_409),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_445),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_446),
.B(n_182),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_446),
.B(n_179),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_478),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_447),
.B(n_187),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_502),
.B(n_366),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_478),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_488),
.B(n_222),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_491),
.B(n_222),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_445),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_493),
.B(n_322),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_445),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_499),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_502),
.Y(n_658)
);

INVxp33_ASAP7_75t_L g659 ( 
.A(n_447),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_483),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_515),
.B(n_527),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_569),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_516),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_556),
.B(n_526),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_606),
.B(n_500),
.Y(n_665)
);

BUFx5_ASAP7_75t_L g666 ( 
.A(n_510),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_556),
.B(n_540),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_509),
.A2(n_434),
.B(n_432),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_536),
.B(n_455),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_634),
.B(n_455),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_553),
.B(n_225),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_634),
.B(n_460),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_524),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_524),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_570),
.B(n_207),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_531),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_620),
.B(n_460),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_553),
.B(n_518),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_523),
.B(n_187),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_570),
.B(n_207),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_R g681 ( 
.A(n_591),
.B(n_299),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_590),
.B(n_239),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_523),
.B(n_193),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_516),
.B(n_193),
.Y(n_684)
);

NOR2x2_ASAP7_75t_L g685 ( 
.A(n_593),
.B(n_229),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_514),
.A2(n_330),
.B1(n_339),
.B2(n_315),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_534),
.B(n_557),
.Y(n_687)
);

O2A1O1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_550),
.A2(n_318),
.B(n_261),
.C(n_238),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_591),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_534),
.Y(n_690)
);

NAND3xp33_ASAP7_75t_L g691 ( 
.A(n_529),
.B(n_205),
.C(n_197),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_531),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_561),
.Y(n_693)
);

AND3x1_ASAP7_75t_L g694 ( 
.A(n_577),
.B(n_229),
.C(n_224),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_561),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_513),
.Y(n_696)
);

OR2x6_ASAP7_75t_L g697 ( 
.A(n_611),
.B(n_519),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_557),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_576),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_576),
.Y(n_700)
);

AO22x1_ASAP7_75t_L g701 ( 
.A1(n_586),
.A2(n_261),
.B1(n_280),
.B2(n_278),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_SL g702 ( 
.A(n_598),
.B(n_234),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_560),
.B(n_195),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_559),
.A2(n_304),
.B1(n_314),
.B2(n_308),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_513),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_560),
.B(n_571),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_581),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_571),
.B(n_195),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_528),
.A2(n_280),
.B1(n_285),
.B2(n_294),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_626),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_655),
.B(n_208),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_582),
.B(n_209),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_567),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_508),
.B(n_420),
.Y(n_714)
);

NAND3xp33_ASAP7_75t_SL g715 ( 
.A(n_547),
.B(n_269),
.C(n_242),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_626),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_659),
.B(n_210),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_528),
.A2(n_238),
.B1(n_327),
.B2(n_294),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_581),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_566),
.B(n_575),
.Y(n_720)
);

O2A1O1Ixp5_ASAP7_75t_L g721 ( 
.A1(n_510),
.A2(n_262),
.B(n_201),
.C(n_190),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_582),
.B(n_209),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_605),
.Y(n_723)
);

NAND2x1_ASAP7_75t_L g724 ( 
.A(n_616),
.B(n_456),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_583),
.B(n_220),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_528),
.A2(n_327),
.B1(n_278),
.B2(n_263),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_535),
.Y(n_727)
);

AND2x6_ASAP7_75t_L g728 ( 
.A(n_511),
.B(n_220),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_583),
.B(n_228),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_565),
.B(n_214),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_L g731 ( 
.A(n_599),
.B(n_74),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_595),
.B(n_228),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_595),
.B(n_233),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_638),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_565),
.B(n_215),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_638),
.Y(n_736)
);

AOI22x1_ASAP7_75t_L g737 ( 
.A1(n_511),
.A2(n_262),
.B1(n_258),
.B2(n_293),
.Y(n_737)
);

INVx8_ASAP7_75t_L g738 ( 
.A(n_593),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_602),
.B(n_608),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_537),
.B(n_420),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_602),
.B(n_233),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_611),
.B(n_199),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_572),
.B(n_217),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_568),
.A2(n_490),
.B(n_483),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_608),
.B(n_287),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_543),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_609),
.B(n_287),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_570),
.B(n_207),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_648),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_605),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_631),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_631),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_609),
.Y(n_753)
);

NAND3xp33_ASAP7_75t_L g754 ( 
.A(n_555),
.B(n_617),
.C(n_623),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_614),
.B(n_295),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_614),
.B(n_295),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_648),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_619),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_578),
.A2(n_333),
.B1(n_310),
.B2(n_342),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_535),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_619),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_652),
.B(n_218),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_624),
.B(n_310),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_544),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_624),
.B(n_316),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_537),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_630),
.B(n_316),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_630),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_537),
.B(n_597),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_570),
.B(n_270),
.Y(n_770)
);

AND2x2_ASAP7_75t_SL g771 ( 
.A(n_512),
.B(n_180),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_570),
.B(n_270),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_570),
.B(n_270),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_632),
.Y(n_774)
);

INVx8_ASAP7_75t_L g775 ( 
.A(n_593),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_613),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_653),
.B(n_223),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_632),
.B(n_331),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_651),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_528),
.A2(n_331),
.B1(n_333),
.B2(n_342),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_544),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_519),
.B(n_224),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_647),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_585),
.B(n_290),
.Y(n_784)
);

INVx5_ASAP7_75t_L g785 ( 
.A(n_532),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_615),
.Y(n_786)
);

AND2x6_ASAP7_75t_SL g787 ( 
.A(n_593),
.B(n_248),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_639),
.Y(n_788)
);

NOR3xp33_ASAP7_75t_SL g789 ( 
.A(n_644),
.B(n_235),
.C(n_226),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_585),
.B(n_290),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_597),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_639),
.B(n_237),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_647),
.B(n_421),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_640),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_585),
.B(n_290),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_640),
.B(n_341),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_641),
.B(n_247),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_641),
.B(n_341),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_585),
.B(n_290),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_647),
.B(n_421),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_585),
.B(n_290),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_643),
.B(n_255),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_647),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_643),
.B(n_190),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_528),
.A2(n_646),
.B1(n_649),
.B2(n_597),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_646),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_658),
.B(n_260),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_528),
.A2(n_201),
.B1(n_258),
.B2(n_276),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_658),
.B(n_276),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_627),
.A2(n_505),
.B(n_498),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_642),
.B(n_239),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_SL g812 ( 
.A(n_545),
.B(n_271),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_528),
.A2(n_312),
.B1(n_318),
.B2(n_317),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_SL g814 ( 
.A(n_629),
.B(n_300),
.C(n_264),
.Y(n_814)
);

AND2x6_ASAP7_75t_L g815 ( 
.A(n_517),
.B(n_293),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_520),
.B(n_505),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_637),
.A2(n_222),
.B1(n_265),
.B2(n_267),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_573),
.B(n_445),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_520),
.B(n_483),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_522),
.B(n_505),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_646),
.B(n_649),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_651),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_649),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_522),
.B(n_490),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_530),
.Y(n_825)
);

NOR2x2_ASAP7_75t_L g826 ( 
.A(n_621),
.B(n_239),
.Y(n_826)
);

INVx4_ASAP7_75t_L g827 ( 
.A(n_532),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_580),
.B(n_445),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_579),
.A2(n_248),
.B1(n_263),
.B2(n_285),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_530),
.B(n_490),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_588),
.B(n_459),
.Y(n_831)
);

INVx5_ASAP7_75t_L g832 ( 
.A(n_728),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_713),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_714),
.Y(n_834)
);

BUFx4f_ASAP7_75t_L g835 ( 
.A(n_738),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_663),
.B(n_637),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_664),
.B(n_592),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_769),
.B(n_545),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_661),
.B(n_533),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_727),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_705),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_661),
.B(n_533),
.Y(n_842)
);

NOR3xp33_ASAP7_75t_SL g843 ( 
.A(n_715),
.B(n_273),
.C(n_266),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_690),
.B(n_769),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_662),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_821),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_821),
.B(n_699),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_698),
.Y(n_848)
);

NOR2x1p5_ASAP7_75t_L g849 ( 
.A(n_814),
.B(n_548),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_667),
.B(n_538),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_682),
.B(n_696),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_805),
.B(n_538),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_689),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_711),
.B(n_541),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_776),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_698),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_R g857 ( 
.A(n_734),
.B(n_548),
.Y(n_857)
);

OAI21xp33_ASAP7_75t_L g858 ( 
.A1(n_711),
.A2(n_621),
.B(n_637),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_709),
.A2(n_512),
.B1(n_311),
.B2(n_312),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_700),
.B(n_707),
.Y(n_860)
);

BUFx4f_ASAP7_75t_L g861 ( 
.A(n_738),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_687),
.B(n_541),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_753),
.B(n_546),
.Y(n_863)
);

NOR3xp33_ASAP7_75t_SL g864 ( 
.A(n_812),
.B(n_281),
.C(n_275),
.Y(n_864)
);

OR2x2_ASAP7_75t_SL g865 ( 
.A(n_691),
.B(n_657),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_727),
.Y(n_866)
);

INVx3_ASAP7_75t_SL g867 ( 
.A(n_736),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_766),
.B(n_618),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_758),
.B(n_546),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_825),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_761),
.B(n_549),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_783),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_768),
.B(n_549),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_673),
.Y(n_874)
);

CKINVDCx11_ASAP7_75t_R g875 ( 
.A(n_787),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_774),
.B(n_552),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_788),
.B(n_552),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_746),
.B(n_621),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_805),
.B(n_554),
.Y(n_879)
);

INVxp67_ASAP7_75t_SL g880 ( 
.A(n_760),
.Y(n_880)
);

INVx1_ASAP7_75t_SL g881 ( 
.A(n_720),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_731),
.B(n_554),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_674),
.Y(n_883)
);

AO22x1_ASAP7_75t_L g884 ( 
.A1(n_762),
.A2(n_618),
.B1(n_283),
.B2(n_337),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_783),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_794),
.B(n_600),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_666),
.B(n_539),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_676),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_692),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_665),
.B(n_621),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_806),
.A2(n_637),
.B1(n_587),
.B2(n_558),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_760),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_719),
.B(n_423),
.Y(n_893)
);

BUFx12f_ASAP7_75t_SL g894 ( 
.A(n_782),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_693),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_803),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_665),
.B(n_539),
.Y(n_897)
);

BUFx8_ASAP7_75t_SL g898 ( 
.A(n_811),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_723),
.B(n_423),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_695),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_806),
.A2(n_558),
.B1(n_587),
.B2(n_563),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_743),
.B(n_601),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_750),
.B(n_424),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_738),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_751),
.B(n_424),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_764),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_743),
.B(n_539),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_752),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_730),
.B(n_563),
.Y(n_909)
);

NAND2xp33_ASAP7_75t_R g910 ( 
.A(n_789),
.B(n_282),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_710),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_791),
.B(n_427),
.Y(n_912)
);

INVx2_ASAP7_75t_SL g913 ( 
.A(n_671),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_764),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_775),
.Y(n_915)
);

AOI21x1_ASAP7_75t_L g916 ( 
.A1(n_818),
.A2(n_607),
.B(n_604),
.Y(n_916)
);

AND2x6_ASAP7_75t_L g917 ( 
.A(n_808),
.B(n_563),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_681),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_706),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_775),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_730),
.B(n_735),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_786),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_666),
.B(n_584),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_823),
.B(n_427),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_803),
.Y(n_925)
);

NAND3xp33_ASAP7_75t_SL g926 ( 
.A(n_702),
.B(n_298),
.C(n_284),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_735),
.B(n_239),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_739),
.B(n_584),
.Y(n_928)
);

AOI22x1_ASAP7_75t_L g929 ( 
.A1(n_781),
.A2(n_716),
.B1(n_757),
.B2(n_749),
.Y(n_929)
);

BUFx10_ASAP7_75t_L g930 ( 
.A(n_762),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_666),
.B(n_584),
.Y(n_931)
);

INVx5_ASAP7_75t_L g932 ( 
.A(n_728),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_670),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_672),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_779),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_793),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_740),
.B(n_428),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_679),
.B(n_594),
.Y(n_938)
);

INVx1_ASAP7_75t_SL g939 ( 
.A(n_681),
.Y(n_939)
);

BUFx4f_ASAP7_75t_L g940 ( 
.A(n_775),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_822),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_683),
.B(n_594),
.Y(n_942)
);

BUFx4f_ASAP7_75t_L g943 ( 
.A(n_697),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_666),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_781),
.Y(n_945)
);

NAND3xp33_ASAP7_75t_SL g946 ( 
.A(n_777),
.B(n_686),
.C(n_759),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_800),
.B(n_636),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_704),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_740),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_669),
.B(n_594),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_684),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_R g952 ( 
.A(n_678),
.B(n_289),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_754),
.B(n_428),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_742),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_785),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_677),
.Y(n_956)
);

OR2x6_ASAP7_75t_L g957 ( 
.A(n_697),
.B(n_636),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_792),
.B(n_603),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_816),
.Y(n_959)
);

INVx4_ASAP7_75t_SL g960 ( 
.A(n_728),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_819),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_792),
.B(n_603),
.Y(n_962)
);

NOR2xp67_ASAP7_75t_L g963 ( 
.A(n_717),
.B(n_777),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_742),
.B(n_429),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_724),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_678),
.A2(n_603),
.B1(n_525),
.B2(n_542),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_797),
.B(n_636),
.Y(n_967)
);

CKINVDCx8_ASAP7_75t_R g968 ( 
.A(n_782),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_666),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_717),
.B(n_650),
.Y(n_970)
);

OR2x6_ASAP7_75t_L g971 ( 
.A(n_697),
.B(n_782),
.Y(n_971)
);

AND3x2_ASAP7_75t_SL g972 ( 
.A(n_694),
.B(n_302),
.C(n_265),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_742),
.B(n_429),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_820),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_827),
.Y(n_975)
);

NOR3xp33_ASAP7_75t_SL g976 ( 
.A(n_797),
.B(n_291),
.C(n_292),
.Y(n_976)
);

NAND2xp33_ASAP7_75t_R g977 ( 
.A(n_802),
.B(n_807),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_824),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_802),
.B(n_302),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_807),
.B(n_521),
.Y(n_980)
);

NOR3xp33_ASAP7_75t_SL g981 ( 
.A(n_688),
.B(n_323),
.C(n_305),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_830),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_703),
.B(n_311),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_685),
.Y(n_984)
);

NAND2xp33_ASAP7_75t_SL g985 ( 
.A(n_708),
.B(n_712),
.Y(n_985)
);

CKINVDCx11_ASAP7_75t_R g986 ( 
.A(n_826),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_771),
.B(n_610),
.Y(n_987)
);

BUFx12f_ASAP7_75t_L g988 ( 
.A(n_728),
.Y(n_988)
);

OR2x2_ASAP7_75t_SL g989 ( 
.A(n_817),
.B(n_317),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_722),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_827),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_771),
.B(n_610),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_701),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_666),
.B(n_610),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_725),
.B(n_628),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_728),
.A2(n_741),
.B1(n_733),
.B2(n_745),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_815),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_804),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_729),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_732),
.Y(n_1000)
);

AND2x6_ASAP7_75t_L g1001 ( 
.A(n_780),
.B(n_532),
.Y(n_1001)
);

NOR2x1_ASAP7_75t_L g1002 ( 
.A(n_747),
.B(n_521),
.Y(n_1002)
);

AO22x1_ASAP7_75t_L g1003 ( 
.A1(n_815),
.A2(n_335),
.B1(n_301),
.B2(n_321),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_755),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_756),
.B(n_763),
.Y(n_1005)
);

AND3x1_ASAP7_75t_L g1006 ( 
.A(n_829),
.B(n_344),
.C(n_418),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_785),
.Y(n_1007)
);

INVx5_ASAP7_75t_L g1008 ( 
.A(n_815),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_765),
.B(n_302),
.Y(n_1009)
);

BUFx4_ASAP7_75t_SL g1010 ( 
.A(n_829),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_767),
.B(n_628),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_785),
.B(n_532),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_778),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_815),
.Y(n_1014)
);

NOR3xp33_ASAP7_75t_SL g1015 ( 
.A(n_796),
.B(n_325),
.C(n_336),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_798),
.B(n_628),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_809),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_818),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_815),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_828),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_828),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_709),
.B(n_633),
.Y(n_1022)
);

OAI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_718),
.A2(n_344),
.B1(n_319),
.B2(n_320),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_902),
.A2(n_574),
.B(n_785),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_921),
.A2(n_831),
.B(n_668),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_956),
.B(n_718),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_967),
.A2(n_831),
.B(n_810),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_919),
.B(n_726),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_907),
.A2(n_574),
.B(n_980),
.Y(n_1029)
);

NAND2x1_ASAP7_75t_L g1030 ( 
.A(n_975),
.B(n_525),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_980),
.A2(n_574),
.B(n_564),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_970),
.B(n_726),
.Y(n_1032)
);

CKINVDCx16_ASAP7_75t_R g1033 ( 
.A(n_855),
.Y(n_1033)
);

NOR2xp67_ASAP7_75t_L g1034 ( 
.A(n_833),
.B(n_813),
.Y(n_1034)
);

OAI21x1_ASAP7_75t_L g1035 ( 
.A1(n_929),
.A2(n_721),
.B(n_737),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_975),
.A2(n_521),
.B(n_564),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_837),
.A2(n_744),
.B(n_680),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_991),
.A2(n_564),
.B(n_654),
.Y(n_1038)
);

AO31x2_ASAP7_75t_L g1039 ( 
.A1(n_970),
.A2(n_660),
.A3(n_654),
.B(n_645),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_846),
.B(n_770),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_963),
.B(n_813),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_933),
.B(n_633),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_846),
.B(n_770),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_936),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_916),
.A2(n_633),
.B(n_799),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_848),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_994),
.A2(n_801),
.B(n_799),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_934),
.B(n_660),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_850),
.A2(n_801),
.B(n_795),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_854),
.A2(n_947),
.B1(n_999),
.B2(n_951),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1000),
.B(n_772),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1000),
.B(n_772),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1013),
.B(n_773),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_837),
.A2(n_748),
.B(n_675),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_850),
.A2(n_795),
.B(n_790),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_839),
.A2(n_790),
.B(n_784),
.Y(n_1056)
);

AO31x2_ASAP7_75t_L g1057 ( 
.A1(n_909),
.A2(n_654),
.A3(n_645),
.B(n_498),
.Y(n_1057)
);

NAND2xp33_ASAP7_75t_L g1058 ( 
.A(n_832),
.B(n_532),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_977),
.A2(n_946),
.B1(n_890),
.B2(n_948),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_897),
.A2(n_773),
.B1(n_784),
.B2(n_748),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_979),
.A2(n_313),
.B(n_340),
.C(n_306),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_987),
.A2(n_680),
.B(n_675),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1013),
.B(n_525),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_881),
.B(n_410),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_990),
.A2(n_324),
.B(n_329),
.C(n_307),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1004),
.B(n_953),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_991),
.A2(n_645),
.B(n_551),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_842),
.A2(n_434),
.B(n_432),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_887),
.A2(n_931),
.B(n_923),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_953),
.B(n_959),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_856),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_961),
.B(n_974),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_851),
.B(n_302),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_944),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_SL g1075 ( 
.A1(n_944),
.A2(n_492),
.B(n_498),
.Y(n_1075)
);

AO31x2_ASAP7_75t_L g1076 ( 
.A1(n_897),
.A2(n_496),
.A3(n_492),
.B(n_434),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_978),
.B(n_525),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_887),
.A2(n_432),
.B(n_496),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_982),
.B(n_542),
.Y(n_1079)
);

OAI22x1_ASAP7_75t_L g1080 ( 
.A1(n_890),
.A2(n_309),
.B1(n_334),
.B2(n_343),
.Y(n_1080)
);

AOI21xp33_ASAP7_75t_L g1081 ( 
.A1(n_977),
.A2(n_927),
.B(n_834),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_860),
.B(n_542),
.Y(n_1082)
);

AND2x2_ASAP7_75t_SL g1083 ( 
.A(n_943),
.B(n_859),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_860),
.B(n_1017),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_992),
.A2(n_496),
.B(n_492),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_923),
.A2(n_456),
.B(n_411),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_870),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_931),
.A2(n_456),
.B(n_411),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_938),
.A2(n_562),
.B(n_551),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_942),
.A2(n_562),
.B(n_551),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_870),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_912),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_882),
.A2(n_456),
.B(n_417),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_969),
.Y(n_1094)
);

BUFx12f_ASAP7_75t_L g1095 ( 
.A(n_845),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_874),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_955),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1005),
.B(n_542),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_882),
.A2(n_410),
.B(n_417),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_852),
.A2(n_596),
.B(n_625),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_852),
.A2(n_596),
.B(n_625),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_859),
.A2(n_265),
.B1(n_267),
.B2(n_418),
.Y(n_1102)
);

NAND2x1p5_ASAP7_75t_L g1103 ( 
.A(n_832),
.B(n_551),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_874),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_969),
.A2(n_1011),
.B(n_995),
.Y(n_1105)
);

AO21x2_ASAP7_75t_L g1106 ( 
.A1(n_958),
.A2(n_589),
.B(n_551),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1016),
.A2(n_562),
.B(n_589),
.Y(n_1107)
);

NOR2xp67_ASAP7_75t_L g1108 ( 
.A(n_913),
.B(n_77),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_950),
.A2(n_962),
.B(n_928),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_1005),
.B(n_562),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1018),
.A2(n_1021),
.B(n_869),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_998),
.A2(n_616),
.A3(n_7),
.B(n_9),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_936),
.B(n_265),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1005),
.B(n_562),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_863),
.A2(n_589),
.B(n_616),
.Y(n_1115)
);

AO31x2_ASAP7_75t_L g1116 ( 
.A1(n_998),
.A2(n_862),
.A3(n_1022),
.B(n_876),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1023),
.A2(n_267),
.B1(n_616),
.B2(n_589),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_858),
.A2(n_589),
.B(n_635),
.C(n_612),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_912),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_908),
.B(n_656),
.Y(n_1120)
);

OAI22x1_ASAP7_75t_L g1121 ( 
.A1(n_954),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_955),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_983),
.B(n_656),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1009),
.B(n_267),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_879),
.A2(n_656),
.B1(n_635),
.B2(n_612),
.Y(n_1125)
);

AOI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1020),
.A2(n_656),
.B(n_635),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_871),
.A2(n_596),
.B(n_635),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_983),
.B(n_656),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_924),
.B(n_635),
.Y(n_1129)
);

AO21x2_ASAP7_75t_L g1130 ( 
.A1(n_996),
.A2(n_612),
.B(n_596),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_855),
.Y(n_1131)
);

NOR2xp67_ASAP7_75t_L g1132 ( 
.A(n_918),
.B(n_169),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_924),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_846),
.B(n_128),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_879),
.A2(n_596),
.B(n_622),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_873),
.A2(n_11),
.A3(n_14),
.B(n_15),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1020),
.A2(n_596),
.B(n_622),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_SL g1138 ( 
.A1(n_891),
.A2(n_167),
.B(n_153),
.Y(n_1138)
);

O2A1O1Ixp5_ASAP7_75t_L g1139 ( 
.A1(n_985),
.A2(n_612),
.B(n_152),
.C(n_149),
.Y(n_1139)
);

NOR2x1_ASAP7_75t_R g1140 ( 
.A(n_875),
.B(n_459),
.Y(n_1140)
);

AOI21x1_ASAP7_75t_L g1141 ( 
.A1(n_877),
.A2(n_612),
.B(n_622),
.Y(n_1141)
);

INVx4_ASAP7_75t_L g1142 ( 
.A(n_846),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_893),
.B(n_899),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1014),
.A2(n_625),
.B(n_622),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1014),
.A2(n_625),
.B(n_622),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1002),
.A2(n_625),
.B(n_622),
.Y(n_1146)
);

NOR2xp67_ASAP7_75t_L g1147 ( 
.A(n_878),
.B(n_139),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_886),
.A2(n_985),
.B(n_1008),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_883),
.Y(n_1149)
);

AOI22x1_ASAP7_75t_L g1150 ( 
.A1(n_883),
.A2(n_459),
.B1(n_114),
.B2(n_135),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_901),
.A2(n_625),
.B(n_459),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1012),
.A2(n_111),
.B(n_132),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1008),
.A2(n_459),
.B(n_126),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_904),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_888),
.A2(n_459),
.B(n_124),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_893),
.B(n_459),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_899),
.B(n_14),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1012),
.A2(n_120),
.B(n_112),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1023),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_840),
.A2(n_107),
.B(n_106),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_903),
.B(n_18),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_888),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_993),
.A2(n_21),
.B(n_22),
.C(n_24),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_889),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1008),
.A2(n_105),
.B(n_89),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_840),
.A2(n_914),
.B(n_906),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_889),
.A2(n_84),
.B(n_24),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_903),
.B(n_22),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_867),
.B(n_25),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_880),
.A2(n_957),
.B1(n_914),
.B2(n_906),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_895),
.A2(n_29),
.B(n_30),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_895),
.A2(n_34),
.B(n_35),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_945),
.A2(n_34),
.B(n_36),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_922),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_900),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_922),
.B(n_38),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_900),
.A2(n_39),
.B(n_41),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_878),
.A2(n_39),
.B(n_43),
.C(n_44),
.Y(n_1178)
);

NOR2x1_ASAP7_75t_SL g1179 ( 
.A(n_832),
.B(n_43),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_843),
.A2(n_44),
.B(n_50),
.C(n_54),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_911),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_911),
.A2(n_54),
.B(n_55),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_941),
.A2(n_55),
.B(n_59),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_941),
.A2(n_64),
.B(n_66),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1032),
.A2(n_966),
.B(n_935),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1096),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1095),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_1097),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1134),
.B(n_1142),
.Y(n_1189)
);

OR2x6_ASAP7_75t_L g1190 ( 
.A(n_1134),
.B(n_904),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1127),
.A2(n_965),
.B(n_849),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1058),
.A2(n_1008),
.B(n_932),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1072),
.B(n_1050),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_1131),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1095),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1058),
.A2(n_932),
.B(n_832),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_1134),
.B(n_847),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1096),
.Y(n_1198)
);

AO21x2_ASAP7_75t_L g1199 ( 
.A1(n_1029),
.A2(n_1118),
.B(n_1137),
.Y(n_1199)
);

BUFx8_ASAP7_75t_L g1200 ( 
.A(n_1174),
.Y(n_1200)
);

OA21x2_ASAP7_75t_L g1201 ( 
.A1(n_1105),
.A2(n_981),
.B(n_976),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1131),
.Y(n_1202)
);

OAI221xp5_ASAP7_75t_L g1203 ( 
.A1(n_1059),
.A2(n_843),
.B1(n_926),
.B2(n_976),
.C(n_910),
.Y(n_1203)
);

AOI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1141),
.A2(n_957),
.B(n_905),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1104),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1159),
.A2(n_864),
.B(n_943),
.C(n_905),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1070),
.A2(n_957),
.B1(n_940),
.B2(n_861),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1104),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1097),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_SL g1210 ( 
.A1(n_1179),
.A2(n_949),
.B(n_865),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1127),
.A2(n_1107),
.B(n_1115),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1097),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_1154),
.Y(n_1213)
);

BUFx10_ASAP7_75t_L g1214 ( 
.A(n_1040),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1074),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1073),
.B(n_937),
.Y(n_1216)
);

NOR2x1_ASAP7_75t_R g1217 ( 
.A(n_1154),
.B(n_853),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1118),
.A2(n_885),
.A3(n_896),
.B(n_925),
.Y(n_1218)
);

OR2x6_ASAP7_75t_L g1219 ( 
.A(n_1142),
.B(n_920),
.Y(n_1219)
);

OA21x2_ASAP7_75t_L g1220 ( 
.A1(n_1105),
.A2(n_981),
.B(n_1015),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1159),
.A2(n_864),
.B(n_973),
.C(n_964),
.Y(n_1221)
);

AOI22x1_ASAP7_75t_L g1222 ( 
.A1(n_1080),
.A2(n_1019),
.B1(n_866),
.B2(n_892),
.Y(n_1222)
);

OA21x2_ASAP7_75t_L g1223 ( 
.A1(n_1068),
.A2(n_1015),
.B(n_964),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1109),
.A2(n_932),
.B(n_1007),
.Y(n_1224)
);

NAND3xp33_ASAP7_75t_L g1225 ( 
.A(n_1061),
.B(n_884),
.C(n_910),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1107),
.A2(n_965),
.B(n_1006),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1066),
.B(n_867),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_SL g1228 ( 
.A1(n_1178),
.A2(n_872),
.B(n_972),
.C(n_841),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1031),
.A2(n_932),
.B(n_1007),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1115),
.A2(n_872),
.B(n_917),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1084),
.B(n_853),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1044),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1097),
.Y(n_1233)
);

OR2x6_ASAP7_75t_L g1234 ( 
.A(n_1142),
.B(n_920),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1083),
.A2(n_1026),
.B1(n_1028),
.B2(n_1034),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1087),
.Y(n_1236)
);

OA21x2_ASAP7_75t_L g1237 ( 
.A1(n_1068),
.A2(n_973),
.B(n_937),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1045),
.A2(n_917),
.B(n_960),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1182),
.A2(n_847),
.B(n_1010),
.C(n_997),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1091),
.Y(n_1240)
);

INVx1_ASAP7_75t_SL g1241 ( 
.A(n_1064),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1046),
.Y(n_1242)
);

AO32x2_ASAP7_75t_L g1243 ( 
.A1(n_1170),
.A2(n_972),
.A3(n_989),
.B1(n_930),
.B2(n_971),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1045),
.A2(n_1166),
.B(n_1126),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1166),
.A2(n_917),
.B(n_960),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1071),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1149),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1162),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1081),
.B(n_939),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1111),
.A2(n_917),
.B(n_960),
.Y(n_1250)
);

AO21x2_ASAP7_75t_L g1251 ( 
.A1(n_1155),
.A2(n_952),
.B(n_868),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1111),
.A2(n_917),
.B(n_841),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1035),
.A2(n_1001),
.B(n_988),
.Y(n_1253)
);

NAND3xp33_ASAP7_75t_L g1254 ( 
.A(n_1061),
.B(n_1003),
.C(n_844),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1092),
.B(n_930),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1035),
.A2(n_1001),
.B(n_988),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1122),
.Y(n_1257)
);

BUFx4_ASAP7_75t_SL g1258 ( 
.A(n_1169),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1143),
.B(n_1033),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1164),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1119),
.B(n_915),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1175),
.Y(n_1262)
);

OAI22xp5_ASAP7_75t_L g1263 ( 
.A1(n_1083),
.A2(n_861),
.B1(n_940),
.B2(n_835),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1167),
.A2(n_997),
.B(n_868),
.C(n_835),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1074),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1181),
.Y(n_1266)
);

AO21x2_ASAP7_75t_L g1267 ( 
.A1(n_1130),
.A2(n_952),
.B(n_868),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1178),
.A2(n_1163),
.B(n_1025),
.C(n_1180),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1041),
.A2(n_844),
.B(n_1001),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1133),
.B(n_898),
.Y(n_1270)
);

INVx4_ASAP7_75t_SL g1271 ( 
.A(n_1122),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_SL g1272 ( 
.A1(n_1138),
.A2(n_971),
.B(n_1001),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1099),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1080),
.A2(n_971),
.B1(n_836),
.B2(n_838),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1099),
.Y(n_1275)
);

BUFx8_ASAP7_75t_L g1276 ( 
.A(n_1122),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_1176),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1124),
.B(n_836),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1048),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1120),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1063),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1113),
.Y(n_1282)
);

AO32x2_ASAP7_75t_L g1283 ( 
.A1(n_1060),
.A2(n_1001),
.A3(n_894),
.B1(n_968),
.B2(n_892),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1074),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1157),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1176),
.B(n_984),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1121),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1040),
.B(n_915),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1069),
.A2(n_892),
.B(n_866),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1094),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1094),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1086),
.Y(n_1292)
);

AO21x1_ASAP7_75t_L g1293 ( 
.A1(n_1148),
.A2(n_838),
.B(n_892),
.Y(n_1293)
);

AO21x1_ASAP7_75t_L g1294 ( 
.A1(n_1110),
.A2(n_838),
.B(n_866),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1140),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_SL g1296 ( 
.A1(n_1161),
.A2(n_857),
.B1(n_898),
.B2(n_894),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1069),
.A2(n_866),
.B(n_1007),
.Y(n_1297)
);

AO21x1_ASAP7_75t_L g1298 ( 
.A1(n_1110),
.A2(n_67),
.B(n_71),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1086),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1168),
.B(n_857),
.Y(n_1300)
);

NAND2x1p5_ASAP7_75t_L g1301 ( 
.A(n_1122),
.B(n_955),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1040),
.B(n_955),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1043),
.B(n_1007),
.Y(n_1303)
);

OA21x2_ASAP7_75t_L g1304 ( 
.A1(n_1027),
.A2(n_67),
.B(n_72),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1102),
.A2(n_986),
.B1(n_875),
.B2(n_73),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1088),
.Y(n_1306)
);

INVxp67_ASAP7_75t_SL g1307 ( 
.A(n_1094),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1062),
.A2(n_986),
.B(n_1054),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1075),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1146),
.A2(n_1078),
.B(n_1144),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1051),
.B(n_1052),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_1082),
.Y(n_1312)
);

AO21x2_ASAP7_75t_L g1313 ( 
.A1(n_1130),
.A2(n_1085),
.B(n_1024),
.Y(n_1313)
);

INVx4_ASAP7_75t_L g1314 ( 
.A(n_1043),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1146),
.A2(n_1078),
.B(n_1144),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1102),
.A2(n_1147),
.B1(n_1150),
.B2(n_1117),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1145),
.A2(n_1047),
.B(n_1088),
.Y(n_1317)
);

OA21x2_ASAP7_75t_L g1318 ( 
.A1(n_1171),
.A2(n_1184),
.B(n_1183),
.Y(n_1318)
);

OAI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1053),
.A2(n_1123),
.B1(n_1128),
.B2(n_1108),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1117),
.A2(n_1043),
.B1(n_1042),
.B2(n_1171),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1065),
.B(n_1156),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1145),
.A2(n_1047),
.B(n_1055),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1049),
.A2(n_1055),
.B(n_1093),
.Y(n_1323)
);

NAND3xp33_ASAP7_75t_L g1324 ( 
.A(n_1180),
.B(n_1065),
.C(n_1163),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1132),
.B(n_1129),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1049),
.A2(n_1093),
.B(n_1089),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1136),
.B(n_1098),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1090),
.A2(n_1160),
.B(n_1037),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1114),
.B(n_1116),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1077),
.B(n_1079),
.Y(n_1330)
);

AOI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1125),
.A2(n_1030),
.B(n_1067),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1112),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1136),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1076),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1136),
.B(n_1173),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1172),
.A2(n_1184),
.B(n_1183),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1172),
.A2(n_1177),
.B(n_1139),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1100),
.A2(n_1101),
.B1(n_1135),
.B2(n_1103),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1112),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1116),
.B(n_1056),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_SL g1341 ( 
.A1(n_1165),
.A2(n_1153),
.B(n_1151),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1160),
.A2(n_1158),
.B(n_1152),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1136),
.B(n_1177),
.Y(n_1343)
);

AO21x2_ASAP7_75t_L g1344 ( 
.A1(n_1106),
.A2(n_1038),
.B(n_1036),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1056),
.A2(n_1158),
.B(n_1152),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1106),
.A2(n_1103),
.B1(n_1116),
.B2(n_1039),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1116),
.B(n_1076),
.Y(n_1347)
);

INVxp67_ASAP7_75t_L g1348 ( 
.A(n_1112),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1057),
.A2(n_1039),
.B(n_1076),
.Y(n_1349)
);

INVxp67_ASAP7_75t_L g1350 ( 
.A(n_1112),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1039),
.B(n_1057),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1287),
.A2(n_1039),
.B1(n_1057),
.B2(n_1076),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1225),
.A2(n_1057),
.B1(n_1324),
.B2(n_1203),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1311),
.B(n_1193),
.Y(n_1354)
);

INVx4_ASAP7_75t_L g1355 ( 
.A(n_1271),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1235),
.B(n_1311),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1249),
.A2(n_1305),
.B1(n_1287),
.B2(n_1308),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1283),
.B(n_1281),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1186),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1246),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1241),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1316),
.A2(n_1249),
.B1(n_1282),
.B2(n_1305),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1283),
.B(n_1279),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1277),
.B(n_1231),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1232),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1312),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1189),
.B(n_1314),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1198),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1349),
.A2(n_1341),
.B(n_1328),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1316),
.A2(n_1206),
.B(n_1221),
.Y(n_1370)
);

OAI221xp5_ASAP7_75t_L g1371 ( 
.A1(n_1206),
.A2(n_1278),
.B1(n_1221),
.B2(n_1274),
.C(n_1285),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1189),
.B(n_1314),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1216),
.B(n_1300),
.Y(n_1373)
);

CKINVDCx6p67_ASAP7_75t_R g1374 ( 
.A(n_1187),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1236),
.Y(n_1375)
);

OAI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1277),
.A2(n_1227),
.B1(n_1202),
.B2(n_1194),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_SL g1377 ( 
.A(n_1319),
.B(n_1239),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1205),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1208),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1283),
.B(n_1189),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1213),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1283),
.B(n_1327),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1280),
.B(n_1240),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1197),
.B(n_1259),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1247),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1248),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1239),
.A2(n_1190),
.B1(n_1274),
.B2(n_1264),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1192),
.A2(n_1196),
.B(n_1264),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1302),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1254),
.A2(n_1286),
.B1(n_1222),
.B2(n_1197),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1197),
.A2(n_1312),
.B1(n_1269),
.B2(n_1321),
.Y(n_1391)
);

INVxp33_ASAP7_75t_L g1392 ( 
.A(n_1255),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1251),
.A2(n_1330),
.B1(n_1210),
.B2(n_1272),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1251),
.A2(n_1330),
.B1(n_1298),
.B2(n_1270),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1215),
.Y(n_1395)
);

CKINVDCx20_ASAP7_75t_R g1396 ( 
.A(n_1200),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1260),
.B(n_1262),
.Y(n_1397)
);

INVx4_ASAP7_75t_SL g1398 ( 
.A(n_1218),
.Y(n_1398)
);

INVx3_ASAP7_75t_L g1399 ( 
.A(n_1302),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1190),
.B(n_1302),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1288),
.B(n_1325),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1213),
.Y(n_1402)
);

AOI221xp5_ASAP7_75t_L g1403 ( 
.A1(n_1268),
.A2(n_1228),
.B1(n_1319),
.B2(n_1207),
.C(n_1185),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1330),
.A2(n_1270),
.B1(n_1263),
.B2(n_1220),
.Y(n_1404)
);

INVx4_ASAP7_75t_L g1405 ( 
.A(n_1271),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1200),
.Y(n_1406)
);

AOI21xp33_ASAP7_75t_L g1407 ( 
.A1(n_1268),
.A2(n_1201),
.B(n_1220),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1266),
.B(n_1215),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1190),
.A2(n_1296),
.B1(n_1320),
.B2(n_1288),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1220),
.A2(n_1200),
.B1(n_1201),
.B2(n_1261),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1288),
.B(n_1261),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1303),
.Y(n_1412)
);

AND2x6_ASAP7_75t_L g1413 ( 
.A(n_1309),
.B(n_1334),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1201),
.A2(n_1261),
.B1(n_1294),
.B2(n_1223),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_SL g1415 ( 
.A(n_1293),
.B(n_1320),
.Y(n_1415)
);

BUFx10_ASAP7_75t_L g1416 ( 
.A(n_1303),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1265),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1223),
.A2(n_1187),
.B1(n_1195),
.B2(n_1303),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1295),
.A2(n_1234),
.B1(n_1219),
.B2(n_1338),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1265),
.Y(n_1420)
);

AOI221xp5_ASAP7_75t_L g1421 ( 
.A1(n_1228),
.A2(n_1335),
.B1(n_1351),
.B2(n_1333),
.C(n_1343),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1223),
.A2(n_1195),
.B1(n_1304),
.B2(n_1214),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1217),
.B(n_1284),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1284),
.B(n_1290),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1252),
.A2(n_1191),
.B(n_1224),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1219),
.B(n_1234),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1290),
.B(n_1291),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1291),
.B(n_1214),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1258),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1276),
.Y(n_1430)
);

INVx4_ASAP7_75t_L g1431 ( 
.A(n_1271),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1214),
.B(n_1307),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_1276),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1219),
.B(n_1234),
.Y(n_1434)
);

INVx4_ASAP7_75t_L g1435 ( 
.A(n_1209),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1334),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1329),
.B(n_1188),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1332),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1243),
.B(n_1304),
.Y(n_1439)
);

BUFx4f_ASAP7_75t_L g1440 ( 
.A(n_1209),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1304),
.A2(n_1267),
.B1(n_1309),
.B2(n_1199),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1346),
.A2(n_1243),
.B1(n_1188),
.B2(n_1257),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1257),
.B(n_1233),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1218),
.B(n_1209),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1276),
.B(n_1218),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1209),
.B(n_1212),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1243),
.B(n_1218),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1212),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1212),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1351),
.A2(n_1348),
.B1(n_1350),
.B2(n_1340),
.C(n_1339),
.Y(n_1450)
);

OR2x6_ASAP7_75t_L g1451 ( 
.A(n_1252),
.B(n_1230),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1243),
.B(n_1347),
.Y(n_1452)
);

INVx3_ASAP7_75t_SL g1453 ( 
.A(n_1212),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1301),
.A2(n_1204),
.B1(n_1229),
.B2(n_1233),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1267),
.B(n_1230),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1199),
.A2(n_1313),
.B1(n_1226),
.B2(n_1191),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1253),
.A2(n_1256),
.B1(n_1250),
.B2(n_1337),
.Y(n_1457)
);

OAI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1233),
.A2(n_1301),
.B1(n_1331),
.B2(n_1273),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1245),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1318),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1233),
.B(n_1318),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1318),
.Y(n_1462)
);

OAI21xp33_ASAP7_75t_SL g1463 ( 
.A1(n_1226),
.A2(n_1256),
.B(n_1253),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1336),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1336),
.B(n_1289),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1289),
.B(n_1297),
.Y(n_1466)
);

AO21x2_ASAP7_75t_L g1467 ( 
.A1(n_1328),
.A2(n_1275),
.B(n_1326),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1323),
.A2(n_1322),
.B(n_1211),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1313),
.B(n_1250),
.Y(n_1469)
);

OAI22x1_ASAP7_75t_L g1470 ( 
.A1(n_1337),
.A2(n_1336),
.B1(n_1345),
.B2(n_1237),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1237),
.B(n_1297),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1245),
.B(n_1238),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1337),
.B(n_1237),
.Y(n_1473)
);

OR2x6_ASAP7_75t_L g1474 ( 
.A(n_1238),
.B(n_1323),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1345),
.B(n_1306),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1292),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1345),
.B(n_1299),
.Y(n_1477)
);

NAND2xp33_ASAP7_75t_SL g1478 ( 
.A(n_1344),
.B(n_1342),
.Y(n_1478)
);

CKINVDCx20_ASAP7_75t_R g1479 ( 
.A(n_1344),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1244),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1244),
.Y(n_1481)
);

AO32x2_ASAP7_75t_L g1482 ( 
.A1(n_1322),
.A2(n_1342),
.A3(n_1211),
.B1(n_1326),
.B2(n_1317),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1317),
.Y(n_1483)
);

NOR3xp33_ASAP7_75t_SL g1484 ( 
.A(n_1310),
.B(n_713),
.C(n_1203),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1310),
.Y(n_1485)
);

INVx6_ASAP7_75t_L g1486 ( 
.A(n_1315),
.Y(n_1486)
);

BUFx4f_ASAP7_75t_SL g1487 ( 
.A(n_1315),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1242),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1225),
.A2(n_946),
.B1(n_711),
.B2(n_514),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1311),
.B(n_713),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1242),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1225),
.A2(n_946),
.B1(n_711),
.B2(n_514),
.Y(n_1492)
);

AOI221xp5_ASAP7_75t_L g1493 ( 
.A1(n_1305),
.A2(n_586),
.B1(n_711),
.B2(n_921),
.C(n_529),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1187),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1186),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1242),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1189),
.B(n_1314),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1242),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1225),
.A2(n_946),
.B1(n_711),
.B2(n_514),
.Y(n_1499)
);

NOR2x1_ASAP7_75t_SL g1500 ( 
.A(n_1263),
.B(n_1193),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1316),
.A2(n_921),
.B(n_529),
.C(n_514),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1242),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1241),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1242),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1189),
.B(n_1314),
.Y(n_1505)
);

OR2x6_ASAP7_75t_L g1506 ( 
.A(n_1272),
.B(n_1252),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_SL g1507 ( 
.A1(n_1362),
.A2(n_1370),
.B1(n_1356),
.B2(n_1371),
.Y(n_1507)
);

OAI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1493),
.A2(n_1492),
.B1(n_1499),
.B2(n_1489),
.C(n_1501),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1440),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1357),
.A2(n_1490),
.B1(n_1501),
.B2(n_1390),
.Y(n_1510)
);

INVxp33_ASAP7_75t_L g1511 ( 
.A(n_1364),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1438),
.Y(n_1512)
);

INVxp67_ASAP7_75t_L g1513 ( 
.A(n_1397),
.Y(n_1513)
);

CKINVDCx14_ASAP7_75t_R g1514 ( 
.A(n_1396),
.Y(n_1514)
);

OR2x6_ASAP7_75t_L g1515 ( 
.A(n_1377),
.B(n_1388),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1402),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1361),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1440),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1356),
.A2(n_1387),
.B1(n_1354),
.B2(n_1500),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1403),
.A2(n_1377),
.B1(n_1353),
.B2(n_1503),
.Y(n_1520)
);

OAI221xp5_ASAP7_75t_L g1521 ( 
.A1(n_1373),
.A2(n_1394),
.B1(n_1484),
.B2(n_1404),
.C(n_1391),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1360),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1376),
.A2(n_1366),
.B1(n_1392),
.B2(n_1409),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1419),
.A2(n_1384),
.B1(n_1396),
.B2(n_1400),
.Y(n_1524)
);

AO31x2_ASAP7_75t_L g1525 ( 
.A1(n_1470),
.A2(n_1475),
.A3(n_1483),
.B(n_1466),
.Y(n_1525)
);

AND2x6_ASAP7_75t_SL g1526 ( 
.A(n_1423),
.B(n_1429),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1381),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1415),
.A2(n_1425),
.B(n_1458),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1392),
.A2(n_1401),
.B1(n_1400),
.B2(n_1399),
.Y(n_1529)
);

AOI222xp33_ASAP7_75t_L g1530 ( 
.A1(n_1415),
.A2(n_1365),
.B1(n_1439),
.B2(n_1406),
.C1(n_1358),
.C2(n_1488),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1389),
.A2(n_1412),
.B1(n_1399),
.B2(n_1434),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1439),
.A2(n_1382),
.B1(n_1479),
.B2(n_1433),
.Y(n_1532)
);

AOI222xp33_ASAP7_75t_L g1533 ( 
.A1(n_1358),
.A2(n_1502),
.B1(n_1491),
.B2(n_1504),
.C1(n_1496),
.C2(n_1498),
.Y(n_1533)
);

OR2x6_ASAP7_75t_L g1534 ( 
.A(n_1506),
.B(n_1434),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1478),
.A2(n_1441),
.B(n_1454),
.Y(n_1535)
);

CKINVDCx6p67_ASAP7_75t_R g1536 ( 
.A(n_1433),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1446),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1478),
.A2(n_1469),
.B(n_1369),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1410),
.A2(n_1418),
.B1(n_1494),
.B2(n_1393),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1411),
.Y(n_1540)
);

AOI21xp33_ASAP7_75t_L g1541 ( 
.A1(n_1352),
.A2(n_1422),
.B(n_1428),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_SL g1542 ( 
.A1(n_1382),
.A2(n_1479),
.B1(n_1447),
.B2(n_1380),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1447),
.A2(n_1380),
.B1(n_1452),
.B2(n_1363),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1383),
.Y(n_1544)
);

NAND3xp33_ASAP7_75t_L g1545 ( 
.A(n_1421),
.B(n_1407),
.C(n_1414),
.Y(n_1545)
);

AOI221xp5_ASAP7_75t_L g1546 ( 
.A1(n_1442),
.A2(n_1450),
.B1(n_1386),
.B2(n_1385),
.C(n_1375),
.Y(n_1546)
);

INVxp33_ASAP7_75t_L g1547 ( 
.A(n_1367),
.Y(n_1547)
);

AOI221x1_ASAP7_75t_SL g1548 ( 
.A1(n_1445),
.A2(n_1437),
.B1(n_1476),
.B2(n_1495),
.C(n_1368),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1412),
.A2(n_1372),
.B1(n_1497),
.B2(n_1367),
.Y(n_1549)
);

OAI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1494),
.A2(n_1374),
.B1(n_1426),
.B2(n_1430),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1359),
.Y(n_1551)
);

A2O1A1Ixp33_ASAP7_75t_SL g1552 ( 
.A1(n_1456),
.A2(n_1459),
.B(n_1379),
.C(n_1495),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1436),
.Y(n_1553)
);

OAI211xp5_ASAP7_75t_L g1554 ( 
.A1(n_1383),
.A2(n_1432),
.B(n_1368),
.C(n_1379),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1367),
.B(n_1497),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1372),
.A2(n_1497),
.B1(n_1505),
.B2(n_1363),
.Y(n_1556)
);

OAI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1374),
.A2(n_1429),
.B1(n_1431),
.B2(n_1355),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1372),
.B(n_1505),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1378),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1369),
.A2(n_1473),
.B(n_1470),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1443),
.B(n_1446),
.Y(n_1561)
);

OAI211xp5_ASAP7_75t_SL g1562 ( 
.A1(n_1444),
.A2(n_1463),
.B(n_1457),
.C(n_1471),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1408),
.B(n_1395),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1424),
.A2(n_1427),
.B1(n_1395),
.B2(n_1420),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1424),
.B(n_1427),
.Y(n_1565)
);

INVx3_ASAP7_75t_L g1566 ( 
.A(n_1355),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1355),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1413),
.A2(n_1405),
.B1(n_1431),
.B2(n_1416),
.Y(n_1568)
);

BUFx12f_ASAP7_75t_L g1569 ( 
.A(n_1448),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1468),
.A2(n_1480),
.B(n_1485),
.Y(n_1570)
);

AOI21xp33_ASAP7_75t_L g1571 ( 
.A1(n_1506),
.A2(n_1455),
.B(n_1481),
.Y(n_1571)
);

OAI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1405),
.A2(n_1431),
.B1(n_1440),
.B2(n_1453),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1413),
.A2(n_1416),
.B1(n_1455),
.B2(n_1506),
.Y(n_1573)
);

OAI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1506),
.A2(n_1405),
.B1(n_1449),
.B2(n_1453),
.C(n_1451),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1443),
.B(n_1446),
.Y(n_1575)
);

OAI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1417),
.A2(n_1420),
.B1(n_1435),
.B2(n_1448),
.Y(n_1576)
);

OAI222xp33_ASAP7_75t_L g1577 ( 
.A1(n_1435),
.A2(n_1451),
.B1(n_1443),
.B2(n_1461),
.C1(n_1477),
.C2(n_1474),
.Y(n_1577)
);

OAI21xp33_ASAP7_75t_L g1578 ( 
.A1(n_1451),
.A2(n_1465),
.B(n_1461),
.Y(n_1578)
);

AOI221xp5_ASAP7_75t_L g1579 ( 
.A1(n_1462),
.A2(n_1472),
.B1(n_1465),
.B2(n_1460),
.C(n_1464),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1413),
.A2(n_1472),
.B1(n_1398),
.B2(n_1435),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1460),
.A2(n_1464),
.B1(n_1459),
.B2(n_1480),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1459),
.A2(n_1487),
.B1(n_1467),
.B2(n_1451),
.Y(n_1582)
);

OAI221xp5_ASAP7_75t_L g1583 ( 
.A1(n_1474),
.A2(n_1486),
.B1(n_1467),
.B2(n_1482),
.C(n_1468),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1467),
.B(n_1474),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1474),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1482),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1486),
.A2(n_1493),
.B1(n_977),
.B2(n_529),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1482),
.A2(n_1493),
.B1(n_1357),
.B2(n_946),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1482),
.A2(n_1493),
.B1(n_1357),
.B2(n_921),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1493),
.A2(n_1357),
.B1(n_946),
.B2(n_1489),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1402),
.Y(n_1591)
);

INVxp33_ASAP7_75t_L g1592 ( 
.A(n_1364),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1493),
.A2(n_977),
.B1(n_529),
.B2(n_514),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1438),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1384),
.B(n_1249),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_SL g1596 ( 
.A1(n_1501),
.A2(n_611),
.B(n_1264),
.Y(n_1596)
);

OAI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1362),
.A2(n_977),
.B1(n_1059),
.B2(n_1493),
.Y(n_1597)
);

AOI221xp5_ASAP7_75t_L g1598 ( 
.A1(n_1493),
.A2(n_1501),
.B1(n_1489),
.B2(n_1499),
.C(n_1492),
.Y(n_1598)
);

CKINVDCx6p67_ASAP7_75t_R g1599 ( 
.A(n_1396),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1490),
.B(n_833),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1493),
.A2(n_977),
.B1(n_529),
.B2(n_514),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1493),
.A2(n_1501),
.B1(n_1489),
.B2(n_1499),
.C(n_1492),
.Y(n_1602)
);

OAI211xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1493),
.A2(n_746),
.B(n_1357),
.C(n_1305),
.Y(n_1603)
);

OR2x6_ASAP7_75t_L g1604 ( 
.A(n_1370),
.B(n_1377),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1384),
.B(n_1437),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1357),
.A2(n_1493),
.B1(n_1490),
.B2(n_1059),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1493),
.A2(n_1357),
.B1(n_946),
.B2(n_1489),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1402),
.Y(n_1608)
);

OAI221xp5_ASAP7_75t_L g1609 ( 
.A1(n_1493),
.A2(n_1492),
.B1(n_1499),
.B2(n_1489),
.C(n_921),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1493),
.A2(n_1357),
.B1(n_946),
.B2(n_1489),
.Y(n_1610)
);

A2O1A1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1493),
.A2(n_514),
.B(n_529),
.C(n_1501),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1493),
.A2(n_1357),
.B1(n_921),
.B2(n_1362),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_SL g1613 ( 
.A1(n_1357),
.A2(n_1305),
.B1(n_1277),
.B2(n_1287),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_SL g1614 ( 
.A1(n_1362),
.A2(n_1370),
.B1(n_1287),
.B2(n_458),
.Y(n_1614)
);

OAI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1493),
.A2(n_1492),
.B1(n_1499),
.B2(n_1489),
.C(n_921),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1534),
.B(n_1585),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1614),
.A2(n_1612),
.B1(n_1590),
.B2(n_1607),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1512),
.Y(n_1618)
);

INVxp67_ASAP7_75t_SL g1619 ( 
.A(n_1553),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1594),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1525),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1570),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1543),
.B(n_1542),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1525),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1543),
.B(n_1542),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1525),
.B(n_1586),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1603),
.A2(n_1614),
.B1(n_1613),
.B2(n_1606),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1525),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1581),
.B(n_1532),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1581),
.B(n_1532),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1553),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1534),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1578),
.B(n_1584),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1604),
.B(n_1582),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1533),
.B(n_1595),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1610),
.A2(n_1612),
.B1(n_1597),
.B2(n_1508),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1551),
.Y(n_1637)
);

AO22x1_ASAP7_75t_L g1638 ( 
.A1(n_1510),
.A2(n_1539),
.B1(n_1547),
.B2(n_1592),
.Y(n_1638)
);

BUFx6f_ASAP7_75t_L g1639 ( 
.A(n_1515),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1534),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1559),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1514),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1593),
.B(n_1601),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1515),
.B(n_1573),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1544),
.B(n_1513),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1604),
.B(n_1582),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1604),
.B(n_1571),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1560),
.B(n_1583),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1516),
.Y(n_1649)
);

INVx1_ASAP7_75t_SL g1650 ( 
.A(n_1527),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1522),
.Y(n_1651)
);

INVxp67_ASAP7_75t_L g1652 ( 
.A(n_1554),
.Y(n_1652)
);

INVx4_ASAP7_75t_L g1653 ( 
.A(n_1515),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1538),
.B(n_1528),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1579),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1513),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1544),
.B(n_1548),
.Y(n_1657)
);

AND3x1_ASAP7_75t_L g1658 ( 
.A(n_1611),
.B(n_1602),
.C(n_1598),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1591),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1530),
.B(n_1519),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1563),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1605),
.B(n_1507),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1565),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1580),
.B(n_1535),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1574),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1597),
.A2(n_1615),
.B1(n_1609),
.B2(n_1589),
.C(n_1588),
.Y(n_1666)
);

NAND3xp33_ASAP7_75t_L g1667 ( 
.A(n_1587),
.B(n_1520),
.C(n_1507),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1519),
.B(n_1556),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1561),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1562),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1545),
.Y(n_1671)
);

BUFx3_ASAP7_75t_L g1672 ( 
.A(n_1608),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1577),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1537),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1596),
.A2(n_1552),
.B(n_1589),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1618),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1618),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_R g1678 ( 
.A(n_1642),
.B(n_1599),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1667),
.A2(n_1521),
.B1(n_1511),
.B2(n_1523),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1648),
.B(n_1517),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1637),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1648),
.B(n_1540),
.Y(n_1682)
);

AOI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1658),
.A2(n_1520),
.B1(n_1523),
.B2(n_1546),
.C(n_1541),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_1649),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1667),
.A2(n_1524),
.B1(n_1529),
.B2(n_1600),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1658),
.B(n_1550),
.C(n_1557),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_SL g1687 ( 
.A1(n_1617),
.A2(n_1558),
.B1(n_1555),
.B2(n_1509),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1663),
.B(n_1564),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1627),
.A2(n_1568),
.B1(n_1550),
.B2(n_1557),
.Y(n_1689)
);

AOI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1617),
.A2(n_1576),
.B1(n_1564),
.B2(n_1572),
.C(n_1531),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1637),
.Y(n_1691)
);

OAI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1622),
.A2(n_1549),
.B(n_1567),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1652),
.A2(n_1572),
.B(n_1576),
.Y(n_1693)
);

OA21x2_ASAP7_75t_L g1694 ( 
.A1(n_1675),
.A2(n_1575),
.B(n_1568),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1663),
.B(n_1526),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1620),
.Y(n_1696)
);

OA21x2_ASAP7_75t_L g1697 ( 
.A1(n_1675),
.A2(n_1569),
.B(n_1566),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1627),
.A2(n_1509),
.B1(n_1518),
.B2(n_1536),
.C(n_1636),
.Y(n_1698)
);

OAI31xp33_ASAP7_75t_L g1699 ( 
.A1(n_1643),
.A2(n_1509),
.A3(n_1518),
.B(n_1636),
.Y(n_1699)
);

A2O1A1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1643),
.A2(n_1666),
.B(n_1660),
.C(n_1652),
.Y(n_1700)
);

OA21x2_ASAP7_75t_L g1701 ( 
.A1(n_1621),
.A2(n_1509),
.B(n_1518),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1671),
.A2(n_1518),
.B1(n_1660),
.B2(n_1666),
.C(n_1655),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1672),
.Y(n_1703)
);

OAI21xp33_ASAP7_75t_L g1704 ( 
.A1(n_1660),
.A2(n_1671),
.B(n_1670),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1620),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1638),
.A2(n_1654),
.B(n_1671),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1641),
.Y(n_1707)
);

OAI31xp33_ASAP7_75t_L g1708 ( 
.A1(n_1670),
.A2(n_1655),
.A3(n_1668),
.B(n_1623),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1672),
.Y(n_1709)
);

A2O1A1Ixp33_ASAP7_75t_L g1710 ( 
.A1(n_1668),
.A2(n_1655),
.B(n_1664),
.C(n_1654),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1633),
.B(n_1634),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1633),
.B(n_1634),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1616),
.B(n_1632),
.Y(n_1713)
);

OAI33xp33_ASAP7_75t_L g1714 ( 
.A1(n_1657),
.A2(n_1635),
.A3(n_1662),
.B1(n_1654),
.B2(n_1645),
.B3(n_1651),
.Y(n_1714)
);

NAND2xp33_ASAP7_75t_R g1715 ( 
.A(n_1669),
.B(n_1635),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1650),
.B(n_1661),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1648),
.B(n_1633),
.Y(n_1717)
);

NAND4xp25_ASAP7_75t_L g1718 ( 
.A(n_1662),
.B(n_1657),
.C(n_1623),
.D(n_1625),
.Y(n_1718)
);

NOR4xp25_ASAP7_75t_SL g1719 ( 
.A(n_1621),
.B(n_1628),
.C(n_1624),
.D(n_1638),
.Y(n_1719)
);

BUFx3_ASAP7_75t_L g1720 ( 
.A(n_1672),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1717),
.B(n_1626),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1717),
.B(n_1626),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1680),
.B(n_1626),
.Y(n_1723)
);

OAI21xp33_ASAP7_75t_L g1724 ( 
.A1(n_1700),
.A2(n_1623),
.B(n_1625),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1711),
.B(n_1647),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1711),
.B(n_1712),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1680),
.B(n_1656),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1681),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1716),
.B(n_1621),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1691),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1706),
.B(n_1656),
.Y(n_1731)
);

NOR4xp25_ASAP7_75t_SL g1732 ( 
.A(n_1715),
.B(n_1628),
.C(n_1624),
.D(n_1619),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1682),
.B(n_1628),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1707),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1713),
.B(n_1647),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1713),
.B(n_1692),
.Y(n_1736)
);

INVx1_ASAP7_75t_SL g1737 ( 
.A(n_1682),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1676),
.B(n_1631),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1676),
.B(n_1631),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1713),
.B(n_1624),
.Y(n_1740)
);

INVx1_ASAP7_75t_SL g1741 ( 
.A(n_1703),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1695),
.B(n_1659),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1677),
.Y(n_1743)
);

NAND2xp33_ASAP7_75t_L g1744 ( 
.A(n_1686),
.B(n_1665),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1713),
.B(n_1647),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1708),
.B(n_1686),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1684),
.B(n_1674),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1684),
.B(n_1646),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1696),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1696),
.B(n_1674),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1701),
.B(n_1646),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1701),
.B(n_1646),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1701),
.B(n_1634),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1705),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1754),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1741),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1735),
.B(n_1673),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1743),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1754),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_SL g1760 ( 
.A1(n_1746),
.A2(n_1710),
.B(n_1704),
.Y(n_1760)
);

AOI31xp33_ASAP7_75t_SL g1761 ( 
.A1(n_1731),
.A2(n_1683),
.A3(n_1702),
.B(n_1679),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1740),
.B(n_1632),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1754),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1742),
.B(n_1718),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1743),
.Y(n_1765)
);

NOR2x1_ASAP7_75t_L g1766 ( 
.A(n_1741),
.B(n_1709),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1735),
.B(n_1673),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1745),
.B(n_1720),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1749),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1749),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1745),
.B(n_1720),
.Y(n_1771)
);

INVxp67_ASAP7_75t_L g1772 ( 
.A(n_1744),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1750),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1737),
.B(n_1650),
.Y(n_1774)
);

AOI21xp33_ASAP7_75t_L g1775 ( 
.A1(n_1724),
.A2(n_1704),
.B(n_1708),
.Y(n_1775)
);

AOI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1724),
.A2(n_1689),
.B1(n_1714),
.B2(n_1718),
.Y(n_1776)
);

OR2x2_ASAP7_75t_SL g1777 ( 
.A(n_1731),
.B(n_1697),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1730),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1750),
.Y(n_1779)
);

AND2x4_ASAP7_75t_SL g1780 ( 
.A(n_1748),
.B(n_1639),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1730),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1738),
.Y(n_1782)
);

NOR2x1_ASAP7_75t_L g1783 ( 
.A(n_1737),
.B(n_1709),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1738),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1727),
.B(n_1665),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1721),
.B(n_1688),
.Y(n_1786)
);

BUFx3_ASAP7_75t_L g1787 ( 
.A(n_1747),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1739),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1728),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_SL g1790 ( 
.A(n_1727),
.B(n_1699),
.Y(n_1790)
);

NAND2x1p5_ASAP7_75t_L g1791 ( 
.A(n_1733),
.B(n_1697),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1759),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1757),
.B(n_1740),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1757),
.B(n_1767),
.Y(n_1794)
);

AOI31xp33_ASAP7_75t_L g1795 ( 
.A1(n_1775),
.A2(n_1776),
.A3(n_1772),
.B(n_1760),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1765),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1783),
.B(n_1736),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1786),
.B(n_1782),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1786),
.B(n_1722),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1759),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_L g1801 ( 
.A(n_1760),
.B(n_1732),
.C(n_1699),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_R g1802 ( 
.A(n_1756),
.B(n_1659),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_1766),
.Y(n_1803)
);

INVx1_ASAP7_75t_SL g1804 ( 
.A(n_1777),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1767),
.B(n_1736),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1762),
.B(n_1740),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1765),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1769),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1769),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1764),
.A2(n_1698),
.B(n_1685),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1770),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1770),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1782),
.B(n_1722),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1784),
.B(n_1723),
.Y(n_1814)
);

NAND3xp33_ASAP7_75t_L g1815 ( 
.A(n_1790),
.B(n_1732),
.C(n_1719),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1784),
.B(n_1723),
.Y(n_1816)
);

OA21x2_ASAP7_75t_L g1817 ( 
.A1(n_1755),
.A2(n_1692),
.B(n_1736),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1787),
.Y(n_1818)
);

OAI21xp33_ASAP7_75t_SL g1819 ( 
.A1(n_1768),
.A2(n_1625),
.B(n_1726),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1758),
.Y(n_1820)
);

AOI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1761),
.A2(n_1690),
.B1(n_1693),
.B2(n_1668),
.C(n_1629),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1787),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1785),
.A2(n_1664),
.B1(n_1644),
.B2(n_1687),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1791),
.B(n_1736),
.Y(n_1824)
);

AOI21xp33_ASAP7_75t_SL g1825 ( 
.A1(n_1791),
.A2(n_1697),
.B(n_1678),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1778),
.Y(n_1826)
);

INVxp67_ASAP7_75t_SL g1827 ( 
.A(n_1778),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1789),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_L g1829 ( 
.A(n_1774),
.B(n_1726),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1788),
.B(n_1729),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1762),
.B(n_1725),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1762),
.B(n_1725),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1789),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1796),
.Y(n_1834)
);

INVx1_ASAP7_75t_SL g1835 ( 
.A(n_1802),
.Y(n_1835)
);

OAI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1801),
.A2(n_1639),
.B1(n_1791),
.B2(n_1653),
.Y(n_1836)
);

AOI21xp33_ASAP7_75t_L g1837 ( 
.A1(n_1795),
.A2(n_1697),
.B(n_1788),
.Y(n_1837)
);

A2O1A1Ixp33_ASAP7_75t_L g1838 ( 
.A1(n_1795),
.A2(n_1780),
.B(n_1753),
.C(n_1751),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1821),
.B(n_1768),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1818),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1821),
.B(n_1771),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1817),
.Y(n_1842)
);

OA21x2_ASAP7_75t_L g1843 ( 
.A1(n_1815),
.A2(n_1781),
.B(n_1755),
.Y(n_1843)
);

AOI21xp33_ASAP7_75t_SL g1844 ( 
.A1(n_1801),
.A2(n_1777),
.B(n_1694),
.Y(n_1844)
);

OAI21xp5_ASAP7_75t_SL g1845 ( 
.A1(n_1810),
.A2(n_1664),
.B(n_1629),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1796),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1807),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1817),
.Y(n_1848)
);

AOI21xp33_ASAP7_75t_L g1849 ( 
.A1(n_1804),
.A2(n_1694),
.B(n_1729),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1817),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1807),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1810),
.B(n_1771),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1808),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1818),
.B(n_1773),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1829),
.B(n_1780),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1817),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1815),
.A2(n_1719),
.B1(n_1664),
.B2(n_1752),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1831),
.B(n_1773),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1831),
.B(n_1779),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1797),
.Y(n_1860)
);

NOR2xp67_ASAP7_75t_L g1861 ( 
.A(n_1825),
.B(n_1763),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1832),
.B(n_1779),
.Y(n_1862)
);

AOI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1804),
.A2(n_1664),
.B1(n_1694),
.B2(n_1630),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1817),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1803),
.A2(n_1639),
.B1(n_1630),
.B2(n_1629),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1823),
.A2(n_1644),
.B1(n_1630),
.B2(n_1639),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1818),
.B(n_1748),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1808),
.Y(n_1868)
);

OAI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1803),
.A2(n_1751),
.B(n_1752),
.Y(n_1869)
);

OAI22xp33_ASAP7_75t_SL g1870 ( 
.A1(n_1839),
.A2(n_1822),
.B1(n_1797),
.B2(n_1798),
.Y(n_1870)
);

NAND2xp33_ASAP7_75t_SL g1871 ( 
.A(n_1841),
.B(n_1852),
.Y(n_1871)
);

INVx1_ASAP7_75t_SL g1872 ( 
.A(n_1835),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1834),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1845),
.A2(n_1822),
.B1(n_1819),
.B2(n_1797),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1834),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1846),
.Y(n_1876)
);

AOI222xp33_ASAP7_75t_L g1877 ( 
.A1(n_1845),
.A2(n_1819),
.B1(n_1822),
.B2(n_1798),
.C1(n_1797),
.C2(n_1799),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1846),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1860),
.Y(n_1879)
);

OAI322xp33_ASAP7_75t_L g1880 ( 
.A1(n_1844),
.A2(n_1825),
.A3(n_1799),
.B1(n_1830),
.B2(n_1820),
.C1(n_1813),
.C2(n_1814),
.Y(n_1880)
);

AOI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1857),
.A2(n_1832),
.B1(n_1806),
.B2(n_1794),
.Y(n_1881)
);

NAND4xp25_ASAP7_75t_L g1882 ( 
.A(n_1838),
.B(n_1824),
.C(n_1794),
.D(n_1805),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1860),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1835),
.B(n_1793),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1863),
.A2(n_1843),
.B1(n_1865),
.B2(n_1861),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1858),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1840),
.B(n_1793),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1847),
.Y(n_1888)
);

INVxp67_ASAP7_75t_L g1889 ( 
.A(n_1843),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1847),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1851),
.Y(n_1891)
);

HB1xp67_ASAP7_75t_L g1892 ( 
.A(n_1843),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_SL g1893 ( 
.A1(n_1843),
.A2(n_1827),
.B1(n_1709),
.B2(n_1720),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1851),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1844),
.B(n_1806),
.Y(n_1895)
);

INVx1_ASAP7_75t_SL g1896 ( 
.A(n_1872),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1892),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_R g1898 ( 
.A(n_1871),
.B(n_1855),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1879),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1892),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1886),
.B(n_1879),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1889),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1884),
.B(n_1858),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1889),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1883),
.B(n_1859),
.Y(n_1905)
);

NAND2x1_ASAP7_75t_L g1906 ( 
.A(n_1885),
.B(n_1861),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_1883),
.Y(n_1907)
);

NAND3xp33_ASAP7_75t_SL g1908 ( 
.A(n_1871),
.B(n_1863),
.C(n_1865),
.Y(n_1908)
);

INVxp67_ASAP7_75t_L g1909 ( 
.A(n_1895),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1870),
.B(n_1859),
.Y(n_1910)
);

XNOR2xp5_ASAP7_75t_L g1911 ( 
.A(n_1881),
.B(n_1836),
.Y(n_1911)
);

INVxp67_ASAP7_75t_SL g1912 ( 
.A(n_1893),
.Y(n_1912)
);

NOR2x1_ASAP7_75t_L g1913 ( 
.A(n_1880),
.B(n_1853),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1887),
.Y(n_1914)
);

INVxp67_ASAP7_75t_L g1915 ( 
.A(n_1877),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1896),
.B(n_1874),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1907),
.B(n_1873),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1899),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1909),
.B(n_1882),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_L g1920 ( 
.A(n_1915),
.B(n_1914),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1903),
.B(n_1910),
.Y(n_1921)
);

INVxp67_ASAP7_75t_L g1922 ( 
.A(n_1905),
.Y(n_1922)
);

INVx2_ASAP7_75t_SL g1923 ( 
.A(n_1899),
.Y(n_1923)
);

AOI221xp5_ASAP7_75t_L g1924 ( 
.A1(n_1908),
.A2(n_1837),
.B1(n_1849),
.B2(n_1869),
.C(n_1894),
.Y(n_1924)
);

NOR3xp33_ASAP7_75t_L g1925 ( 
.A(n_1912),
.B(n_1878),
.C(n_1890),
.Y(n_1925)
);

OAI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1906),
.A2(n_1866),
.B1(n_1869),
.B2(n_1867),
.Y(n_1926)
);

AOI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1906),
.A2(n_1854),
.B1(n_1862),
.B2(n_1876),
.Y(n_1927)
);

NAND2xp33_ASAP7_75t_R g1928 ( 
.A(n_1920),
.B(n_1898),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1922),
.B(n_1907),
.Y(n_1929)
);

NAND2xp33_ASAP7_75t_L g1930 ( 
.A(n_1925),
.B(n_1913),
.Y(n_1930)
);

OAI211xp5_ASAP7_75t_SL g1931 ( 
.A1(n_1916),
.A2(n_1913),
.B(n_1904),
.C(n_1897),
.Y(n_1931)
);

NAND3xp33_ASAP7_75t_SL g1932 ( 
.A(n_1924),
.B(n_1900),
.C(n_1897),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_R g1933 ( 
.A(n_1917),
.B(n_1899),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1919),
.B(n_1901),
.Y(n_1934)
);

OAI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1927),
.A2(n_1911),
.B(n_1901),
.Y(n_1935)
);

OAI221xp5_ASAP7_75t_L g1936 ( 
.A1(n_1926),
.A2(n_1911),
.B1(n_1904),
.B2(n_1900),
.C(n_1902),
.Y(n_1936)
);

NOR3xp33_ASAP7_75t_SL g1937 ( 
.A(n_1921),
.B(n_1875),
.C(n_1888),
.Y(n_1937)
);

OAI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1918),
.A2(n_1905),
.B(n_1902),
.Y(n_1938)
);

XNOR2xp5_ASAP7_75t_L g1939 ( 
.A(n_1936),
.B(n_1923),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1935),
.A2(n_1934),
.B1(n_1937),
.B2(n_1929),
.Y(n_1940)
);

NAND3xp33_ASAP7_75t_L g1941 ( 
.A(n_1930),
.B(n_1902),
.C(n_1899),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1938),
.Y(n_1942)
);

NAND4xp75_ASAP7_75t_L g1943 ( 
.A(n_1931),
.B(n_1891),
.C(n_1868),
.D(n_1853),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1933),
.Y(n_1944)
);

NAND2xp33_ASAP7_75t_L g1945 ( 
.A(n_1928),
.B(n_1868),
.Y(n_1945)
);

INVx2_ASAP7_75t_SL g1946 ( 
.A(n_1944),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1941),
.B(n_1862),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1945),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1939),
.B(n_1932),
.Y(n_1949)
);

NAND4xp75_ASAP7_75t_L g1950 ( 
.A(n_1942),
.B(n_1824),
.C(n_1856),
.D(n_1850),
.Y(n_1950)
);

NOR3x1_ASAP7_75t_L g1951 ( 
.A(n_1943),
.B(n_1940),
.C(n_1827),
.Y(n_1951)
);

AOI221xp5_ASAP7_75t_SL g1952 ( 
.A1(n_1949),
.A2(n_1864),
.B1(n_1856),
.B2(n_1850),
.C(n_1848),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_SL g1953 ( 
.A1(n_1948),
.A2(n_1864),
.B1(n_1856),
.B2(n_1850),
.Y(n_1953)
);

NOR3xp33_ASAP7_75t_SL g1954 ( 
.A(n_1950),
.B(n_1830),
.C(n_1816),
.Y(n_1954)
);

INVxp67_ASAP7_75t_SL g1955 ( 
.A(n_1951),
.Y(n_1955)
);

AOI221xp5_ASAP7_75t_L g1956 ( 
.A1(n_1947),
.A2(n_1864),
.B1(n_1848),
.B2(n_1842),
.C(n_1824),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_L g1957 ( 
.A(n_1955),
.B(n_1946),
.Y(n_1957)
);

AOI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1956),
.A2(n_1947),
.B1(n_1848),
.B2(n_1842),
.Y(n_1958)
);

NOR2x1_ASAP7_75t_L g1959 ( 
.A(n_1954),
.B(n_1809),
.Y(n_1959)
);

OAI21x1_ASAP7_75t_L g1960 ( 
.A1(n_1959),
.A2(n_1953),
.B(n_1952),
.Y(n_1960)
);

AOI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1960),
.A2(n_1957),
.B1(n_1958),
.B2(n_1826),
.Y(n_1961)
);

AOI221xp5_ASAP7_75t_R g1962 ( 
.A1(n_1961),
.A2(n_1842),
.B1(n_1640),
.B2(n_1734),
.C(n_1805),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1961),
.Y(n_1963)
);

XNOR2xp5_ASAP7_75t_L g1964 ( 
.A(n_1963),
.B(n_1805),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1962),
.Y(n_1965)
);

AOI222xp33_ASAP7_75t_SL g1966 ( 
.A1(n_1965),
.A2(n_1809),
.B1(n_1811),
.B2(n_1812),
.C1(n_1828),
.C2(n_1833),
.Y(n_1966)
);

AOI22xp33_ASAP7_75t_L g1967 ( 
.A1(n_1964),
.A2(n_1826),
.B1(n_1792),
.B2(n_1800),
.Y(n_1967)
);

AOI22xp5_ASAP7_75t_SL g1968 ( 
.A1(n_1966),
.A2(n_1812),
.B1(n_1811),
.B2(n_1833),
.Y(n_1968)
);

AOI221xp5_ASAP7_75t_L g1969 ( 
.A1(n_1968),
.A2(n_1967),
.B1(n_1820),
.B2(n_1828),
.C(n_1826),
.Y(n_1969)
);

AOI211xp5_ASAP7_75t_L g1970 ( 
.A1(n_1969),
.A2(n_1792),
.B(n_1800),
.C(n_1816),
.Y(n_1970)
);


endmodule