module fake_jpeg_871_n_610 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_610);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_610;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_58),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_59),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_60),
.Y(n_170)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_61),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_63),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_30),
.Y(n_64)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_64),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_65),
.Y(n_175)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_31),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_99),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_23),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_68),
.B(n_76),
.Y(n_157)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_70),
.Y(n_184)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_23),
.B(n_0),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_81),
.Y(n_160)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_83),
.Y(n_171)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_85),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_28),
.B(n_33),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_86),
.B(n_89),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_28),
.B(n_1),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_43),
.B(n_1),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_41),
.Y(n_120)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_31),
.B(n_2),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_98),
.B(n_34),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_20),
.B(n_2),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_35),
.Y(n_100)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_29),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_113),
.Y(n_168)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_29),
.Y(n_114)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_120),
.B(n_3),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_121),
.B(n_163),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_64),
.A2(n_30),
.B1(n_41),
.B2(n_48),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_124),
.A2(n_136),
.B1(n_146),
.B2(n_166),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_57),
.A2(n_30),
.B1(n_48),
.B2(n_41),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_125),
.A2(n_127),
.B1(n_162),
.B2(n_56),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_30),
.B1(n_48),
.B2(n_53),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_58),
.A2(n_25),
.B1(n_47),
.B2(n_26),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_59),
.A2(n_25),
.B1(n_26),
.B2(n_47),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_87),
.A2(n_53),
.B1(n_26),
.B2(n_47),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_62),
.B(n_44),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_77),
.B(n_39),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_164),
.B(n_36),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_70),
.A2(n_56),
.B1(n_45),
.B2(n_25),
.Y(n_166)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_87),
.Y(n_167)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_176),
.Y(n_192)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_72),
.A2(n_56),
.B1(n_34),
.B2(n_53),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_173),
.A2(n_181),
.B1(n_37),
.B2(n_42),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_60),
.B(n_51),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_73),
.A2(n_56),
.B1(n_51),
.B2(n_54),
.Y(n_181)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_185),
.Y(n_290)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

INVxp67_ASAP7_75t_SL g273 ( 
.A(n_188),
.Y(n_273)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_189),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_181),
.A2(n_65),
.B1(n_114),
.B2(n_111),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_190),
.A2(n_208),
.B1(n_83),
.B2(n_78),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_50),
.B1(n_54),
.B2(n_52),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_191),
.A2(n_160),
.B1(n_156),
.B2(n_134),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_46),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_193),
.B(n_196),
.Y(n_269)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_194),
.Y(n_266)
);

INVx3_ASAP7_75t_SL g195 ( 
.A(n_129),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_46),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_197),
.Y(n_275)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_198),
.Y(n_284)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_200),
.Y(n_260)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_202),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_152),
.Y(n_203)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_203),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_119),
.B(n_50),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_204),
.B(n_216),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_129),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_205),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_135),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g289 ( 
.A(n_206),
.B(n_217),
.C(n_219),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_120),
.A2(n_91),
.B1(n_158),
.B2(n_122),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_SL g272 ( 
.A1(n_207),
.A2(n_213),
.B(n_223),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_166),
.A2(n_92),
.B1(n_107),
.B2(n_100),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_117),
.Y(n_209)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_209),
.Y(n_281)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_142),
.Y(n_210)
);

BUFx8_ASAP7_75t_L g297 ( 
.A(n_210),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_140),
.Y(n_211)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_211),
.Y(n_287)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_137),
.Y(n_212)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_212),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_122),
.A2(n_91),
.B1(n_110),
.B2(n_108),
.Y(n_213)
);

INVx11_ASAP7_75t_L g214 ( 
.A(n_142),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_214),
.Y(n_305)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_131),
.Y(n_215)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_215),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_128),
.A2(n_36),
.B(n_52),
.C(n_44),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_135),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_145),
.Y(n_218)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_218),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_142),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_152),
.Y(n_220)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_220),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_130),
.B(n_113),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_221),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_147),
.B(n_141),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_226),
.Y(n_254)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_118),
.Y(n_224)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_224),
.Y(n_310)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_150),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_225),
.B(n_229),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_123),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_230),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_228),
.B(n_233),
.Y(n_296)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_180),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_132),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_182),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_235),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_140),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_232),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_155),
.B(n_42),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_144),
.B(n_37),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_234),
.B(n_247),
.Y(n_301)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_115),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_236),
.A2(n_175),
.B1(n_170),
.B2(n_184),
.Y(n_259)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_115),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_239),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_153),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_238),
.Y(n_256)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_124),
.B(n_97),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_244),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_125),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_242),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_153),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_243),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_154),
.B(n_96),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_116),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_245),
.B(n_248),
.Y(n_292)
);

AND2x2_ASAP7_75t_SL g252 ( 
.A(n_246),
.B(n_148),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_168),
.B(n_3),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_116),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_154),
.B(n_85),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_250),
.Y(n_298)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_134),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_139),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_251),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_252),
.B(n_8),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_216),
.A2(n_127),
.B(n_162),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_253),
.A2(n_300),
.B(n_195),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_259),
.A2(n_264),
.B1(n_268),
.B2(n_283),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_192),
.B(n_139),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_263),
.B(n_270),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_184),
.B1(n_175),
.B2(n_170),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_160),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_186),
.B(n_75),
.C(n_81),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_274),
.B(n_282),
.C(n_302),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_187),
.B(n_71),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_236),
.A2(n_242),
.B1(n_221),
.B2(n_223),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_285),
.A2(n_303),
.B1(n_306),
.B2(n_194),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_229),
.B(n_156),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_295),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_231),
.B(n_3),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_207),
.A2(n_165),
.B(n_55),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_225),
.B(n_174),
.C(n_171),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_223),
.A2(n_171),
.B1(n_174),
.B2(n_55),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_221),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_304),
.A2(n_232),
.B1(n_211),
.B2(n_243),
.Y(n_322)
);

OAI22xp33_ASAP7_75t_L g306 ( 
.A1(n_223),
.A2(n_213),
.B1(n_248),
.B2(n_245),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_290),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_311),
.B(n_323),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_312),
.A2(n_316),
.B1(n_329),
.B2(n_335),
.Y(n_405)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_313),
.Y(n_367)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_292),
.Y(n_314)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_314),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_283),
.A2(n_237),
.B1(n_235),
.B2(n_250),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_317),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_269),
.B(n_215),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_318),
.B(n_336),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_269),
.B(n_296),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_319),
.B(n_340),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_320),
.Y(n_384)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_287),
.Y(n_321)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_321),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_322),
.A2(n_267),
.B1(n_271),
.B2(n_309),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_290),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_261),
.Y(n_324)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_324),
.Y(n_377)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_281),
.Y(n_325)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_325),
.Y(n_381)
);

INVx5_ASAP7_75t_L g328 ( 
.A(n_278),
.Y(n_328)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_328),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_276),
.A2(n_239),
.B1(n_185),
.B2(n_197),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_263),
.B(n_198),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_330),
.B(n_358),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_282),
.B(n_205),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_331),
.B(n_337),
.C(n_345),
.Y(n_379)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_281),
.Y(n_332)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_332),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_303),
.A2(n_272),
.B1(n_256),
.B2(n_294),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_333),
.A2(n_361),
.B1(n_305),
.B2(n_308),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_286),
.A2(n_188),
.B(n_226),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_334),
.A2(n_338),
.B(n_300),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_253),
.A2(n_238),
.B1(n_220),
.B2(n_203),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_301),
.B(n_212),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_252),
.B(n_218),
.Y(n_337)
);

O2A1O1Ixp33_ASAP7_75t_SL g338 ( 
.A1(n_306),
.A2(n_214),
.B(n_199),
.C(n_210),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_280),
.B(n_199),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_339),
.B(n_352),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_289),
.B(n_4),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_290),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_341),
.B(n_348),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_259),
.A2(n_285),
.B1(n_265),
.B2(n_298),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_342),
.A2(n_349),
.B1(n_360),
.B2(n_362),
.Y(n_363)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_344),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_252),
.B(n_5),
.Y(n_345)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_266),
.Y(n_347)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_299),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_265),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_299),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_350),
.B(n_353),
.Y(n_404)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_310),
.Y(n_351)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_258),
.B(n_6),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_258),
.B(n_8),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_297),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_354),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_359),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_299),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_356),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_297),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_357),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_257),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_260),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_270),
.A2(n_17),
.B1(n_10),
.B2(n_11),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_260),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_268),
.A2(n_17),
.B1(n_10),
.B2(n_11),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_346),
.A2(n_254),
.B1(n_256),
.B2(n_294),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_364),
.A2(n_389),
.B(n_397),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_312),
.A2(n_274),
.B1(n_302),
.B2(n_295),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_369),
.A2(n_382),
.B1(n_255),
.B2(n_291),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_313),
.A2(n_304),
.B1(n_262),
.B2(n_279),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_375),
.A2(n_406),
.B1(n_322),
.B2(n_359),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_380),
.A2(n_391),
.B(n_401),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_331),
.B(n_279),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_383),
.B(n_399),
.Y(n_422)
);

OAI32xp33_ASAP7_75t_L g386 ( 
.A1(n_315),
.A2(n_262),
.A3(n_293),
.B1(n_273),
.B2(n_284),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_386),
.B(n_393),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_320),
.A2(n_348),
.B(n_350),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_326),
.B(n_337),
.C(n_315),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_390),
.B(n_392),
.C(n_395),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_334),
.A2(n_297),
.B(n_305),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_326),
.B(n_266),
.C(n_277),
.Y(n_392)
);

OAI32xp33_ASAP7_75t_L g393 ( 
.A1(n_330),
.A2(n_293),
.A3(n_275),
.B1(n_284),
.B2(n_308),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_314),
.B(n_277),
.C(n_309),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_327),
.B(n_307),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_338),
.A2(n_307),
.B(n_255),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_328),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_403),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_342),
.A2(n_278),
.B1(n_267),
.B2(n_275),
.Y(n_406)
);

A2O1A1O1Ixp25_ASAP7_75t_L g409 ( 
.A1(n_390),
.A2(n_327),
.B(n_355),
.C(n_324),
.D(n_358),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_409),
.B(n_423),
.Y(n_467)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_371),
.Y(n_410)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_410),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_384),
.A2(n_335),
.B1(n_316),
.B2(n_362),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_411),
.A2(n_425),
.B1(n_434),
.B2(n_442),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_395),
.Y(n_412)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_412),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_373),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_413),
.B(n_416),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_379),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_414),
.B(n_421),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_415),
.A2(n_420),
.B1(n_426),
.B2(n_428),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_388),
.B(n_361),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_371),
.Y(n_417)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_417),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_376),
.Y(n_418)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_418),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_369),
.A2(n_338),
.B1(n_355),
.B2(n_317),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_379),
.B(n_345),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_394),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_394),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_424),
.B(n_429),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_384),
.A2(n_321),
.B1(n_360),
.B2(n_332),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_363),
.A2(n_351),
.B1(n_343),
.B2(n_325),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_363),
.A2(n_311),
.B1(n_323),
.B2(n_341),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_404),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_430),
.Y(n_471)
);

XNOR2x2_ASAP7_75t_SL g431 ( 
.A(n_389),
.B(n_349),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_380),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_388),
.B(n_347),
.Y(n_432)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_432),
.Y(n_472)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_433),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_364),
.A2(n_357),
.B1(n_354),
.B2(n_344),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_435),
.A2(n_439),
.B1(n_441),
.B2(n_443),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_402),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_436),
.Y(n_470)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_381),
.Y(n_437)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_437),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_367),
.B(n_291),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_438),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_400),
.B(n_9),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_381),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_440),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_402),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_385),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_402),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_392),
.B(n_399),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_365),
.Y(n_462)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_385),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_446),
.A2(n_387),
.B1(n_398),
.B2(n_375),
.Y(n_452)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_452),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_422),
.B(n_377),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_454),
.B(n_465),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_447),
.B(n_367),
.C(n_377),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_455),
.B(n_458),
.C(n_460),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_456),
.A2(n_478),
.B1(n_482),
.B2(n_444),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_370),
.C(n_378),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_445),
.B(n_370),
.C(n_396),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_462),
.B(n_464),
.C(n_480),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_414),
.B(n_396),
.C(n_366),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_422),
.B(n_365),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_421),
.B(n_365),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_466),
.B(n_469),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_434),
.A2(n_374),
.B1(n_406),
.B2(n_405),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_468),
.A2(n_426),
.B(n_415),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_374),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_408),
.B(n_386),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_476),
.B(n_479),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_420),
.A2(n_401),
.B1(n_382),
.B2(n_403),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_409),
.B(n_398),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_423),
.B(n_366),
.C(n_387),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_408),
.A2(n_391),
.B1(n_368),
.B2(n_393),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_448),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_484),
.B(n_498),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_457),
.B(n_427),
.C(n_444),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_486),
.B(n_510),
.C(n_466),
.Y(n_518)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_481),
.Y(n_488)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_488),
.Y(n_514)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_475),
.Y(n_489)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_489),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_461),
.B(n_429),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_490),
.B(n_506),
.Y(n_525)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_475),
.Y(n_491)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_491),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_492),
.A2(n_509),
.B1(n_493),
.B2(n_487),
.Y(n_527)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_480),
.Y(n_493)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_493),
.Y(n_520)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_450),
.Y(n_496)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_496),
.Y(n_521)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_472),
.Y(n_497)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_497),
.Y(n_513)
);

A2O1A1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_467),
.A2(n_427),
.B(n_425),
.C(n_411),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_499),
.A2(n_482),
.B(n_470),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_463),
.A2(n_428),
.B1(n_419),
.B2(n_433),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_500),
.A2(n_508),
.B1(n_478),
.B2(n_512),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_453),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_501),
.B(n_507),
.Y(n_530)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_471),
.Y(n_502)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_502),
.Y(n_529)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_473),
.Y(n_503)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_503),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_468),
.A2(n_446),
.B1(n_417),
.B2(n_440),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_504),
.B(n_512),
.Y(n_532)
);

NAND3xp33_ASAP7_75t_L g506 ( 
.A(n_467),
.B(n_437),
.C(n_430),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_474),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_451),
.A2(n_438),
.B1(n_442),
.B2(n_410),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_477),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_509),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_457),
.B(n_368),
.C(n_407),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_464),
.B(n_407),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_511),
.B(n_462),
.Y(n_528)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_459),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_515),
.A2(n_505),
.B1(n_508),
.B2(n_469),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_518),
.B(n_528),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_500),
.B(n_459),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_522),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_485),
.B(n_460),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_524),
.B(n_526),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_485),
.B(n_455),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_527),
.A2(n_496),
.B1(n_10),
.B2(n_11),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_511),
.B(n_479),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_531),
.B(n_536),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_483),
.B(n_449),
.C(n_458),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_534),
.B(n_483),
.C(n_510),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_535),
.A2(n_498),
.B(n_499),
.Y(n_538)
);

XNOR2x1_ASAP7_75t_L g536 ( 
.A(n_486),
.B(n_456),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_489),
.B(n_476),
.Y(n_537)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_537),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_SL g561 ( 
.A(n_538),
.B(n_552),
.Y(n_561)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_540),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_544),
.B(n_545),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_526),
.B(n_524),
.C(n_534),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_528),
.B(n_505),
.C(n_495),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_546),
.B(n_550),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_515),
.A2(n_491),
.B1(n_497),
.B2(n_495),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_547),
.B(n_554),
.Y(n_560)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_525),
.Y(n_548)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_548),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_520),
.B(n_494),
.C(n_454),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_530),
.Y(n_551)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_551),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_516),
.B(n_484),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_518),
.B(n_494),
.C(n_465),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_553),
.B(n_556),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_535),
.A2(n_9),
.B(n_10),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_555),
.B(n_521),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_531),
.B(n_12),
.C(n_13),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_513),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_557),
.B(n_513),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_545),
.B(n_527),
.C(n_536),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_558),
.B(n_559),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_544),
.B(n_542),
.C(n_541),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_541),
.B(n_522),
.C(n_537),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_562),
.B(n_563),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_549),
.B(n_522),
.C(n_532),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_SL g564 ( 
.A(n_539),
.B(n_514),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_564),
.B(n_573),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_567),
.B(n_555),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_549),
.B(n_532),
.C(n_523),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_568),
.B(n_571),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_547),
.B(n_523),
.C(n_517),
.Y(n_571)
);

XOR2x1_ASAP7_75t_SL g574 ( 
.A(n_538),
.B(n_519),
.Y(n_574)
);

INVxp33_ASAP7_75t_L g583 ( 
.A(n_574),
.Y(n_583)
);

MAJx2_ASAP7_75t_L g577 ( 
.A(n_558),
.B(n_546),
.C(n_540),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_577),
.B(n_581),
.C(n_587),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_562),
.B(n_550),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_578),
.B(n_586),
.Y(n_593)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_580),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_559),
.B(n_553),
.C(n_552),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_568),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_582),
.B(n_569),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_565),
.B(n_519),
.Y(n_585)
);

NAND3xp33_ASAP7_75t_L g594 ( 
.A(n_585),
.B(n_561),
.C(n_572),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_563),
.B(n_556),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_566),
.B(n_554),
.C(n_543),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_589),
.B(n_590),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_582),
.B(n_570),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_594),
.A2(n_595),
.B(n_596),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_588),
.B(n_575),
.C(n_574),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_576),
.B(n_571),
.C(n_560),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_591),
.B(n_584),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_598),
.B(n_599),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_593),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_592),
.A2(n_583),
.B(n_577),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_601),
.Y(n_603)
);

A2O1A1O1Ixp25_ASAP7_75t_L g602 ( 
.A1(n_597),
.A2(n_583),
.B(n_589),
.C(n_579),
.D(n_578),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_602),
.A2(n_600),
.B(n_586),
.Y(n_605)
);

OAI321xp33_ASAP7_75t_L g607 ( 
.A1(n_605),
.A2(n_606),
.A3(n_603),
.B1(n_543),
.B2(n_529),
.C(n_533),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_604),
.B(n_560),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_607),
.A2(n_14),
.B(n_15),
.Y(n_608)
);

OAI211xp5_ASAP7_75t_L g609 ( 
.A1(n_608),
.A2(n_14),
.B(n_16),
.C(n_17),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_SL g610 ( 
.A1(n_609),
.A2(n_16),
.B(n_340),
.Y(n_610)
);


endmodule