module fake_jpeg_20962_n_141 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_19),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_14),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_0),
.B(n_1),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_73),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_1),
.B(n_2),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_2),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_55),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_79),
.Y(n_83)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_51),
.B1(n_57),
.B2(n_67),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_88),
.B1(n_48),
.B2(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_87),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_70),
.B1(n_59),
.B2(n_68),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_64),
.B1(n_54),
.B2(n_52),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_71),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_71),
.B1(n_67),
.B2(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_60),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_102),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_49),
.B1(n_50),
.B2(n_69),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_103),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_3),
.B(n_4),
.Y(n_98)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_98),
.B(n_9),
.CI(n_10),
.CON(n_106),
.SN(n_106)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_31),
.Y(n_115)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_62),
.B1(n_61),
.B2(n_5),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_7),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_25),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_100),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_109),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

OAI32xp33_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_13),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_22),
.Y(n_110)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_28),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_114),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_125)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_125),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_117),
.A2(n_37),
.B1(n_39),
.B2(n_43),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_126),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_108),
.B(n_113),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_129),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_120),
.B1(n_111),
.B2(n_127),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

NAND4xp25_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_130),
.C(n_106),
.D(n_123),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_121),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_121),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_136),
.A2(n_122),
.B(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_118),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_140),
.Y(n_141)
);


endmodule