module fake_jpeg_22777_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx4_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_3),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g17 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_20),
.B(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_15),
.B(n_11),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_29),
.C(n_34),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_15),
.C(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_30),
.B(n_5),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_10),
.B1(n_21),
.B2(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_11),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_6),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_25),
.A2(n_12),
.B(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVxp33_ASAP7_75t_SL g43 ( 
.A(n_36),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_12),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_24),
.C(n_29),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_24),
.C(n_37),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_38),
.B(n_44),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_46),
.C(n_12),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_27),
.Y(n_52)
);

OAI21x1_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_50),
.B(n_10),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_10),
.B1(n_26),
.B2(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_27),
.Y(n_55)
);


endmodule