module real_aes_16083_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_0), .Y(n_557) );
AND2x4_ASAP7_75t_L g116 ( .A(n_1), .B(n_117), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_2), .A2(n_4), .B1(n_273), .B2(n_274), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_3), .A2(n_23), .B1(n_222), .B2(n_256), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g158 ( .A1(n_5), .A2(n_53), .B1(n_159), .B2(n_160), .Y(n_158) );
BUFx3_ASAP7_75t_L g610 ( .A(n_6), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_7), .A2(n_14), .B1(n_174), .B2(n_175), .Y(n_173) );
INVx1_ASAP7_75t_L g117 ( .A(n_8), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_9), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g847 ( .A(n_10), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_11), .B(n_199), .Y(n_588) );
BUFx2_ASAP7_75t_L g108 ( .A(n_12), .Y(n_108) );
OR2x2_ASAP7_75t_L g131 ( .A(n_12), .B(n_32), .Y(n_131) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_13), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_15), .B(n_150), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_16), .B(n_190), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_17), .A2(n_86), .B1(n_150), .B2(n_256), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_18), .A2(n_19), .B1(n_842), .B2(n_843), .Y(n_841) );
INVx1_ASAP7_75t_L g843 ( .A(n_18), .Y(n_843) );
INVx1_ASAP7_75t_L g842 ( .A(n_19), .Y(n_842) );
OAI21x1_ASAP7_75t_L g164 ( .A1(n_20), .A2(n_49), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_21), .B(n_501), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_22), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_24), .B(n_222), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_25), .B(n_147), .Y(n_214) );
INVx4_ASAP7_75t_R g198 ( .A(n_26), .Y(n_198) );
AO32x1_ASAP7_75t_L g526 ( .A1(n_27), .A2(n_210), .A3(n_211), .B1(n_527), .B2(n_530), .Y(n_526) );
AO32x2_ASAP7_75t_L g618 ( .A1(n_27), .A2(n_210), .A3(n_211), .B1(n_527), .B2(n_530), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_28), .B(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g278 ( .A(n_29), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_SL g253 ( .A1(n_30), .A2(n_146), .B(n_174), .C(n_254), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_31), .A2(n_46), .B1(n_174), .B2(n_178), .Y(n_262) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_32), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_33), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_34), .A2(n_52), .B1(n_200), .B2(n_222), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_35), .A2(n_91), .B1(n_178), .B2(n_256), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_36), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_37), .B(n_538), .Y(n_542) );
INVx1_ASAP7_75t_L g218 ( .A(n_38), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_39), .B(n_174), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_40), .A2(n_68), .B1(n_178), .B2(n_566), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_41), .Y(n_232) );
INVx2_ASAP7_75t_L g122 ( .A(n_42), .Y(n_122) );
INVx1_ASAP7_75t_L g111 ( .A(n_43), .Y(n_111) );
BUFx3_ASAP7_75t_L g507 ( .A(n_43), .Y(n_507) );
INVx1_ASAP7_75t_L g494 ( .A(n_44), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_45), .B(n_544), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_47), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_48), .A2(n_85), .B1(n_174), .B2(n_178), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_50), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_51), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_54), .A2(n_79), .B1(n_153), .B2(n_538), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_55), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_56), .A2(n_83), .B1(n_150), .B2(n_256), .Y(n_606) );
INVx1_ASAP7_75t_L g165 ( .A(n_57), .Y(n_165) );
AND2x4_ASAP7_75t_L g168 ( .A(n_58), .B(n_169), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g134 ( .A1(n_59), .A2(n_78), .B1(n_135), .B2(n_136), .Y(n_134) );
INVx1_ASAP7_75t_L g136 ( .A(n_59), .Y(n_136) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_60), .A2(n_90), .B1(n_178), .B2(n_271), .Y(n_270) );
AO22x1_ASAP7_75t_L g148 ( .A1(n_61), .A2(n_73), .B1(n_149), .B2(n_152), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_62), .B(n_256), .Y(n_587) );
INVx1_ASAP7_75t_L g169 ( .A(n_63), .Y(n_169) );
AND2x2_ASAP7_75t_L g257 ( .A(n_64), .B(n_210), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_65), .B(n_210), .Y(n_593) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_66), .A2(n_156), .B(n_159), .C(n_556), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_67), .B(n_256), .C(n_591), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_69), .B(n_159), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_70), .Y(n_248) );
AND2x2_ASAP7_75t_L g558 ( .A(n_71), .B(n_204), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_72), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_74), .B(n_222), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_75), .A2(n_96), .B1(n_150), .B2(n_153), .Y(n_600) );
INVx2_ASAP7_75t_L g147 ( .A(n_76), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_77), .B(n_234), .Y(n_579) );
INVx1_ASAP7_75t_L g135 ( .A(n_78), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_80), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_81), .B(n_210), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_82), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_84), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_87), .B(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_88), .A2(n_100), .B1(n_178), .B2(n_200), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_89), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_92), .B(n_210), .Y(n_229) );
INVx1_ASAP7_75t_L g115 ( .A(n_93), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_93), .B(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_94), .B(n_190), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_95), .A2(n_159), .B(n_180), .C(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g203 ( .A(n_97), .B(n_204), .Y(n_203) );
NAND2xp33_ASAP7_75t_L g237 ( .A(n_98), .B(n_199), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_99), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_118), .B(n_846), .Y(n_101) );
CKINVDCx12_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx5_ASAP7_75t_L g848 ( .A(n_103), .Y(n_848) );
OR2x6_ASAP7_75t_L g103 ( .A(n_104), .B(n_109), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NOR2x1p5_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g129 ( .A(n_111), .Y(n_129) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_116), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g505 ( .A(n_115), .Y(n_505) );
OR2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_508), .Y(n_118) );
OAI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_123), .B(n_498), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x6_ASAP7_75t_SL g512 ( .A(n_121), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_122), .B(n_503), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_132), .B(n_493), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
CKINVDCx8_ASAP7_75t_R g497 ( .A(n_127), .Y(n_497) );
AND2x6_ASAP7_75t_SL g127 ( .A(n_128), .B(n_130), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_130), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2x1_ASAP7_75t_L g506 ( .A(n_131), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
XNOR2x1_ASAP7_75t_L g133 ( .A(n_134), .B(n_137), .Y(n_133) );
AO22x2_ASAP7_75t_L g516 ( .A1(n_137), .A2(n_517), .B1(n_837), .B2(n_839), .Y(n_516) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_403), .Y(n_137) );
NOR3xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_332), .C(n_374), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_306), .Y(n_139) );
AOI22xp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_205), .B1(n_281), .B2(n_292), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_186), .Y(n_142) );
AOI21xp33_ASAP7_75t_L g325 ( .A1(n_143), .A2(n_326), .B(n_328), .Y(n_325) );
AOI21xp33_ASAP7_75t_L g398 ( .A1(n_143), .A2(n_399), .B(n_400), .Y(n_398) );
OR2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_170), .Y(n_143) );
INVx2_ASAP7_75t_L g318 ( .A(n_144), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_144), .B(n_171), .Y(n_348) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_148), .B(n_154), .C(n_166), .Y(n_145) );
INVx6_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_146), .A2(n_237), .B(n_238), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_146), .B(n_148), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_146), .A2(n_252), .B1(n_528), .B2(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_146), .A2(n_587), .B(n_588), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_146), .A2(n_176), .B1(n_606), .B2(n_607), .Y(n_605) );
BUFx8_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g157 ( .A(n_147), .Y(n_157) );
INVx1_ASAP7_75t_L g180 ( .A(n_147), .Y(n_180) );
INVx1_ASAP7_75t_L g217 ( .A(n_147), .Y(n_217) );
INVxp67_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g544 ( .A(n_150), .Y(n_544) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g153 ( .A(n_151), .Y(n_153) );
INVx1_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
INVx1_ASAP7_75t_L g161 ( .A(n_151), .Y(n_161) );
INVx3_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_151), .Y(n_178) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_151), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_151), .Y(n_200) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_151), .Y(n_222) );
INVx1_ASAP7_75t_L g250 ( .A(n_151), .Y(n_250) );
INVx2_ASAP7_75t_L g256 ( .A(n_151), .Y(n_256) );
OAI21xp33_ASAP7_75t_SL g213 ( .A1(n_152), .A2(n_214), .B(n_215), .Y(n_213) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_153), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g289 ( .A(n_154), .Y(n_289) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_158), .B(n_162), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_155), .A2(n_220), .B(n_221), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g260 ( .A1(n_155), .A2(n_176), .B1(n_261), .B2(n_262), .Y(n_260) );
AOI21x1_ASAP7_75t_L g536 ( .A1(n_155), .A2(n_537), .B(n_539), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_155), .A2(n_176), .B1(n_565), .B2(n_567), .Y(n_564) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g235 ( .A(n_157), .Y(n_235) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_161), .B(n_195), .Y(n_194) );
OAI21xp33_ASAP7_75t_L g166 ( .A1(n_162), .A2(n_163), .B(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g181 ( .A(n_163), .Y(n_181) );
INVx2_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
INVx2_ASAP7_75t_L g191 ( .A(n_163), .Y(n_191) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_164), .Y(n_211) );
INVx1_ASAP7_75t_L g291 ( .A(n_166), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_167), .A2(n_246), .B(n_253), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_167), .A2(n_550), .B(n_555), .Y(n_549) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx10_ASAP7_75t_L g182 ( .A(n_168), .Y(n_182) );
BUFx10_ASAP7_75t_L g224 ( .A(n_168), .Y(n_224) );
INVx1_ASAP7_75t_L g276 ( .A(n_168), .Y(n_276) );
AO31x2_ASAP7_75t_L g562 ( .A1(n_168), .A2(n_563), .A3(n_564), .B(n_568), .Y(n_562) );
AND2x2_ASAP7_75t_L g388 ( .A(n_170), .B(n_227), .Y(n_388) );
INVx1_ASAP7_75t_L g421 ( .A(n_170), .Y(n_421) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g283 ( .A(n_171), .B(n_228), .Y(n_283) );
AND2x2_ASAP7_75t_L g314 ( .A(n_171), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g323 ( .A(n_171), .Y(n_323) );
OR2x2_ASAP7_75t_L g342 ( .A(n_171), .B(n_188), .Y(n_342) );
AND2x2_ASAP7_75t_L g357 ( .A(n_171), .B(n_188), .Y(n_357) );
AO31x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_181), .A3(n_182), .B(n_183), .Y(n_171) );
OAI22x1_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_176), .B1(n_177), .B2(n_179), .Y(n_172) );
INVx4_ASAP7_75t_L g175 ( .A(n_174), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_175), .A2(n_232), .B(n_233), .C(n_234), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_176), .A2(n_179), .B1(n_270), .B2(n_272), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_176), .A2(n_542), .B(n_543), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_176), .A2(n_598), .B1(n_599), .B2(n_600), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_178), .B(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g273 ( .A(n_178), .Y(n_273) );
INVx2_ASAP7_75t_L g540 ( .A(n_178), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_179), .B(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g554 ( .A(n_180), .Y(n_554) );
INVx1_ASAP7_75t_SL g599 ( .A(n_180), .Y(n_599) );
INVx2_ASAP7_75t_L g584 ( .A(n_181), .Y(n_584) );
INVx2_ASAP7_75t_L g202 ( .A(n_182), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
INVx2_ASAP7_75t_L g204 ( .A(n_185), .Y(n_204) );
BUFx2_ASAP7_75t_L g244 ( .A(n_185), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_185), .B(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_185), .B(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_185), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_187), .B(n_356), .Y(n_399) );
OR2x2_ASAP7_75t_L g487 ( .A(n_187), .B(n_348), .Y(n_487) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g315 ( .A(n_188), .Y(n_315) );
AND2x2_ASAP7_75t_L g324 ( .A(n_188), .B(n_287), .Y(n_324) );
AND2x2_ASAP7_75t_L g327 ( .A(n_188), .B(n_228), .Y(n_327) );
AND2x2_ASAP7_75t_L g346 ( .A(n_188), .B(n_227), .Y(n_346) );
AND2x4_ASAP7_75t_L g365 ( .A(n_188), .B(n_288), .Y(n_365) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_192), .B(n_203), .Y(n_188) );
AOI21x1_ASAP7_75t_L g548 ( .A1(n_189), .A2(n_549), .B(n_558), .Y(n_548) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_196), .B(n_202), .Y(n_192) );
OAI22xp33_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B1(n_200), .B2(n_201), .Y(n_197) );
INVx2_ASAP7_75t_L g271 ( .A(n_199), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_200), .A2(n_222), .B1(n_552), .B2(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g580 ( .A(n_200), .Y(n_580) );
OAI21xp33_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_225), .B(n_266), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_206), .B(n_360), .Y(n_463) );
CKINVDCx14_ASAP7_75t_R g206 ( .A(n_207), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_208), .B(n_280), .Y(n_279) );
INVx3_ASAP7_75t_L g296 ( .A(n_208), .Y(n_296) );
OR2x2_ASAP7_75t_L g304 ( .A(n_208), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_208), .B(n_297), .Y(n_329) );
AND2x2_ASAP7_75t_L g354 ( .A(n_208), .B(n_268), .Y(n_354) );
AND2x2_ASAP7_75t_L g372 ( .A(n_208), .B(n_302), .Y(n_372) );
INVx1_ASAP7_75t_L g411 ( .A(n_208), .Y(n_411) );
AND2x2_ASAP7_75t_L g413 ( .A(n_208), .B(n_414), .Y(n_413) );
NAND2x1p5_ASAP7_75t_SL g432 ( .A(n_208), .B(n_353), .Y(n_432) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_212), .Y(n_208) );
NOR2x1_ASAP7_75t_L g239 ( .A(n_210), .B(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g263 ( .A(n_210), .Y(n_263) );
INVx4_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g223 ( .A(n_211), .B(n_224), .Y(n_223) );
INVx2_ASAP7_75t_SL g534 ( .A(n_211), .Y(n_534) );
BUFx3_ASAP7_75t_L g563 ( .A(n_211), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_211), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g573 ( .A(n_211), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_211), .B(n_609), .Y(n_608) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_219), .B(n_223), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
BUFx4f_ASAP7_75t_L g252 ( .A(n_217), .Y(n_252) );
INVx1_ASAP7_75t_L g591 ( .A(n_217), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_222), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g566 ( .A(n_222), .Y(n_566) );
INVx1_ASAP7_75t_L g240 ( .A(n_224), .Y(n_240) );
AO31x2_ASAP7_75t_L g259 ( .A1(n_224), .A2(n_260), .A3(n_263), .B(n_264), .Y(n_259) );
OAI21x1_ASAP7_75t_L g574 ( .A1(n_224), .A2(n_575), .B(n_578), .Y(n_574) );
OAI21x1_ASAP7_75t_L g585 ( .A1(n_224), .A2(n_586), .B(n_589), .Y(n_585) );
AOI31xp67_ASAP7_75t_L g604 ( .A1(n_224), .A2(n_263), .A3(n_605), .B(n_608), .Y(n_604) );
OAI32xp33_ASAP7_75t_L g316 ( .A1(n_225), .A2(n_308), .A3(n_317), .B1(n_319), .B2(n_321), .Y(n_316) );
OR2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_241), .Y(n_225) );
INVx1_ASAP7_75t_L g356 ( .A(n_226), .Y(n_356) );
AND2x2_ASAP7_75t_L g364 ( .A(n_226), .B(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g363 ( .A(n_227), .B(n_287), .Y(n_363) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
BUFx3_ASAP7_75t_L g313 ( .A(n_228), .Y(n_313) );
AND2x2_ASAP7_75t_L g322 ( .A(n_228), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g428 ( .A(n_228), .Y(n_428) );
NAND2x1p5_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
OAI21x1_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_236), .B(n_239), .Y(n_230) );
INVx2_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_235), .A2(n_579), .B1(n_580), .B2(n_581), .Y(n_578) );
INVx2_ASAP7_75t_L g298 ( .A(n_241), .Y(n_298) );
OR2x2_ASAP7_75t_L g308 ( .A(n_241), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g430 ( .A(n_241), .Y(n_430) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_258), .Y(n_241) );
AND2x2_ASAP7_75t_L g331 ( .A(n_242), .B(n_259), .Y(n_331) );
INVx2_ASAP7_75t_L g353 ( .A(n_242), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_242), .B(n_268), .Y(n_373) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g280 ( .A(n_243), .Y(n_280) );
AOI21x1_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_257), .Y(n_243) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_244), .A2(n_269), .A3(n_275), .B(n_277), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_249), .B(n_252), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx2_ASAP7_75t_L g274 ( .A(n_250), .Y(n_274) );
O2A1O1Ixp5_ASAP7_75t_L g575 ( .A1(n_252), .A2(n_274), .B(n_576), .C(n_577), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx2_ASAP7_75t_SL g538 ( .A(n_256), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_258), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g362 ( .A(n_258), .Y(n_362) );
INVx2_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
BUFx2_ASAP7_75t_L g302 ( .A(n_259), .Y(n_302) );
OR2x2_ASAP7_75t_L g368 ( .A(n_259), .B(n_268), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_259), .B(n_268), .Y(n_401) );
INVx2_ASAP7_75t_L g349 ( .A(n_266), .Y(n_349) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_279), .Y(n_266) );
OR2x2_ASAP7_75t_L g336 ( .A(n_267), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g414 ( .A(n_267), .Y(n_414) );
INVx1_ASAP7_75t_L g297 ( .A(n_268), .Y(n_297) );
INVx1_ASAP7_75t_L g305 ( .A(n_268), .Y(n_305) );
INVx1_ASAP7_75t_L g320 ( .A(n_268), .Y(n_320) );
AO31x2_ASAP7_75t_L g596 ( .A1(n_275), .A2(n_563), .A3(n_597), .B(n_601), .Y(n_596) );
INVx2_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_SL g530 ( .A(n_276), .Y(n_530) );
OR2x2_ASAP7_75t_L g424 ( .A(n_279), .B(n_401), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_280), .B(n_296), .Y(n_337) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_280), .Y(n_339) );
OR2x2_ASAP7_75t_L g438 ( .A(n_280), .B(n_362), .Y(n_438) );
INVxp67_ASAP7_75t_L g462 ( .A(n_280), .Y(n_462) );
INVx2_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
NAND2x1_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_283), .B(n_324), .Y(n_391) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g340 ( .A(n_285), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g453 ( .A(n_286), .Y(n_453) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g482 ( .A(n_287), .B(n_315), .Y(n_482) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g408 ( .A(n_288), .B(n_315), .Y(n_408) );
AOI21x1_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_290), .B(n_291), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_299), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_295), .B(n_331), .Y(n_445) );
AND2x4_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx2_ASAP7_75t_L g309 ( .A(n_296), .Y(n_309) );
AND2x2_ASAP7_75t_L g359 ( .A(n_296), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_296), .B(n_353), .Y(n_402) );
OR2x2_ASAP7_75t_L g474 ( .A(n_296), .B(n_361), .Y(n_474) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g394 ( .A(n_300), .B(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx2_ASAP7_75t_L g385 ( .A(n_301), .Y(n_385) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g375 ( .A(n_304), .B(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_SL g386 ( .A(n_304), .Y(n_386) );
OR2x2_ASAP7_75t_L g437 ( .A(n_304), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g492 ( .A(n_304), .Y(n_492) );
AOI211xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_310), .B(n_316), .C(n_325), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g381 ( .A(n_309), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_309), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g454 ( .A(n_309), .B(n_331), .Y(n_454) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_312), .B(n_357), .Y(n_379) );
NAND2x1p5_ASAP7_75t_L g396 ( .A(n_312), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g464 ( .A(n_312), .B(n_465), .Y(n_464) );
INVx3_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx2_ASAP7_75t_L g407 ( .A(n_313), .Y(n_407) );
AND2x2_ASAP7_75t_L g435 ( .A(n_314), .B(n_363), .Y(n_435) );
INVx2_ASAP7_75t_L g458 ( .A(n_314), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_314), .B(n_356), .Y(n_490) );
AND2x4_ASAP7_75t_SL g444 ( .A(n_317), .B(n_322), .Y(n_444) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g397 ( .A(n_318), .B(n_323), .Y(n_397) );
OR2x2_ASAP7_75t_L g449 ( .A(n_318), .B(n_342), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_319), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_319), .B(n_331), .Y(n_485) );
BUFx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g433 ( .A(n_320), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g416 ( .A(n_322), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_322), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g466 ( .A(n_323), .Y(n_466) );
BUFx2_ASAP7_75t_L g334 ( .A(n_324), .Y(n_334) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g452 ( .A(n_327), .B(n_453), .Y(n_452) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g376 ( .A(n_331), .Y(n_376) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_331), .Y(n_393) );
NAND3xp33_ASAP7_75t_SL g332 ( .A(n_333), .B(n_343), .C(n_358), .Y(n_332) );
AOI22xp33_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_335), .B1(n_338), .B2(n_340), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_340), .A2(n_366), .B1(n_447), .B2(n_450), .C1(n_452), .C2(n_454), .Y(n_446) );
AND2x2_ASAP7_75t_L g478 ( .A(n_341), .B(n_427), .Y(n_478) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g426 ( .A(n_342), .B(n_427), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_349), .B1(n_350), .B2(n_355), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx2_ASAP7_75t_SL g422 ( .A(n_346), .Y(n_422) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_354), .Y(n_350) );
AND2x2_ASAP7_75t_L g409 ( .A(n_351), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g367 ( .A(n_352), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g361 ( .A(n_353), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g476 ( .A(n_354), .Y(n_476) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_357), .B(n_453), .Y(n_472) );
INVx1_ASAP7_75t_L g489 ( .A(n_357), .Y(n_489) );
AOI222xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_363), .B1(n_364), .B2(n_366), .C1(n_369), .C2(n_370), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_365), .Y(n_369) );
AND2x2_ASAP7_75t_L g387 ( .A(n_365), .B(n_388), .Y(n_387) );
INVx3_ASAP7_75t_L g418 ( .A(n_365), .Y(n_418) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g382 ( .A(n_368), .Y(n_382) );
OR2x2_ASAP7_75t_L g451 ( .A(n_368), .B(n_432), .Y(n_451) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
OAI211xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_377), .B(n_380), .C(n_389), .Y(n_374) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI21xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_383), .B(n_387), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_381), .A2(n_419), .B1(n_468), .B2(n_471), .C(n_473), .Y(n_467) );
AND2x4_ASAP7_75t_L g410 ( .A(n_382), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g441 ( .A(n_388), .Y(n_441) );
AOI211x1_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B(n_394), .C(n_398), .Y(n_389) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g459 ( .A(n_397), .Y(n_459) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_400), .B(n_448), .C(n_449), .Y(n_447) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g483 ( .A(n_401), .Y(n_483) );
NOR2x1_ASAP7_75t_L g403 ( .A(n_404), .B(n_455), .Y(n_403) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_405), .B(n_412), .C(n_434), .D(n_446), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_409), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
AND2x2_ASAP7_75t_L g465 ( .A(n_408), .B(n_466), .Y(n_465) );
AOI221x1_ASAP7_75t_L g434 ( .A1(n_410), .A2(n_435), .B1(n_436), .B2(n_439), .C(n_442), .Y(n_434) );
AND2x2_ASAP7_75t_L g460 ( .A(n_410), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g470 ( .A(n_411), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B1(n_419), .B2(n_423), .C(n_425), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_417), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_422), .A2(n_426), .B1(n_429), .B2(n_431), .Y(n_425) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_426), .A2(n_443), .B(n_445), .Y(n_442) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g448 ( .A(n_428), .Y(n_448) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g469 ( .A(n_438), .Y(n_469) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_451), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_467), .C(n_479), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_460), .B1(n_463), .B2(n_464), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVxp67_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g475 ( .A(n_462), .B(n_476), .Y(n_475) );
NAND2x1_ASAP7_75t_L g491 ( .A(n_462), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVx2_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_477), .Y(n_473) );
INVx1_ASAP7_75t_SL g477 ( .A(n_478), .Y(n_477) );
AOI221xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_483), .B1(n_484), .B2(n_486), .C(n_488), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx3_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_493), .B(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx4_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
BUFx10_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g838 ( .A(n_505), .Y(n_838) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_505), .Y(n_840) );
INVx1_ASAP7_75t_L g514 ( .A(n_507), .Y(n_514) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_515), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx5_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OAI22xp33_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_841), .B1(n_844), .B2(n_845), .Y(n_515) );
INVx1_ASAP7_75t_L g844 ( .A(n_516), .Y(n_844) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_724), .Y(n_517) );
AND4x1_ASAP7_75t_L g518 ( .A(n_519), .B(n_633), .C(n_671), .D(n_709), .Y(n_518) );
NOR2x1_ASAP7_75t_L g519 ( .A(n_520), .B(n_611), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_559), .B(n_570), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_523), .B(n_531), .Y(n_522) );
NAND2xp5_ASAP7_75t_R g682 ( .A(n_523), .B(n_630), .Y(n_682) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g783 ( .A(n_525), .B(n_661), .Y(n_783) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g561 ( .A(n_526), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g644 ( .A(n_526), .Y(n_644) );
AND2x2_ASAP7_75t_L g658 ( .A(n_526), .B(n_562), .Y(n_658) );
OAI21x1_ASAP7_75t_L g535 ( .A1(n_530), .A2(n_536), .B(n_541), .Y(n_535) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_546), .Y(n_531) );
BUFx2_ASAP7_75t_L g560 ( .A(n_532), .Y(n_560) );
AND2x2_ASAP7_75t_L g616 ( .A(n_532), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g631 ( .A(n_532), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_532), .B(n_562), .Y(n_648) );
INVx3_ASAP7_75t_L g661 ( .A(n_532), .Y(n_661) );
AND2x2_ASAP7_75t_L g696 ( .A(n_532), .B(n_618), .Y(n_696) );
INVx2_ASAP7_75t_L g708 ( .A(n_532), .Y(n_708) );
INVx1_ASAP7_75t_L g712 ( .A(n_532), .Y(n_712) );
INVxp67_ASAP7_75t_L g749 ( .A(n_532), .Y(n_749) );
OR2x2_ASAP7_75t_L g762 ( .A(n_532), .B(n_645), .Y(n_762) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OAI21x1_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B(n_545), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_540), .A2(n_590), .B(n_592), .Y(n_589) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g614 ( .A(n_547), .Y(n_614) );
INVx1_ASAP7_75t_L g701 ( .A(n_547), .Y(n_701) );
AND2x2_ASAP7_75t_L g716 ( .A(n_547), .B(n_562), .Y(n_716) );
INVx1_ASAP7_75t_L g731 ( .A(n_547), .Y(n_731) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g645 ( .A(n_548), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_551), .B(n_554), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_559), .A2(n_820), .B1(n_822), .B2(n_824), .Y(n_819) );
OR2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_560), .B(n_700), .Y(n_777) );
BUFx2_ASAP7_75t_L g791 ( .A(n_560), .Y(n_791) );
AND2x2_ASAP7_75t_L g809 ( .A(n_560), .B(n_665), .Y(n_809) );
INVx2_ASAP7_75t_L g691 ( .A(n_561), .Y(n_691) );
OR2x2_ASAP7_75t_L g707 ( .A(n_561), .B(n_708), .Y(n_707) );
INVx3_ASAP7_75t_L g615 ( .A(n_562), .Y(n_615) );
AND2x2_ASAP7_75t_L g700 ( .A(n_562), .B(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_594), .Y(n_570) );
OR2x2_ASAP7_75t_L g756 ( .A(n_571), .B(n_713), .Y(n_756) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_583), .Y(n_571) );
AND2x2_ASAP7_75t_L g627 ( .A(n_572), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g668 ( .A(n_572), .Y(n_668) );
INVx2_ASAP7_75t_SL g676 ( .A(n_572), .Y(n_676) );
BUFx2_ASAP7_75t_L g688 ( .A(n_572), .Y(n_688) );
OR2x2_ASAP7_75t_L g776 ( .A(n_572), .B(n_596), .Y(n_776) );
OA21x2_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B(n_582), .Y(n_572) );
OA21x2_ASAP7_75t_L g641 ( .A1(n_573), .A2(n_574), .B(n_582), .Y(n_641) );
AND2x2_ASAP7_75t_L g620 ( .A(n_583), .B(n_603), .Y(n_620) );
AND2x2_ASAP7_75t_L g656 ( .A(n_583), .B(n_641), .Y(n_656) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B(n_593), .Y(n_583) );
OAI21x1_ASAP7_75t_L g626 ( .A1(n_584), .A2(n_585), .B(n_593), .Y(n_626) );
INVx1_ASAP7_75t_L g694 ( .A(n_594), .Y(n_694) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_595), .B(n_688), .Y(n_687) );
AND2x4_ASAP7_75t_L g800 ( .A(n_595), .B(n_780), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_595), .B(n_623), .Y(n_824) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_603), .Y(n_595) );
INVx1_ASAP7_75t_L g628 ( .A(n_596), .Y(n_628) );
INVx2_ASAP7_75t_L g638 ( .A(n_596), .Y(n_638) );
AND2x2_ASAP7_75t_L g652 ( .A(n_596), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g667 ( .A(n_596), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g681 ( .A(n_596), .B(n_641), .Y(n_681) );
OR2x2_ASAP7_75t_L g713 ( .A(n_596), .B(n_653), .Y(n_713) );
INVx1_ASAP7_75t_L g797 ( .A(n_596), .Y(n_797) );
AND2x2_ASAP7_75t_L g640 ( .A(n_603), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g678 ( .A(n_603), .Y(n_678) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g654 ( .A(n_604), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g609 ( .A(n_610), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_619), .B1(n_621), .B2(n_629), .Y(n_611) );
NAND2x1p5_ASAP7_75t_L g612 ( .A(n_613), .B(n_616), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g758 ( .A(n_614), .Y(n_758) );
INVx1_ASAP7_75t_L g632 ( .A(n_615), .Y(n_632) );
AND2x4_ASAP7_75t_L g665 ( .A(n_615), .B(n_618), .Y(n_665) );
AND2x2_ASAP7_75t_L g774 ( .A(n_615), .B(n_645), .Y(n_774) );
AND2x2_ASAP7_75t_L g826 ( .A(n_616), .B(n_700), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_616), .B(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g680 ( .A(n_620), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g813 ( .A(n_620), .B(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_627), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_623), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g732 ( .A(n_623), .Y(n_732) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g798 ( .A(n_624), .Y(n_798) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g685 ( .A(n_625), .Y(n_685) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g670 ( .A(n_626), .B(n_654), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_627), .B(n_669), .Y(n_785) );
AND2x2_ASAP7_75t_L g677 ( .A(n_628), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx1_ASAP7_75t_L g817 ( .A(n_632), .Y(n_817) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_642), .B1(n_649), .B2(n_657), .C(n_662), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_639), .Y(n_635) );
AND2x2_ASAP7_75t_L g735 ( .A(n_636), .B(n_656), .Y(n_735) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_637), .B(n_656), .Y(n_704) );
OR2x2_ASAP7_75t_L g719 ( .A(n_637), .B(n_670), .Y(n_719) );
INVx2_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g684 ( .A(n_638), .B(n_685), .Y(n_684) );
INVxp67_ASAP7_75t_L g795 ( .A(n_640), .Y(n_795) );
INVx1_ASAP7_75t_L g755 ( .A(n_641), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_646), .Y(n_642) );
AND2x2_ASAP7_75t_L g815 ( .A(n_643), .B(n_816), .Y(n_815) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
AND2x2_ASAP7_75t_L g769 ( .A(n_644), .B(n_731), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_645), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g690 ( .A(n_645), .Y(n_690) );
INVx1_ASAP7_75t_L g742 ( .A(n_645), .Y(n_742) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI21xp33_ASAP7_75t_L g710 ( .A1(n_650), .A2(n_676), .B(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_655), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g705 ( .A(n_652), .B(n_688), .Y(n_705) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_652), .Y(n_745) );
AND2x2_ASAP7_75t_L g829 ( .A(n_652), .B(n_766), .Y(n_829) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g836 ( .A(n_655), .B(n_753), .Y(n_836) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx2_ASAP7_75t_SL g737 ( .A(n_658), .Y(n_737) );
AND2x2_ASAP7_75t_L g741 ( .A(n_658), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g801 ( .A(n_658), .B(n_661), .Y(n_801) );
AND2x2_ASAP7_75t_L g823 ( .A(n_658), .B(n_748), .Y(n_823) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g720 ( .A(n_661), .B(n_665), .Y(n_720) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
BUFx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x4_ASAP7_75t_L g714 ( .A(n_665), .B(n_690), .Y(n_714) );
AND2x2_ASAP7_75t_L g747 ( .A(n_665), .B(n_748), .Y(n_747) );
INVx3_ASAP7_75t_L g764 ( .A(n_665), .Y(n_764) );
INVx1_ASAP7_75t_L g833 ( .A(n_666), .Y(n_833) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
AND2x4_ASAP7_75t_L g697 ( .A(n_667), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g739 ( .A(n_669), .B(n_688), .Y(n_739) );
AND2x2_ASAP7_75t_L g765 ( .A(n_669), .B(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g775 ( .A(n_670), .B(n_776), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_692), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_679), .B(n_682), .C(n_683), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_675), .B(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_676), .B(n_723), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_676), .B(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_677), .B(n_780), .Y(n_779) );
AND2x2_ASAP7_75t_L g698 ( .A(n_678), .B(n_685), .Y(n_698) );
INVx1_ASAP7_75t_L g753 ( .A(n_678), .Y(n_753) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_686), .B(n_689), .Y(n_683) );
NAND2x1p5_ASAP7_75t_L g754 ( .A(n_685), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g766 ( .A(n_688), .Y(n_766) );
AND2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
AND2x4_ASAP7_75t_L g790 ( .A(n_691), .B(n_758), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_702), .Y(n_692) );
A2O1A1Ixp33_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B(n_697), .C(n_699), .Y(n_693) );
BUFx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g757 ( .A(n_696), .B(n_758), .Y(n_757) );
BUFx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI21xp5_ASAP7_75t_SL g702 ( .A1(n_703), .A2(n_705), .B(n_706), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_708), .Y(n_717) );
OR2x2_ASAP7_75t_L g736 ( .A(n_708), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g818 ( .A(n_708), .Y(n_818) );
AOI222xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_714), .B1(n_715), .B2(n_718), .C1(n_720), .C2(n_721), .Y(n_709) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_711), .B(n_728), .Y(n_727) );
OR2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
NAND2x1p5_ASAP7_75t_L g768 ( .A(n_712), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g723 ( .A(n_713), .Y(n_723) );
INVx1_ASAP7_75t_L g821 ( .A(n_713), .Y(n_821) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_716), .B(n_782), .Y(n_781) );
BUFx2_ASAP7_75t_L g799 ( .A(n_716), .Y(n_799) );
AND2x4_ASAP7_75t_L g806 ( .A(n_716), .B(n_783), .Y(n_806) );
INVx2_ASAP7_75t_L g835 ( .A(n_716), .Y(n_835) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g771 ( .A1(n_719), .A2(n_772), .B1(n_775), .B2(n_777), .Y(n_771) );
AOI211xp5_ASAP7_75t_L g825 ( .A1(n_721), .A2(n_826), .B(n_827), .C(n_831), .Y(n_825) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NOR2xp67_ASAP7_75t_SL g724 ( .A(n_725), .B(n_786), .Y(n_724) );
NAND4xp25_ASAP7_75t_L g725 ( .A(n_726), .B(n_743), .C(n_750), .D(n_770), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_732), .B(n_733), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_736), .B1(n_738), .B2(n_740), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_737), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_738), .B(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g748 ( .A(n_742), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .Y(n_743) );
AND2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_749), .Y(n_746) );
INVx1_ASAP7_75t_L g773 ( .A(n_749), .Y(n_773) );
AOI221xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_757), .B1(n_759), .B2(n_765), .C(n_767), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_756), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_752), .B(n_768), .Y(n_767) );
OR2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
AND2x2_ASAP7_75t_L g805 ( .A(n_753), .B(n_780), .Y(n_805) );
INVx2_ASAP7_75t_L g780 ( .A(n_754), .Y(n_780) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
NAND2x1_ASAP7_75t_SL g760 ( .A(n_761), .B(n_763), .Y(n_760) );
INVx1_ASAP7_75t_L g830 ( .A(n_761), .Y(n_830) );
INVx3_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g832 ( .A(n_769), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_771), .B(n_778), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
INVx1_ASAP7_75t_L g814 ( .A(n_776), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_781), .B1(n_784), .B2(n_785), .Y(n_778) );
AND2x2_ASAP7_75t_L g811 ( .A(n_780), .B(n_797), .Y(n_811) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g792 ( .A(n_785), .Y(n_792) );
NAND3xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_802), .C(n_825), .Y(n_786) );
AOI222xp33_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_792), .B1(n_793), .B2(n_799), .C1(n_800), .C2(n_801), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_789), .B(n_791), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
OR2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
AOI211xp5_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_806), .B(n_807), .C(n_819), .Y(n_802) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_810), .B1(n_812), .B2(n_815), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_818), .Y(n_816) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_828), .B(n_830), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_833), .B1(n_834), .B2(n_836), .Y(n_831) );
INVx4_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_SL g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g845 ( .A(n_841), .Y(n_845) );
NOR2xp33_ASAP7_75t_R g846 ( .A(n_847), .B(n_848), .Y(n_846) );
endmodule