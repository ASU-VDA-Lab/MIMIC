module fake_jpeg_600_n_674 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_674);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_674;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_6),
.B(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_59),
.Y(n_172)
);

INVx2_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_60),
.B(n_121),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_61),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_62),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_65),
.Y(n_231)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_67),
.Y(n_174)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_68),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_69),
.B(n_79),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_70),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_71),
.Y(n_208)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_74),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_47),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_75),
.Y(n_185)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_78),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_8),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_81),
.B(n_88),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_82),
.Y(n_156)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_85),
.B(n_103),
.Y(n_145)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_54),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_92),
.Y(n_140)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_41),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_93),
.Y(n_177)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_94),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_95),
.Y(n_173)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_96),
.Y(n_187)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_98),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_99),
.Y(n_190)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_101),
.Y(n_196)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_24),
.B(n_8),
.Y(n_103)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_38),
.Y(n_104)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_104),
.Y(n_209)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_105),
.Y(n_195)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_22),
.Y(n_106)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_107),
.Y(n_221)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_35),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_113),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_110),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_111),
.Y(n_183)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_33),
.Y(n_112)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_39),
.B(n_7),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_114),
.Y(n_217)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_35),
.Y(n_115)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_53),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_24),
.B(n_15),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_127),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_118),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_41),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_39),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_122),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_55),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_42),
.Y(n_124)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_124),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_126),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_42),
.B(n_7),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_39),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_128),
.Y(n_215)
);

BUFx12_ASAP7_75t_L g129 ( 
.A(n_38),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_129),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_26),
.B(n_40),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_44),
.Y(n_157)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_48),
.Y(n_131)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_131),
.Y(n_201)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_43),
.Y(n_132)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_113),
.A2(n_43),
.B1(n_57),
.B2(n_30),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_139),
.A2(n_179),
.B1(n_177),
.B2(n_228),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_93),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g236 ( 
.A1(n_146),
.A2(n_160),
.B1(n_205),
.B2(n_214),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_107),
.A2(n_55),
.B1(n_43),
.B2(n_23),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_148),
.A2(n_188),
.B1(n_192),
.B2(n_222),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_40),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_153),
.B(n_168),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_157),
.B(n_165),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_83),
.A2(n_23),
.B1(n_25),
.B2(n_30),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_76),
.B(n_48),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_91),
.B(n_44),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_60),
.B(n_56),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_169),
.B(n_171),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_56),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_80),
.A2(n_57),
.B1(n_38),
.B2(n_50),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_26),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_181),
.B(n_202),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_102),
.A2(n_57),
.B1(n_50),
.B2(n_28),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_110),
.A2(n_118),
.B1(n_126),
.B2(n_125),
.Y(n_192)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

INVx4_ASAP7_75t_SL g267 ( 
.A(n_194),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_111),
.B(n_132),
.C(n_119),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_95),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_106),
.B(n_28),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_198),
.B(n_216),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_101),
.B(n_104),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_63),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_207),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_98),
.A2(n_25),
.B1(n_58),
.B2(n_36),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_114),
.B(n_36),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_64),
.A2(n_65),
.B1(n_94),
.B2(n_58),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_129),
.Y(n_250)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_67),
.Y(n_213)
);

INVx4_ASAP7_75t_SL g300 ( 
.A(n_213),
.Y(n_300)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_115),
.A2(n_27),
.B1(n_58),
.B2(n_46),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_120),
.B(n_27),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_84),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_9),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_59),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_68),
.Y(n_223)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_61),
.A2(n_37),
.B1(n_9),
.B2(n_10),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_225),
.B1(n_3),
.B2(n_4),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_62),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_96),
.A2(n_37),
.B(n_10),
.C(n_11),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_226),
.B(n_14),
.Y(n_284)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_77),
.Y(n_227)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

AND2x4_ASAP7_75t_SL g228 ( 
.A(n_70),
.B(n_99),
.Y(n_228)
);

INVx4_ASAP7_75t_SL g310 ( 
.A(n_228),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_71),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_229)
);

OA22x2_ASAP7_75t_L g281 ( 
.A1(n_229),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_155),
.A2(n_73),
.B1(n_78),
.B2(n_74),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_232),
.Y(n_372)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_233),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_149),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_234),
.B(n_244),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_235),
.B(n_250),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_172),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_239),
.Y(n_320)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_240),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_141),
.B(n_0),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_241),
.B(n_246),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_155),
.Y(n_244)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_245),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_145),
.B(n_3),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_247),
.A2(n_253),
.B1(n_305),
.B2(n_313),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_135),
.A2(n_129),
.B1(n_10),
.B2(n_6),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_248),
.A2(n_296),
.B1(n_306),
.B2(n_307),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_152),
.B(n_4),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_251),
.B(n_252),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_136),
.B(n_4),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_148),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_255),
.Y(n_373)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_134),
.Y(n_256)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_256),
.Y(n_317)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_178),
.Y(n_257)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_257),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_173),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_258),
.A2(n_276),
.B1(n_281),
.B2(n_286),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_133),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_259),
.B(n_266),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_183),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_260),
.Y(n_349)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_183),
.Y(n_261)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_261),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_204),
.B(n_5),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_262),
.B(n_264),
.Y(n_332)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_150),
.Y(n_263)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_263),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_140),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_177),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_268),
.B(n_278),
.Y(n_330)
);

O2A1O1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_214),
.A2(n_187),
.B(n_199),
.C(n_164),
.Y(n_269)
);

O2A1O1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_269),
.A2(n_277),
.B(n_294),
.C(n_261),
.Y(n_366)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_174),
.Y(n_270)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_270),
.Y(n_374)
);

INVx8_ASAP7_75t_L g271 ( 
.A(n_172),
.Y(n_271)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_271),
.Y(n_336)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_196),
.Y(n_273)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_273),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_185),
.B(n_12),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_275),
.B(n_288),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_173),
.A2(n_156),
.B1(n_144),
.B2(n_159),
.Y(n_276)
);

INVx6_ASAP7_75t_SL g277 ( 
.A(n_187),
.Y(n_277)
);

BUFx24_ASAP7_75t_L g343 ( 
.A(n_277),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g278 ( 
.A(n_195),
.B(n_12),
.Y(n_278)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_212),
.Y(n_279)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_279),
.Y(n_339)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_184),
.Y(n_280)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_280),
.Y(n_367)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_201),
.Y(n_282)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_282),
.Y(n_333)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_209),
.Y(n_283)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_283),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_284),
.B(n_287),
.Y(n_337)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_180),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_285),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_204),
.A2(n_5),
.B1(n_15),
.B2(n_215),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_209),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_137),
.B(n_15),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_154),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_289),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_161),
.B(n_5),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_303),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_154),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_291),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_160),
.A2(n_146),
.B1(n_231),
.B2(n_163),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_292),
.A2(n_208),
.B(n_206),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_142),
.B(n_158),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_293),
.B(n_294),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_230),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_295),
.B(n_297),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_215),
.A2(n_214),
.B1(n_231),
.B2(n_176),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_219),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_230),
.B(n_162),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_298),
.B(n_299),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_211),
.B(n_163),
.Y(n_299)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_186),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_301),
.B(n_302),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_211),
.B(n_151),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_151),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_180),
.Y(n_304)
);

INVx8_ASAP7_75t_L g345 ( 
.A(n_304),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_192),
.A2(n_225),
.B1(n_222),
.B2(n_229),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_205),
.A2(n_221),
.B1(n_218),
.B2(n_193),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_221),
.A2(n_143),
.B1(n_167),
.B2(n_190),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_217),
.B(n_147),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_308),
.B(n_311),
.Y(n_368)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_175),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_309),
.B(n_314),
.Y(n_334)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_217),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_200),
.Y(n_312)
);

BUFx8_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_L g313 ( 
.A1(n_143),
.A2(n_190),
.B1(n_189),
.B2(n_167),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_189),
.B(n_206),
.Y(n_314)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_147),
.Y(n_315)
);

BUFx8_ASAP7_75t_L g352 ( 
.A(n_315),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_138),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_316),
.B(n_312),
.Y(n_341)
);

OAI21xp33_ASAP7_75t_SL g401 ( 
.A1(n_324),
.A2(n_366),
.B(n_287),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_264),
.A2(n_310),
.B1(n_292),
.B2(n_274),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_328),
.A2(n_350),
.B1(n_351),
.B2(n_357),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_341),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_252),
.B(n_200),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_344),
.B(n_364),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_310),
.A2(n_208),
.B1(n_182),
.B2(n_138),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_250),
.A2(n_182),
.B1(n_170),
.B2(n_166),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_237),
.A2(n_175),
.B1(n_269),
.B2(n_305),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_353),
.A2(n_377),
.B1(n_242),
.B2(n_249),
.Y(n_393)
);

A2O1A1Ixp33_ASAP7_75t_L g355 ( 
.A1(n_241),
.A2(n_272),
.B(n_265),
.C(n_246),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_355),
.B(n_315),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_235),
.A2(n_236),
.B1(n_314),
.B2(n_290),
.Y(n_357)
);

NOR3xp33_ASAP7_75t_SL g360 ( 
.A(n_251),
.B(n_238),
.C(n_243),
.Y(n_360)
);

NAND3xp33_ASAP7_75t_L g423 ( 
.A(n_360),
.B(n_330),
.C(n_364),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_235),
.B(n_254),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_361),
.B(n_370),
.C(n_335),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_262),
.B(n_278),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_236),
.A2(n_253),
.B1(n_262),
.B2(n_263),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_365),
.A2(n_369),
.B1(n_376),
.B2(n_372),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_236),
.A2(n_282),
.B1(n_281),
.B2(n_313),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_256),
.B(n_259),
.C(n_266),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_236),
.A2(n_234),
.B1(n_281),
.B2(n_285),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_281),
.A2(n_280),
.B1(n_301),
.B2(n_257),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_372),
.A2(n_300),
.B1(n_316),
.B2(n_233),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_379),
.Y(n_442)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_331),
.Y(n_380)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_380),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_267),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_381),
.B(n_382),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_356),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_321),
.B(n_303),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_383),
.B(n_385),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_346),
.A2(n_239),
.B1(n_304),
.B2(n_295),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_384),
.A2(n_390),
.B1(n_401),
.B2(n_419),
.Y(n_437)
);

AO21x1_ASAP7_75t_L g385 ( 
.A1(n_332),
.A2(n_297),
.B(n_309),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_331),
.Y(n_386)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_386),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_267),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_387),
.B(n_388),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_300),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_346),
.A2(n_271),
.B1(n_245),
.B2(n_240),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_326),
.A2(n_291),
.B(n_289),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_391),
.A2(n_392),
.B(n_408),
.Y(n_435)
);

NAND2xp33_ASAP7_75t_SL g392 ( 
.A(n_326),
.B(n_273),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_393),
.A2(n_427),
.B1(n_367),
.B2(n_325),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_356),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_394),
.B(n_395),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_283),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_336),
.Y(n_396)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_396),
.Y(n_438)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_336),
.Y(n_397)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_397),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_343),
.Y(n_398)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_398),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_327),
.B(n_242),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_399),
.B(n_406),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_356),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_400),
.B(n_409),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_329),
.Y(n_403)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_403),
.Y(n_452)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_340),
.Y(n_404)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_404),
.Y(n_459)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_333),
.Y(n_405)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_405),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_327),
.B(n_249),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_333),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_407),
.B(n_411),
.Y(n_451)
);

OAI21xp33_ASAP7_75t_SL g408 ( 
.A1(n_326),
.A2(n_311),
.B(n_279),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_340),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_322),
.B(n_270),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_410),
.B(n_412),
.Y(n_447)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_348),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_329),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_413),
.B(n_414),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_322),
.B(n_344),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_334),
.B(n_321),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_415),
.B(n_424),
.Y(n_463)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_334),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_417),
.B(n_418),
.Y(n_457)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_317),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_332),
.A2(n_365),
.B1(n_347),
.B2(n_357),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_359),
.B(n_318),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_420),
.B(n_423),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_332),
.A2(n_361),
.B1(n_377),
.B2(n_369),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_421),
.A2(n_426),
.B1(n_339),
.B2(n_378),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_328),
.B(n_354),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_422),
.B(n_368),
.C(n_337),
.Y(n_431)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_425),
.B(n_355),
.Y(n_429)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_317),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_385),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_428),
.B(n_458),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_429),
.B(n_440),
.C(n_448),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_426),
.A2(n_419),
.B1(n_421),
.B2(n_417),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_430),
.A2(n_444),
.B1(n_445),
.B2(n_427),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_431),
.B(n_345),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_385),
.A2(n_366),
.B(n_324),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_433),
.A2(n_323),
.B(n_352),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_425),
.B(n_362),
.C(n_349),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_416),
.A2(n_358),
.B1(n_337),
.B2(n_341),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_416),
.A2(n_337),
.B1(n_348),
.B2(n_360),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_415),
.B(n_351),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_342),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_450),
.B(n_453),
.C(n_460),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_349),
.C(n_342),
.Y(n_453)
);

O2A1O1Ixp33_ASAP7_75t_L g455 ( 
.A1(n_393),
.A2(n_343),
.B(n_339),
.C(n_323),
.Y(n_455)
);

AO22x2_ASAP7_75t_L g479 ( 
.A1(n_455),
.A2(n_323),
.B1(n_343),
.B2(n_352),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_402),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_389),
.B(n_410),
.C(n_411),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_389),
.A2(n_363),
.B1(n_374),
.B2(n_320),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_461),
.A2(n_384),
.B1(n_390),
.B2(n_405),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_391),
.Y(n_462)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_399),
.Y(n_465)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_465),
.Y(n_486)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_468),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_469),
.A2(n_437),
.B1(n_433),
.B2(n_467),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_470),
.B(n_471),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_457),
.B(n_406),
.Y(n_471)
);

OAI22xp33_ASAP7_75t_SL g472 ( 
.A1(n_437),
.A2(n_402),
.B1(n_400),
.B2(n_394),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_472),
.A2(n_483),
.B1(n_505),
.B2(n_451),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_430),
.A2(n_383),
.B1(n_382),
.B2(n_403),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_473),
.A2(n_484),
.B1(n_489),
.B2(n_501),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_386),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_474),
.B(n_487),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_428),
.A2(n_413),
.B1(n_398),
.B2(n_407),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_475),
.Y(n_525)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_434),
.Y(n_477)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_477),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_462),
.A2(n_392),
.B(n_398),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_478),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_479),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_441),
.A2(n_404),
.B(n_380),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_481),
.B(n_495),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_SL g484 ( 
.A1(n_442),
.A2(n_409),
.B1(n_412),
.B2(n_424),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_447),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_456),
.B(n_418),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_488),
.B(n_492),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_444),
.A2(n_397),
.B1(n_396),
.B2(n_363),
.Y(n_489)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_434),
.Y(n_491)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_491),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_459),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_465),
.B(n_458),
.Y(n_493)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_493),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_447),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_494),
.B(n_500),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_441),
.A2(n_352),
.B(n_378),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_429),
.B(n_325),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_440),
.Y(n_516)
);

INVxp33_ASAP7_75t_L g497 ( 
.A(n_454),
.Y(n_497)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_497),
.Y(n_521)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_436),
.Y(n_498)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_498),
.Y(n_524)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_436),
.Y(n_499)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_499),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_464),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_469),
.A2(n_345),
.B1(n_320),
.B2(n_371),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_502),
.A2(n_503),
.B1(n_443),
.B2(n_452),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_SL g503 ( 
.A1(n_443),
.A2(n_371),
.B1(n_319),
.B2(n_338),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_451),
.A2(n_338),
.B(n_367),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_504),
.B(n_508),
.Y(n_510)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_467),
.Y(n_506)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_506),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_450),
.B(n_319),
.Y(n_507)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_507),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_493),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_509),
.B(n_523),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_514),
.A2(n_494),
.B1(n_489),
.B2(n_470),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_516),
.B(n_518),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_482),
.B(n_431),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_482),
.B(n_453),
.C(n_432),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_519),
.B(n_526),
.C(n_527),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_485),
.B(n_460),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_520),
.B(n_522),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_485),
.B(n_456),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_492),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_463),
.C(n_449),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_496),
.B(n_463),
.C(n_449),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_476),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_528),
.B(n_544),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_507),
.B(n_448),
.C(n_446),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_531),
.B(n_537),
.C(n_504),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_488),
.B(n_466),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_532),
.B(n_534),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_480),
.B(n_445),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_480),
.B(n_446),
.C(n_435),
.Y(n_537)
);

INVxp33_ASAP7_75t_L g571 ( 
.A(n_538),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_473),
.A2(n_435),
.B1(n_452),
.B2(n_455),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_542),
.A2(n_543),
.B1(n_505),
.B2(n_483),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_487),
.A2(n_455),
.B1(n_466),
.B2(n_461),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_500),
.B(n_474),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_530),
.B(n_536),
.Y(n_547)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_547),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_513),
.A2(n_476),
.B(n_495),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_548),
.A2(n_535),
.B(n_530),
.Y(n_585)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_541),
.Y(n_549)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_549),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_550),
.A2(n_574),
.B1(n_540),
.B2(n_525),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_551),
.B(n_553),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_518),
.B(n_478),
.C(n_486),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_552),
.B(n_556),
.C(n_560),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_517),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_555),
.B(n_557),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_520),
.B(n_486),
.C(n_471),
.Y(n_556)
);

AND2x6_ASAP7_75t_L g557 ( 
.A(n_532),
.B(n_501),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_517),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_559),
.B(n_565),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_516),
.B(n_519),
.C(n_522),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_561),
.A2(n_564),
.B1(n_525),
.B2(n_543),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_526),
.B(n_481),
.C(n_499),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_563),
.B(n_566),
.C(n_568),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_514),
.A2(n_502),
.B1(n_490),
.B2(n_506),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_510),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_510),
.B(n_498),
.C(n_491),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_541),
.Y(n_567)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_567),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_527),
.B(n_477),
.C(n_459),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_531),
.B(n_438),
.C(n_439),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_569),
.B(n_576),
.Y(n_581)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_536),
.Y(n_570)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_570),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_521),
.B(n_438),
.Y(n_573)
);

NOR3xp33_ASAP7_75t_L g591 ( 
.A(n_573),
.B(n_575),
.C(n_511),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_533),
.A2(n_515),
.B1(n_542),
.B2(n_512),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_515),
.B(n_439),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_537),
.B(n_490),
.C(n_479),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_578),
.A2(n_593),
.B1(n_479),
.B2(n_558),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_579),
.B(n_585),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_568),
.B(n_545),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_SL g617 ( 
.A(n_583),
.B(n_558),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_553),
.B(n_534),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_584),
.B(n_552),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_588),
.A2(n_598),
.B1(n_599),
.B2(n_600),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_562),
.B(n_539),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_590),
.B(n_556),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_591),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_547),
.B(n_524),
.Y(n_592)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_592),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_574),
.A2(n_535),
.B1(n_533),
.B2(n_538),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_554),
.Y(n_595)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_595),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_555),
.B(n_529),
.Y(n_597)
);

CKINVDCx14_ASAP7_75t_R g621 ( 
.A(n_597),
.Y(n_621)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_559),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_564),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_576),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_571),
.A2(n_479),
.B1(n_550),
.B2(n_548),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_601),
.A2(n_571),
.B1(n_566),
.B2(n_572),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g625 ( 
.A(n_602),
.B(n_586),
.Y(n_625)
);

BUFx24_ASAP7_75t_SL g603 ( 
.A(n_582),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_603),
.B(n_604),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_595),
.B(n_569),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_606),
.B(n_607),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_596),
.B(n_546),
.C(n_560),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_584),
.B(n_563),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g628 ( 
.A(n_609),
.B(n_611),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_SL g611 ( 
.A(n_579),
.B(n_572),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_577),
.B(n_546),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_612),
.B(n_580),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_614),
.A2(n_589),
.B1(n_594),
.B2(n_479),
.Y(n_635)
);

FAx1_ASAP7_75t_SL g616 ( 
.A(n_585),
.B(n_557),
.CI(n_551),
.CON(n_616),
.SN(n_616)
);

FAx1_ASAP7_75t_SL g623 ( 
.A(n_616),
.B(n_577),
.CI(n_596),
.CON(n_623),
.SN(n_623)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_617),
.B(n_618),
.Y(n_636)
);

CKINVDCx16_ASAP7_75t_R g618 ( 
.A(n_597),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_600),
.B(n_565),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_619),
.A2(n_592),
.B(n_594),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_620),
.A2(n_601),
.B1(n_588),
.B2(n_599),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_610),
.A2(n_593),
.B1(n_578),
.B2(n_615),
.Y(n_622)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_622),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_623),
.B(n_634),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_612),
.B(n_581),
.C(n_582),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_624),
.B(n_627),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_625),
.B(n_629),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_626),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_607),
.B(n_586),
.C(n_598),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_608),
.B(n_587),
.C(n_589),
.Y(n_629)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_608),
.B(n_580),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_630),
.B(n_633),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_632),
.B(n_635),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_615),
.B(n_587),
.Y(n_633)
);

XOR2xp5_ASAP7_75t_L g637 ( 
.A(n_602),
.B(n_479),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_637),
.B(n_620),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_624),
.A2(n_613),
.B(n_621),
.Y(n_640)
);

OAI21x1_ASAP7_75t_SL g659 ( 
.A1(n_640),
.A2(n_651),
.B(n_633),
.Y(n_659)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_641),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_627),
.B(n_605),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_644),
.B(n_645),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_631),
.B(n_609),
.C(n_611),
.Y(n_645)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_629),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_649),
.B(n_625),
.Y(n_652)
);

AOI221x1_ASAP7_75t_L g651 ( 
.A1(n_636),
.A2(n_605),
.B1(n_610),
.B2(n_616),
.C(n_635),
.Y(n_651)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_652),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_643),
.B(n_638),
.Y(n_654)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_654),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_SL g655 ( 
.A1(n_639),
.A2(n_623),
.B(n_616),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_SL g661 ( 
.A1(n_655),
.A2(n_660),
.B(n_640),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_646),
.B(n_632),
.Y(n_657)
);

XOR2xp5_ASAP7_75t_L g663 ( 
.A(n_657),
.B(n_658),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_639),
.B(n_630),
.C(n_628),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_659),
.B(n_642),
.C(n_650),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_SL g660 ( 
.A1(n_648),
.A2(n_633),
.B(n_623),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_661),
.B(n_666),
.C(n_646),
.Y(n_669)
);

A2O1A1Ixp33_ASAP7_75t_SL g668 ( 
.A1(n_662),
.A2(n_664),
.B(n_642),
.C(n_663),
.Y(n_668)
);

MAJx2_ASAP7_75t_L g666 ( 
.A(n_653),
.B(n_647),
.C(n_645),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_665),
.A2(n_656),
.B(n_652),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_667),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_668),
.B(n_669),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_671),
.B(n_666),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_672),
.A2(n_670),
.B(n_628),
.Y(n_673)
);

FAx1_ASAP7_75t_SL g674 ( 
.A(n_673),
.B(n_637),
.CI(n_624),
.CON(n_674),
.SN(n_674)
);


endmodule