module fake_jpeg_16023_n_292 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_292);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_292;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_181;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_35),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_36),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_12),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_16),
.Y(n_36)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_13),
.C(n_16),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_15),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_22),
.B1(n_24),
.B2(n_17),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_29),
.B1(n_22),
.B2(n_24),
.Y(n_58)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_60),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_70),
.B1(n_41),
.B2(n_42),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_15),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_65),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_22),
.B1(n_17),
.B2(n_26),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_17),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_40),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_50),
.A2(n_22),
.B1(n_25),
.B2(n_14),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_71),
.A2(n_25),
.B1(n_56),
.B2(n_27),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_46),
.B1(n_42),
.B2(n_37),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_61),
.B1(n_63),
.B2(n_36),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_45),
.B1(n_19),
.B2(n_38),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_76),
.A2(n_82),
.B1(n_15),
.B2(n_20),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_28),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_45),
.B1(n_38),
.B2(n_25),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_20),
.B(n_23),
.Y(n_107)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_90),
.Y(n_106)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_67),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_60),
.B1(n_55),
.B2(n_42),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_94),
.B1(n_97),
.B2(n_99),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_88),
.A2(n_64),
.B1(n_47),
.B2(n_37),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_39),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_107),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_63),
.B(n_47),
.C(n_69),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_100),
.B(n_20),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_47),
.B1(n_55),
.B2(n_61),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_98),
.A2(n_32),
.B(n_34),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_25),
.B(n_14),
.C(n_33),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_48),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_53),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_111),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_85),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_77),
.A2(n_32),
.B1(n_27),
.B2(n_28),
.Y(n_109)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_32),
.B1(n_27),
.B2(n_28),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_48),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_118),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_86),
.B(n_53),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_90),
.B(n_100),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_116),
.Y(n_145)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_74),
.Y(n_121)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_73),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_81),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_102),
.C(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_74),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_126),
.B(n_104),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_142),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_154),
.C(n_114),
.Y(n_162)
);

XOR2x1_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_94),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_141),
.A2(n_144),
.B(n_23),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_97),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_99),
.B1(n_110),
.B2(n_101),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_157),
.B1(n_135),
.B2(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_72),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_100),
.Y(n_152)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_124),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_72),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_83),
.B1(n_78),
.B2(n_73),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_84),
.Y(n_171)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_169),
.C(n_183),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_163),
.A2(n_170),
.B1(n_176),
.B2(n_186),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_159),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_150),
.B(n_148),
.C(n_151),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_156),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_181),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_130),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_178),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_149),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_130),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_117),
.B1(n_133),
.B2(n_128),
.Y(n_170)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_128),
.B(n_119),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_78),
.Y(n_180)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_153),
.B(n_140),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_144),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_89),
.B1(n_84),
.B2(n_23),
.Y(n_186)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_138),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_200),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_SL g191 ( 
.A(n_172),
.B(n_152),
.C(n_145),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_191),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_195),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_180),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_157),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_146),
.C(n_148),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_176),
.C(n_163),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_143),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_89),
.Y(n_219)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

XOR2x1_ASAP7_75t_SL g205 ( 
.A(n_178),
.B(n_150),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_205),
.B(n_170),
.Y(n_211)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_184),
.B1(n_164),
.B2(n_177),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_208),
.A2(n_210),
.B1(n_212),
.B2(n_223),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_207),
.A2(n_164),
.B1(n_174),
.B2(n_167),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_211),
.B(n_224),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_201),
.B1(n_205),
.B2(n_182),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_216),
.C(n_13),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_186),
.B1(n_146),
.B2(n_173),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_195),
.B1(n_193),
.B2(n_9),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_84),
.C(n_48),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_13),
.Y(n_236)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_221),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_189),
.A2(n_14),
.B1(n_9),
.B2(n_11),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_222),
.Y(n_238)
);

XOR2x2_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_13),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_224),
.A2(n_202),
.B1(n_197),
.B2(n_195),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_230),
.A2(n_233),
.B1(n_235),
.B2(n_0),
.Y(n_251)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_232),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_195),
.B(n_193),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_193),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_236),
.B(n_239),
.Y(n_243)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_242),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_217),
.A2(n_10),
.B1(n_11),
.B2(n_4),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_10),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_241),
.C(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_250),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_241),
.A2(n_216),
.B1(n_225),
.B2(n_219),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_245),
.A2(n_255),
.B1(n_230),
.B2(n_238),
.Y(n_256)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_218),
.C(n_223),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_227),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_10),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_254),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_34),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_234),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_256),
.B(n_259),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_236),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_260),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_34),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_227),
.B(n_5),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_264),
.B1(n_243),
.B2(n_251),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_16),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_265),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_3),
.B(n_5),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_33),
.Y(n_265)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_250),
.B1(n_247),
.B2(n_252),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_268),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_33),
.C(n_31),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_274),
.C(n_5),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_258),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_271),
.B(n_273),
.Y(n_277)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_3),
.C(n_5),
.Y(n_274)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_278),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_273),
.B(n_6),
.Y(n_279)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_279),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_275),
.A2(n_8),
.B(n_6),
.Y(n_280)
);

NAND4xp25_ASAP7_75t_SL g283 ( 
.A(n_280),
.B(n_274),
.C(n_272),
.D(n_8),
.Y(n_283)
);

AO21x1_ASAP7_75t_L g285 ( 
.A1(n_283),
.A2(n_269),
.B(n_281),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_285),
.A2(n_286),
.B(n_284),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_277),
.B(n_276),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_287),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_270),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_6),
.B(n_7),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_7),
.C(n_8),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_8),
.Y(n_292)
);


endmodule