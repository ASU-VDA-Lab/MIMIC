module fake_netlist_6_1302_n_434 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_125, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_434);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_434;

wire n_326;
wire n_256;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_148;
wire n_208;
wire n_161;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_392;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_246;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_141;
wire n_383;
wire n_200;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_360;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_397;
wire n_155;
wire n_425;
wire n_218;
wire n_234;
wire n_381;
wire n_236;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_417;
wire n_374;
wire n_366;
wire n_407;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_293;
wire n_334;
wire n_370;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_265;
wire n_260;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_152;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_406;
wire n_204;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_164;
wire n_292;
wire n_307;
wire n_433;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_282;
wire n_211;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_136;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_128;
wire n_241;
wire n_275;
wire n_276;
wire n_221;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_277;
wire n_418;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_328;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_412;
wire n_267;
wire n_339;
wire n_315;
wire n_288;
wire n_427;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_259;
wire n_177;
wire n_391;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g126 ( 
.A(n_22),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_1),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_82),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_120),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_69),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_18),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_63),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_2),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_51),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_16),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g142 ( 
.A(n_40),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

AND2x4_ASAP7_75t_L g144 ( 
.A(n_35),
.B(n_15),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_11),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_45),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_48),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_17),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_33),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_25),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_44),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVxp67_ASAP7_75t_SL g157 ( 
.A(n_38),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

INVxp33_ASAP7_75t_SL g159 ( 
.A(n_122),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

INVxp67_ASAP7_75t_SL g162 ( 
.A(n_99),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_30),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_85),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_62),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_53),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_21),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_26),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_65),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_27),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_36),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_5),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_80),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_57),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_39),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_74),
.Y(n_181)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_72),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_5),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_43),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_1),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_34),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_71),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_94),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_67),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_3),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_9),
.Y(n_192)
);

INVxp33_ASAP7_75t_SL g193 ( 
.A(n_70),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_77),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_91),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_75),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_78),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_114),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_4),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_102),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_0),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_50),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_105),
.Y(n_203)
);

OR2x6_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_128),
.A2(n_137),
.B1(n_201),
.B2(n_199),
.Y(n_206)
);

NAND2xp33_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_0),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_130),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_2),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_140),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_139),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_139),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_139),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_132),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_129),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_173),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_133),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_178),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_127),
.B(n_160),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_134),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_167),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_135),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_138),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_141),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g230 ( 
.A(n_144),
.B(n_12),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_143),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_145),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_136),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_131),
.B(n_3),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_196),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_146),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_167),
.B(n_4),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_147),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_221),
.B(n_159),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_217),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_193),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_157),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_6),
.Y(n_246)
);

AO22x2_ASAP7_75t_L g247 ( 
.A1(n_225),
.A2(n_144),
.B1(n_157),
.B2(n_162),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_213),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

AND2x6_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_197),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_222),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_210),
.B(n_239),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_214),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_215),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_218),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_224),
.B(n_162),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_209),
.B(n_153),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_151),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_153),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_164),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_230),
.A2(n_190),
.B1(n_202),
.B2(n_195),
.Y(n_268)
);

AO22x2_ASAP7_75t_L g269 ( 
.A1(n_238),
.A2(n_156),
.B1(n_171),
.B2(n_172),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_204),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_232),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_204),
.Y(n_274)
);

AO22x2_ASAP7_75t_L g275 ( 
.A1(n_231),
.A2(n_179),
.B1(n_200),
.B2(n_198),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_204),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_230),
.Y(n_278)
);

AND2x4_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_230),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_244),
.B(n_266),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_237),
.Y(n_281)
);

BUFx12f_ASAP7_75t_SL g282 ( 
.A(n_241),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_230),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_233),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_246),
.Y(n_285)
);

AND2x4_ASAP7_75t_SL g286 ( 
.A(n_268),
.B(n_234),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_249),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_247),
.A2(n_206),
.B1(n_216),
.B2(n_207),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_L g289 ( 
.A1(n_245),
.A2(n_174),
.B1(n_148),
.B2(n_203),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_241),
.B(n_216),
.Y(n_290)
);

NAND2x1p5_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_271),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_253),
.Y(n_294)
);

NOR2x2_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_206),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_254),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_251),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_247),
.B(n_142),
.Y(n_299)
);

AO22x1_ASAP7_75t_L g300 ( 
.A1(n_271),
.A2(n_182),
.B1(n_149),
.B2(n_169),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_275),
.Y(n_301)
);

NAND2xp33_ASAP7_75t_L g302 ( 
.A(n_253),
.B(n_197),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_251),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_243),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_245),
.A2(n_263),
.B1(n_269),
.B2(n_240),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_269),
.A2(n_197),
.B1(n_177),
.B2(n_170),
.Y(n_306)
);

AND2x4_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_248),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_263),
.B(n_150),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_253),
.B(n_186),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_265),
.B(n_187),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_253),
.B(n_152),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_267),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_260),
.B(n_154),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_258),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_280),
.A2(n_275),
.B1(n_267),
.B2(n_155),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_242),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_278),
.A2(n_242),
.B(n_270),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

O2A1O1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_305),
.A2(n_273),
.B(n_184),
.C(n_180),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_299),
.A2(n_189),
.B1(n_161),
.B2(n_163),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_278),
.A2(n_272),
.B(n_262),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_315),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_299),
.A2(n_289),
.B1(n_306),
.B2(n_284),
.Y(n_324)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_303),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_285),
.B(n_158),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_165),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_310),
.B(n_166),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_304),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_283),
.A2(n_261),
.B(n_250),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_279),
.A2(n_194),
.B1(n_188),
.B2(n_168),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_297),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_281),
.A2(n_257),
.B(n_251),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_294),
.B(n_13),
.Y(n_337)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_294),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_257),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_282),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_14),
.Y(n_341)
);

NAND3x1_ASAP7_75t_L g342 ( 
.A(n_290),
.B(n_6),
.C(n_7),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_303),
.B(n_19),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_314),
.Y(n_344)
);

BUFx4f_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_301),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_295),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_276),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_307),
.Y(n_349)
);

A2O1A1Ixp33_ASAP7_75t_L g350 ( 
.A1(n_311),
.A2(n_8),
.B(n_10),
.C(n_20),
.Y(n_350)
);

BUFx8_ASAP7_75t_L g351 ( 
.A(n_347),
.Y(n_351)
);

OAI21x1_ASAP7_75t_L g352 ( 
.A1(n_322),
.A2(n_311),
.B(n_313),
.Y(n_352)
);

OAI21x1_ASAP7_75t_L g353 ( 
.A1(n_318),
.A2(n_313),
.B(n_287),
.Y(n_353)
);

AO21x1_ASAP7_75t_L g354 ( 
.A1(n_320),
.A2(n_309),
.B(n_302),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_317),
.B(n_286),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_288),
.Y(n_356)
);

AOI21x1_ASAP7_75t_L g357 ( 
.A1(n_332),
.A2(n_298),
.B(n_296),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_334),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_319),
.Y(n_359)
);

OA21x2_ASAP7_75t_L g360 ( 
.A1(n_341),
.A2(n_293),
.B(n_276),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_346),
.A2(n_307),
.B1(n_300),
.B2(n_10),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

AO21x2_ASAP7_75t_L g363 ( 
.A1(n_336),
.A2(n_125),
.B(n_23),
.Y(n_363)
);

CKINVDCx11_ASAP7_75t_R g364 ( 
.A(n_331),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_324),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_324),
.A2(n_31),
.B(n_32),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_37),
.Y(n_367)
);

OAI21x1_ASAP7_75t_L g368 ( 
.A1(n_343),
.A2(n_339),
.B(n_323),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_327),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_326),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_349),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_325),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_344),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_316),
.A2(n_41),
.B(n_42),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_325),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_325),
.Y(n_376)
);

AOI211xp5_ASAP7_75t_L g377 ( 
.A1(n_356),
.A2(n_329),
.B(n_321),
.C(n_350),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_L g378 ( 
.A1(n_367),
.A2(n_321),
.B1(n_316),
.B2(n_345),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_369),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_374),
.A2(n_337),
.B(n_338),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_355),
.A2(n_333),
.B1(n_340),
.B2(n_342),
.Y(n_381)
);

OAI221xp5_ASAP7_75t_L g382 ( 
.A1(n_361),
.A2(n_355),
.B1(n_367),
.B2(n_366),
.C(n_362),
.Y(n_382)
);

AOI221xp5_ASAP7_75t_SL g383 ( 
.A1(n_361),
.A2(n_345),
.B1(n_337),
.B2(n_338),
.C(n_335),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_358),
.A2(n_335),
.B1(n_46),
.B2(n_47),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_370),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_373),
.A2(n_49),
.B1(n_52),
.B2(n_55),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_58),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_372),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_353),
.A2(n_59),
.B(n_60),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_61),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_364),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_365),
.A2(n_66),
.B(n_68),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_379),
.Y(n_393)
);

INVx5_ASAP7_75t_L g394 ( 
.A(n_388),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_385),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_391),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_375),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_387),
.Y(n_398)
);

AOI221xp5_ASAP7_75t_L g399 ( 
.A1(n_378),
.A2(n_354),
.B1(n_363),
.B2(n_376),
.C(n_372),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_390),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_376),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_383),
.B(n_392),
.Y(n_402)
);

AO31x2_ASAP7_75t_L g403 ( 
.A1(n_380),
.A2(n_368),
.A3(n_360),
.B(n_353),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_398),
.A2(n_384),
.B1(n_351),
.B2(n_389),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_400),
.B(n_363),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_393),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_395),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_401),
.B(n_389),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_397),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_394),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_402),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_394),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_409),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_406),
.B(n_403),
.Y(n_414)
);

OAI211xp5_ASAP7_75t_SL g415 ( 
.A1(n_404),
.A2(n_399),
.B(n_386),
.C(n_396),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_411),
.B(n_403),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_407),
.Y(n_417)
);

NOR2x1_ASAP7_75t_L g418 ( 
.A(n_410),
.B(n_412),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_405),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_403),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_352),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_417),
.B(n_81),
.Y(n_422)
);

AOI211x1_ASAP7_75t_SL g423 ( 
.A1(n_422),
.A2(n_415),
.B(n_419),
.C(n_418),
.Y(n_423)
);

OAI221xp5_ASAP7_75t_SL g424 ( 
.A1(n_423),
.A2(n_421),
.B1(n_416),
.B2(n_419),
.C(n_420),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_424),
.B(n_414),
.Y(n_425)
);

AOI31xp33_ASAP7_75t_L g426 ( 
.A1(n_425),
.A2(n_414),
.A3(n_84),
.B(n_90),
.Y(n_426)
);

NOR3xp33_ASAP7_75t_L g427 ( 
.A(n_426),
.B(n_357),
.C(n_352),
.Y(n_427)
);

OAI211xp5_ASAP7_75t_SL g428 ( 
.A1(n_427),
.A2(n_93),
.B(n_95),
.C(n_96),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_428),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_429),
.A2(n_372),
.B1(n_100),
.B2(n_103),
.Y(n_430)
);

AOI211xp5_ASAP7_75t_L g431 ( 
.A1(n_430),
.A2(n_98),
.B(n_107),
.C(n_108),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_431),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_432),
.A2(n_116),
.B(n_117),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_433),
.A2(n_119),
.B1(n_121),
.B2(n_123),
.Y(n_434)
);


endmodule