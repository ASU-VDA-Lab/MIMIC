module fake_jpeg_7552_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_24),
.B(n_16),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_36),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_39),
.B(n_43),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx9p33_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_27),
.Y(n_73)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_50),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_23),
.B(n_0),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_54),
.B(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_62),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_59),
.B(n_64),
.Y(n_97)
);

AO22x2_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_19),
.B1(n_31),
.B2(n_17),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_60),
.A2(n_29),
.B1(n_22),
.B2(n_34),
.Y(n_107)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_69),
.Y(n_94)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_74),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_77),
.Y(n_109)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_26),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_79),
.B(n_88),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_60),
.A2(n_32),
.B1(n_31),
.B2(n_46),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_81),
.A2(n_90),
.B1(n_95),
.B2(n_96),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_84),
.Y(n_134)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_60),
.A2(n_73),
.B(n_53),
.C(n_67),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_87),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_45),
.C(n_15),
.Y(n_88)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_108),
.Y(n_132)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_51),
.A2(n_32),
.B1(n_49),
.B2(n_35),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_67),
.B(n_47),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_119),
.C(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_66),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_21),
.B1(n_28),
.B2(n_27),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_21),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_14),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_33),
.A3(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_47),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_63),
.A2(n_44),
.B1(n_22),
.B2(n_29),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_33),
.B1(n_17),
.B2(n_30),
.Y(n_135)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_66),
.B(n_33),
.Y(n_114)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_56),
.A2(n_44),
.B1(n_28),
.B2(n_34),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_93),
.B1(n_80),
.B2(n_85),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_68),
.B(n_48),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_26),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_121),
.A2(n_123),
.B1(n_128),
.B2(n_135),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_79),
.B(n_94),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_122),
.A2(n_97),
.B(n_109),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_87),
.A2(n_44),
.B1(n_34),
.B2(n_17),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_1),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_142),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_48),
.C(n_40),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_100),
.C(n_104),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_48),
.B1(n_40),
.B2(n_30),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_139),
.A2(n_105),
.B1(n_90),
.B2(n_95),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_141),
.B(n_151),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_1),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_102),
.Y(n_152)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_152),
.B(n_164),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_92),
.B(n_107),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_153),
.A2(n_160),
.B(n_167),
.Y(n_189)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_157),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_155),
.A2(n_159),
.B1(n_177),
.B2(n_160),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_107),
.B1(n_103),
.B2(n_118),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_156),
.A2(n_171),
.B1(n_178),
.B2(n_142),
.Y(n_194)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_158),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_139),
.A2(n_86),
.B1(n_120),
.B2(n_92),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_121),
.A2(n_86),
.B1(n_108),
.B2(n_117),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_138),
.B(n_124),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_108),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_166),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_123),
.A2(n_113),
.B(n_30),
.C(n_112),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_174),
.B(n_149),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_6),
.C(n_8),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_106),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_128),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_150),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_168),
.A2(n_180),
.B(n_126),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_116),
.B(n_12),
.C(n_14),
.D(n_13),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_141),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_91),
.B1(n_117),
.B2(n_84),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_175),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_132),
.A2(n_91),
.B(n_3),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_111),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_176),
.B(n_181),
.Y(n_215)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_179),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_132),
.A2(n_13),
.B1(n_12),
.B2(n_83),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_1),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_83),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_142),
.Y(n_182)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_130),
.B(n_83),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_184),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_SL g185 ( 
.A(n_172),
.B(n_131),
.C(n_141),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_193),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_137),
.B1(n_151),
.B2(n_147),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_186),
.A2(n_198),
.B1(n_206),
.B2(n_216),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_124),
.B1(n_146),
.B2(n_137),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_188),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_190),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_209),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_194),
.A2(n_199),
.B1(n_208),
.B2(n_204),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_SL g220 ( 
.A(n_195),
.B(n_163),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_153),
.A2(n_146),
.B1(n_125),
.B2(n_148),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_161),
.A2(n_149),
.B1(n_126),
.B2(n_130),
.Y(n_199)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_125),
.B(n_150),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_210),
.B(n_212),
.Y(n_225)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_214),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_205),
.B(n_169),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_159),
.A2(n_129),
.B1(n_4),
.B2(n_5),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_13),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_213),
.C(n_174),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_156),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_163),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_4),
.B(n_6),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_152),
.A2(n_6),
.B(n_7),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_173),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_155),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_175),
.Y(n_218)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_218),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_235),
.B1(n_208),
.B2(n_194),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_165),
.Y(n_221)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_179),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_169),
.Y(n_227)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_233),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_169),
.Y(n_231)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_231),
.Y(n_262)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_201),
.A2(n_168),
.B1(n_154),
.B2(n_180),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_234),
.A2(n_240),
.B1(n_216),
.B2(n_203),
.Y(n_265)
);

O2A1O1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_199),
.A2(n_163),
.B(n_178),
.C(n_170),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_238),
.Y(n_266)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_242),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_192),
.B(n_164),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_192),
.C(n_187),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_166),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_241),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_163),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_244),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_190),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_211),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_SL g270 ( 
.A(n_246),
.B(n_254),
.C(n_255),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_248),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_191),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_189),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_256),
.Y(n_284)
);

NAND3xp33_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_185),
.C(n_193),
.Y(n_254)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_187),
.C(n_212),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_207),
.C(n_195),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_213),
.C(n_201),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_229),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_210),
.Y(n_261)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_223),
.A2(n_203),
.B1(n_211),
.B2(n_209),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_263),
.A2(n_226),
.B1(n_230),
.B2(n_235),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_265),
.A2(n_223),
.B(n_263),
.Y(n_274)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_218),
.Y(n_269)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_224),
.Y(n_271)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_252),
.C(n_247),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_273),
.A2(n_277),
.B(n_278),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_274),
.B(n_265),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_249),
.A2(n_232),
.B1(n_244),
.B2(n_245),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_275),
.A2(n_276),
.B1(n_281),
.B2(n_282),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_219),
.B1(n_240),
.B2(n_224),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_250),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_250),
.A2(n_225),
.B1(n_242),
.B2(n_222),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_246),
.A2(n_225),
.B1(n_237),
.B2(n_233),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_230),
.B1(n_220),
.B2(n_221),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_286),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_285),
.A2(n_236),
.B(n_9),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_258),
.Y(n_286)
);

OAI322xp33_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_251),
.A3(n_255),
.B1(n_253),
.B2(n_262),
.C1(n_259),
.C2(n_256),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_288),
.A2(n_269),
.B(n_284),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_271),
.Y(n_290)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_291),
.B(n_298),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_259),
.B(n_248),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_292),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_293),
.B(n_274),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_266),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_268),
.C(n_279),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_235),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_280),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_232),
.Y(n_298)
);

A2O1A1O1Ixp25_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_261),
.B(n_228),
.C(n_266),
.D(n_205),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_284),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_10),
.B(n_294),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_305),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_296),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_290),
.A2(n_280),
.B1(n_273),
.B2(n_278),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_306),
.A2(n_297),
.B1(n_289),
.B2(n_293),
.Y(n_321)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_307),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_8),
.C(n_9),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_313),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_311),
.A2(n_310),
.B1(n_312),
.B2(n_308),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_10),
.C(n_291),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_319),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_318),
.B(n_320),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_303),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_311),
.A2(n_287),
.B1(n_301),
.B2(n_297),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_307),
.Y(n_325)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_325),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_313),
.C(n_306),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_326),
.B(n_327),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_305),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_322),
.B(n_300),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_328),
.A2(n_322),
.B(n_315),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_316),
.Y(n_329)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_329),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_331),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_334)
);

AO21x1_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_332),
.B(n_330),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_333),
.B(n_289),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_336),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_302),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_299),
.B(n_10),
.Y(n_339)
);


endmodule