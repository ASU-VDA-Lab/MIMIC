module fake_ariane_458_n_1701 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1701);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1701;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_263;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_99),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_126),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_6),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_78),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_12),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_51),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_59),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_0),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_121),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_105),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_45),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_39),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_71),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_72),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_67),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_21),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_5),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_81),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_35),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_44),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_97),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_120),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_64),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_2),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_66),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_54),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_38),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_12),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_98),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_76),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_127),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_122),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_1),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_96),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_31),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_28),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_83),
.Y(n_195)
);

INVxp33_ASAP7_75t_SL g196 ( 
.A(n_48),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_27),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_102),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_62),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_18),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_70),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_68),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_135),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_147),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_111),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_89),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_1),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_24),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_2),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_43),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_137),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_0),
.Y(n_215)
);

BUFx8_ASAP7_75t_SL g216 ( 
.A(n_118),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_44),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_146),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_10),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_117),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_60),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_136),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_133),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_24),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_149),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_140),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_74),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_57),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_16),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_130),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_148),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_15),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_42),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_58),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_37),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_41),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_141),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_92),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_82),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_28),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_80),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_113),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_48),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_123),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_51),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_65),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_26),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_132),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_155),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_41),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_138),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_43),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_104),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_110),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_153),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_22),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_23),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_151),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_91),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_107),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_19),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_100),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_31),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_20),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_33),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_139),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_131),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_10),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_77),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_144),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_106),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_30),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_39),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_103),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_13),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_47),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_79),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_69),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_128),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_87),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_142),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_34),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_40),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_94),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_112),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_73),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_90),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_8),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_88),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_4),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_45),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_108),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_5),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_8),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_49),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_53),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_37),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_20),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_14),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_42),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_63),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_15),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_19),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_55),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_27),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_129),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_85),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_61),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_52),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_124),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_161),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_204),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_216),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_190),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_161),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_160),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_244),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_266),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_161),
.Y(n_319)
);

INVxp33_ASAP7_75t_SL g320 ( 
.A(n_275),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_161),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_250),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_196),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_161),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_186),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_193),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_273),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_225),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_198),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_201),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_273),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_273),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_273),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_163),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_210),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_163),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_264),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_264),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_250),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_213),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_175),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_178),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_182),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_191),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_194),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_212),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_209),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_224),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_217),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_229),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_203),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_203),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_205),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_205),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_221),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_159),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_221),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_226),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_215),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_232),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_235),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_251),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_247),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_251),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_271),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_271),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_256),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_226),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_291),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_240),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_257),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_211),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_243),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_262),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_265),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_268),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_282),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_219),
.Y(n_379)
);

INVxp33_ASAP7_75t_SL g380 ( 
.A(n_159),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_288),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_293),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_311),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_311),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_322),
.B(n_262),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_319),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_315),
.Y(n_387)
);

AND3x2_ASAP7_75t_L g388 ( 
.A(n_379),
.B(n_248),
.C(n_228),
.Y(n_388)
);

AO22x1_ASAP7_75t_L g389 ( 
.A1(n_320),
.A2(n_219),
.B1(n_303),
.B2(n_294),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_357),
.Y(n_390)
);

AND2x2_ASAP7_75t_SL g391 ( 
.A(n_314),
.B(n_286),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_373),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_375),
.A2(n_380),
.B1(n_328),
.B2(n_323),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_312),
.B(n_179),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_315),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_317),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_359),
.B(n_156),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_319),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_321),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_313),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_321),
.Y(n_402)
);

AND2x6_ASAP7_75t_L g403 ( 
.A(n_359),
.B(n_211),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_330),
.A2(n_233),
.B1(n_336),
.B2(n_331),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_373),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_341),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_324),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_324),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_327),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_360),
.B(n_269),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_361),
.A2(n_303),
.B1(n_283),
.B2(n_169),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_371),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_327),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_374),
.B(n_269),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_329),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_329),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_369),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_325),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_316),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_332),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_332),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_347),
.A2(n_236),
.B1(n_283),
.B2(n_177),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_369),
.B(n_297),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_333),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_333),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_346),
.B(n_348),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_373),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_350),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_R g429 ( 
.A(n_318),
.B(n_195),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_334),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_334),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_352),
.Y(n_432)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_373),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_373),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_362),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_364),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_352),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_353),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_340),
.B(n_162),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_353),
.B(n_164),
.Y(n_440)
);

AND2x6_ASAP7_75t_L g441 ( 
.A(n_354),
.B(n_211),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_354),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_370),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_368),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_368),
.B(n_262),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_355),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_355),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_445),
.A2(n_166),
.B1(n_290),
.B2(n_236),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_402),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_402),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_383),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_397),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_417),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_445),
.B(n_372),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_383),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_433),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_385),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_384),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_410),
.B(n_356),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_442),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_413),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_413),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_414),
.B(n_356),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_420),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_442),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_384),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_420),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_424),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_424),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_386),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_387),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_386),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_391),
.A2(n_309),
.B1(n_305),
.B2(n_302),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_385),
.B(n_358),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_403),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_387),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_399),
.Y(n_477)
);

NAND2xp33_ASAP7_75t_L g478 ( 
.A(n_444),
.B(n_157),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_429),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_395),
.B(n_358),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_399),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_403),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_396),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_404),
.B(n_157),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_396),
.Y(n_485)
);

BUFx8_ASAP7_75t_SL g486 ( 
.A(n_418),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_400),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_433),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_400),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_407),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_407),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_404),
.B(n_158),
.Y(n_492)
);

INVxp33_ASAP7_75t_L g493 ( 
.A(n_443),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_442),
.Y(n_494)
);

OAI22xp33_ASAP7_75t_L g495 ( 
.A1(n_411),
.A2(n_299),
.B1(n_298),
.B2(n_185),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_394),
.B(n_158),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_426),
.B(n_363),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_423),
.B(n_372),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_390),
.B(n_406),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_417),
.B(n_363),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_408),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_408),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_412),
.B(n_365),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_417),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_409),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_409),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_415),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_415),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_433),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_403),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_416),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_398),
.B(n_432),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_428),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_391),
.A2(n_169),
.B1(n_299),
.B2(n_298),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_416),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_435),
.Y(n_516)
);

CKINVDCx6p67_ASAP7_75t_R g517 ( 
.A(n_391),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_421),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_436),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_433),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_392),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_421),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_432),
.B(n_365),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_425),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_438),
.B(n_366),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_392),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_442),
.Y(n_527)
);

NOR3xp33_ASAP7_75t_L g528 ( 
.A(n_422),
.B(n_389),
.C(n_401),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_423),
.A2(n_300),
.B1(n_366),
.B2(n_367),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_419),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_425),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_430),
.Y(n_532)
);

AO22x2_ASAP7_75t_L g533 ( 
.A1(n_423),
.A2(n_367),
.B1(n_381),
.B2(n_378),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_430),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_431),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_431),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_437),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_442),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_437),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_422),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_437),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_447),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_447),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_438),
.B(n_376),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_447),
.Y(n_545)
);

NAND3xp33_ASAP7_75t_L g546 ( 
.A(n_447),
.B(n_167),
.C(n_165),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_423),
.B(n_376),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_447),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_392),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_393),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_L g551 ( 
.A(n_441),
.B(n_168),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_392),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_405),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_446),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_446),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_388),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_389),
.A2(n_290),
.B1(n_295),
.B2(n_166),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_440),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_393),
.B(n_342),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_439),
.B(n_377),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_392),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_405),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_405),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_427),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_427),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_427),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_434),
.B(n_168),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_434),
.Y(n_568)
);

NAND3xp33_ASAP7_75t_L g569 ( 
.A(n_434),
.B(n_174),
.C(n_170),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_441),
.Y(n_570)
);

OAI22x1_ASAP7_75t_L g571 ( 
.A1(n_441),
.A2(n_170),
.B1(n_295),
.B2(n_174),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_441),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_441),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_441),
.A2(n_177),
.B1(n_185),
.B2(n_263),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_403),
.A2(n_382),
.B1(n_345),
.B2(n_344),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_441),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_403),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_403),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_403),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_433),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_383),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_391),
.A2(n_343),
.B1(n_349),
.B2(n_351),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_404),
.B(n_171),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_433),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_383),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_426),
.B(n_381),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_383),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_402),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_402),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_433),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_383),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_433),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_L g593 ( 
.A(n_444),
.B(n_171),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_445),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_402),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_594),
.B(n_172),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_451),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_451),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_594),
.B(n_172),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_540),
.A2(n_378),
.B1(n_377),
.B2(n_339),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_455),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_470),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_448),
.A2(n_276),
.B1(n_272),
.B2(n_261),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_453),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_455),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_459),
.B(n_173),
.Y(n_606)
);

BUFx6f_ASAP7_75t_SL g607 ( 
.A(n_556),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_458),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_458),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_558),
.B(n_173),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g611 ( 
.A(n_452),
.B(n_245),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_453),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_448),
.A2(n_252),
.B1(n_310),
.B2(n_308),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_463),
.B(n_181),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_479),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_470),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_472),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_558),
.B(n_181),
.Y(n_618)
);

NAND2x1_ASAP7_75t_L g619 ( 
.A(n_456),
.B(n_488),
.Y(n_619)
);

CKINVDCx16_ASAP7_75t_R g620 ( 
.A(n_513),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_457),
.B(n_183),
.Y(n_621)
);

NAND2x1_ASAP7_75t_L g622 ( 
.A(n_456),
.B(n_211),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_497),
.B(n_183),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_466),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_472),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_457),
.B(n_335),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_486),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_466),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_480),
.B(n_560),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_471),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_471),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_454),
.B(n_335),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_476),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_560),
.B(n_512),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_586),
.B(n_184),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_477),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_454),
.B(n_184),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_586),
.B(n_503),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_476),
.Y(n_639)
);

AND3x1_ASAP7_75t_L g640 ( 
.A(n_528),
.B(n_339),
.C(n_338),
.Y(n_640)
);

NAND2xp33_ASAP7_75t_L g641 ( 
.A(n_456),
.B(n_188),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_483),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_477),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_499),
.B(n_337),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_489),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_481),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_484),
.B(n_188),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_474),
.B(n_189),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_498),
.B(n_189),
.Y(n_649)
);

BUFx5_ASAP7_75t_L g650 ( 
.A(n_577),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_489),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_490),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_490),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_479),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_456),
.A2(n_200),
.B(n_238),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_498),
.B(n_284),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_491),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_481),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_460),
.B(n_284),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_504),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_475),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_491),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_547),
.B(n_285),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_501),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_547),
.B(n_285),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_530),
.Y(n_666)
);

BUFx5_ASAP7_75t_L g667 ( 
.A(n_577),
.Y(n_667)
);

OAI221xp5_ASAP7_75t_L g668 ( 
.A1(n_557),
.A2(n_514),
.B1(n_473),
.B2(n_582),
.C(n_492),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_504),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_554),
.B(n_289),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_514),
.A2(n_289),
.B1(n_310),
.B2(n_308),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_449),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_554),
.B(n_292),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_583),
.B(n_292),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_485),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_555),
.B(n_296),
.Y(n_676)
);

O2A1O1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_555),
.A2(n_338),
.B(n_337),
.C(n_187),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_496),
.B(n_296),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_537),
.A2(n_176),
.B(n_304),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_533),
.B(n_301),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_501),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_449),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_488),
.A2(n_180),
.B(n_197),
.Y(n_683)
);

OR2x6_ASAP7_75t_L g684 ( 
.A(n_556),
.B(n_218),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_460),
.B(n_301),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_488),
.A2(n_223),
.B(n_237),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_537),
.A2(n_287),
.B(n_220),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_475),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_557),
.A2(n_227),
.B(n_234),
.C(n_254),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_559),
.B(n_3),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_460),
.B(n_306),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_450),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_516),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_559),
.B(n_306),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_533),
.B(n_307),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_533),
.B(n_307),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_533),
.B(n_199),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_517),
.B(n_3),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_538),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_544),
.B(n_202),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_539),
.B(n_206),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_SL g702 ( 
.A(n_571),
.B(n_207),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_460),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_L g704 ( 
.A(n_488),
.B(n_192),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_460),
.B(n_192),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_505),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_519),
.B(n_550),
.Y(n_707)
);

NOR2xp67_ASAP7_75t_L g708 ( 
.A(n_569),
.B(n_208),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_465),
.B(n_494),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_505),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_507),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_485),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_539),
.B(n_214),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_507),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_508),
.A2(n_535),
.B1(n_591),
.B2(n_534),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_541),
.B(n_222),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_465),
.B(n_192),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_465),
.B(n_192),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_487),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_509),
.A2(n_281),
.B(n_280),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_538),
.Y(n_721)
);

AND2x6_ASAP7_75t_SL g722 ( 
.A(n_519),
.B(n_4),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_500),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_487),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_478),
.A2(n_279),
.B1(n_278),
.B2(n_277),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_475),
.B(n_6),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_465),
.Y(n_727)
);

NAND3xp33_ASAP7_75t_L g728 ( 
.A(n_593),
.B(n_249),
.C(n_230),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_493),
.B(n_7),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_502),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_465),
.B(n_192),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_508),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_509),
.B(n_7),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_509),
.B(n_9),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_494),
.B(n_192),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_523),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_450),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_494),
.B(n_192),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_511),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_461),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_509),
.B(n_9),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_494),
.B(n_192),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_541),
.B(n_274),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_494),
.B(n_270),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_511),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_517),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_515),
.B(n_231),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_520),
.B(n_11),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_571),
.A2(n_270),
.B1(n_211),
.B2(n_260),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_515),
.Y(n_750)
);

BUFx6f_ASAP7_75t_SL g751 ( 
.A(n_542),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_525),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_565),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_527),
.B(n_270),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_518),
.B(n_267),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_529),
.B(n_574),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_SL g757 ( 
.A1(n_574),
.A2(n_253),
.B1(n_259),
.B2(n_258),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_518),
.B(n_255),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_520),
.B(n_11),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_522),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_522),
.B(n_246),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_520),
.B(n_13),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_527),
.B(n_270),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_527),
.B(n_270),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_531),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_527),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_693),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_602),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_SL g769 ( 
.A1(n_668),
.A2(n_495),
.B1(n_546),
.B2(n_551),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_638),
.B(n_531),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_726),
.B(n_527),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_629),
.B(n_534),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_746),
.B(n_475),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_597),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_634),
.A2(n_592),
.B1(n_520),
.B2(n_590),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_703),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_615),
.Y(n_777)
);

INVx4_ASAP7_75t_L g778 ( 
.A(n_726),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_602),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_635),
.B(n_644),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_615),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_694),
.B(n_580),
.Y(n_782)
);

AND2x2_ASAP7_75t_SL g783 ( 
.A(n_749),
.B(n_482),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_598),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_601),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_620),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_654),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_635),
.B(n_535),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_606),
.B(n_581),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_625),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_756),
.A2(n_749),
.B1(n_690),
.B2(n_694),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_757),
.A2(n_536),
.B1(n_506),
.B2(n_524),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_605),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_661),
.B(n_580),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_614),
.B(n_580),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_608),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_689),
.A2(n_591),
.B(n_581),
.C(n_587),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_703),
.Y(n_798)
);

OAI22x1_ASAP7_75t_L g799 ( 
.A1(n_671),
.A2(n_546),
.B1(n_567),
.B2(n_506),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_609),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_736),
.B(n_585),
.Y(n_801)
);

NAND2x1_ASAP7_75t_L g802 ( 
.A(n_661),
.B(n_580),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_624),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_610),
.B(n_584),
.Y(n_804)
);

OR2x6_ASAP7_75t_L g805 ( 
.A(n_666),
.B(n_482),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_628),
.Y(n_806)
);

AND2x6_ASAP7_75t_SL g807 ( 
.A(n_647),
.B(n_674),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_753),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_626),
.A2(n_536),
.B1(n_532),
.B2(n_524),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_684),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_688),
.B(n_584),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_610),
.B(n_584),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_600),
.B(n_502),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_688),
.B(n_584),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_625),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_752),
.B(n_590),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_636),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_623),
.B(n_585),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_632),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_632),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_630),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_618),
.B(n_587),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_723),
.B(n_590),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_631),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_633),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_639),
.Y(n_826)
);

INVx6_ASAP7_75t_L g827 ( 
.A(n_626),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_621),
.B(n_590),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_684),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_619),
.A2(n_592),
.B(n_548),
.Y(n_830)
);

INVxp67_ASAP7_75t_SL g831 ( 
.A(n_703),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_715),
.B(n_592),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_642),
.A2(n_645),
.B1(n_652),
.B2(n_651),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_707),
.B(n_637),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_703),
.B(n_592),
.Y(n_835)
);

NOR2x2_ASAP7_75t_L g836 ( 
.A(n_684),
.B(n_532),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_621),
.B(n_461),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_648),
.B(n_595),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_647),
.B(n_542),
.Y(n_839)
);

BUFx8_ASAP7_75t_L g840 ( 
.A(n_607),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_674),
.B(n_543),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_640),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_653),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_657),
.B(n_462),
.Y(n_844)
);

INVx5_ASAP7_75t_L g845 ( 
.A(n_766),
.Y(n_845)
);

AO22x1_ASAP7_75t_L g846 ( 
.A1(n_698),
.A2(n_573),
.B1(n_576),
.B2(n_570),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_627),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_596),
.B(n_543),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_672),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_766),
.B(n_548),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_672),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_600),
.B(n_462),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_766),
.B(n_545),
.Y(n_853)
);

NOR2x2_ASAP7_75t_L g854 ( 
.A(n_611),
.B(n_545),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_662),
.B(n_464),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_727),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_682),
.Y(n_857)
);

INVx3_ASAP7_75t_SL g858 ( 
.A(n_729),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_679),
.A2(n_595),
.B1(n_589),
.B2(n_588),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_607),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_664),
.B(n_589),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_682),
.Y(n_862)
);

BUFx12f_ASAP7_75t_L g863 ( 
.A(n_722),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_766),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_649),
.B(n_464),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_727),
.B(n_482),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_687),
.A2(n_588),
.B1(n_469),
.B2(n_468),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_681),
.B(n_469),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_706),
.Y(n_869)
);

INVx4_ASAP7_75t_L g870 ( 
.A(n_751),
.Y(n_870)
);

AOI21xp33_ASAP7_75t_L g871 ( 
.A1(n_678),
.A2(n_613),
.B(n_656),
.Y(n_871)
);

AND2x6_ASAP7_75t_SL g872 ( 
.A(n_678),
.B(n_562),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_710),
.B(n_711),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_663),
.B(n_467),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_714),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_732),
.A2(n_561),
.B1(n_552),
.B2(n_521),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_739),
.B(n_467),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_745),
.B(n_468),
.Y(n_878)
);

INVx5_ASAP7_75t_L g879 ( 
.A(n_699),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_596),
.A2(n_570),
.B1(n_573),
.B2(n_576),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_750),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_692),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_665),
.B(n_575),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_760),
.B(n_765),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_675),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_712),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_599),
.B(n_561),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_689),
.A2(n_562),
.B(n_564),
.C(n_566),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_670),
.B(n_564),
.Y(n_889)
);

INVxp67_ASAP7_75t_SL g890 ( 
.A(n_699),
.Y(n_890)
);

NOR3xp33_ASAP7_75t_L g891 ( 
.A(n_603),
.B(n_552),
.C(n_561),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_719),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_673),
.B(n_566),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_676),
.B(n_561),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_733),
.A2(n_552),
.B(n_521),
.C(n_526),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_604),
.B(n_482),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_700),
.B(n_526),
.Y(n_897)
);

NOR2x1p5_ASAP7_75t_L g898 ( 
.A(n_680),
.B(n_521),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_724),
.A2(n_572),
.B1(n_510),
.B2(n_579),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_721),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_599),
.B(n_521),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_702),
.A2(n_510),
.B1(n_572),
.B2(n_552),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_737),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_660),
.B(n_526),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_733),
.A2(n_734),
.B1(n_762),
.B2(n_748),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_612),
.B(n_510),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_751),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_721),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_730),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_737),
.Y(n_910)
);

CKINVDCx20_ASAP7_75t_R g911 ( 
.A(n_725),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_669),
.B(n_526),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_740),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_740),
.A2(n_510),
.B1(n_578),
.B2(n_579),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_695),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_616),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_617),
.Y(n_917)
);

NOR2xp67_ASAP7_75t_L g918 ( 
.A(n_728),
.B(n_578),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_709),
.Y(n_919)
);

INVx4_ASAP7_75t_L g920 ( 
.A(n_650),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_643),
.Y(n_921)
);

OR2x2_ASAP7_75t_SL g922 ( 
.A(n_696),
.B(n_568),
.Y(n_922)
);

NOR2x1p5_ASAP7_75t_L g923 ( 
.A(n_697),
.B(n_242),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_709),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_747),
.B(n_568),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_646),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_755),
.B(n_563),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_758),
.B(n_563),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_658),
.A2(n_553),
.B1(n_241),
.B2(n_239),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_761),
.B(n_553),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_650),
.Y(n_931)
);

NOR2x2_ASAP7_75t_L g932 ( 
.A(n_708),
.B(n_14),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_734),
.B(n_549),
.Y(n_933)
);

INVxp67_ASAP7_75t_L g934 ( 
.A(n_701),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_650),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_677),
.Y(n_936)
);

NAND2xp33_ASAP7_75t_L g937 ( 
.A(n_650),
.B(n_549),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_650),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_659),
.B(n_685),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_741),
.B(n_549),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_713),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_741),
.B(n_549),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_716),
.B(n_549),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_SL g944 ( 
.A(n_748),
.B(n_16),
.C(n_17),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_743),
.Y(n_945)
);

AND2x6_ASAP7_75t_L g946 ( 
.A(n_759),
.B(n_154),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_759),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_650),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_667),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_762),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_667),
.Y(n_951)
);

NAND2xp33_ASAP7_75t_SL g952 ( 
.A(n_659),
.B(n_17),
.Y(n_952)
);

OA22x2_ASAP7_75t_L g953 ( 
.A1(n_819),
.A2(n_691),
.B1(n_685),
.B2(n_718),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_780),
.B(n_691),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_871),
.A2(n_655),
.B(n_683),
.C(n_686),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_819),
.B(n_18),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_770),
.B(n_667),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_905),
.A2(n_704),
.B(n_641),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_787),
.B(n_667),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_788),
.A2(n_622),
.B(n_731),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_795),
.A2(n_735),
.B(n_705),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_776),
.Y(n_962)
);

AOI221xp5_ASAP7_75t_L g963 ( 
.A1(n_791),
.A2(n_720),
.B1(n_705),
.B2(n_731),
.C(n_717),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_795),
.A2(n_738),
.B(n_717),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_834),
.B(n_667),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_839),
.A2(n_742),
.B(n_718),
.C(n_735),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_772),
.B(n_667),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_813),
.B(n_742),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_820),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_828),
.A2(n_738),
.B(n_763),
.Y(n_970)
);

OAI22x1_ASAP7_75t_L g971 ( 
.A1(n_829),
.A2(n_764),
.B1(n_763),
.B2(n_754),
.Y(n_971)
);

NAND3xp33_ASAP7_75t_SL g972 ( 
.A(n_911),
.B(n_764),
.C(n_754),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_776),
.Y(n_973)
);

INVx5_ASAP7_75t_L g974 ( 
.A(n_773),
.Y(n_974)
);

O2A1O1Ixp5_ASAP7_75t_L g975 ( 
.A1(n_940),
.A2(n_832),
.B(n_950),
.C(n_947),
.Y(n_975)
);

INVx5_ASAP7_75t_L g976 ( 
.A(n_773),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_840),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_937),
.A2(n_942),
.B(n_933),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_895),
.A2(n_744),
.B(n_22),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_842),
.B(n_744),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_786),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_832),
.A2(n_152),
.B(n_150),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_777),
.B(n_778),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_842),
.B(n_21),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_776),
.Y(n_985)
);

INVx4_ASAP7_75t_L g986 ( 
.A(n_778),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_827),
.B(n_23),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_777),
.B(n_25),
.Y(n_988)
);

INVx4_ASAP7_75t_L g989 ( 
.A(n_845),
.Y(n_989)
);

AOI221x1_ASAP7_75t_L g990 ( 
.A1(n_799),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.C(n_30),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_774),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_820),
.B(n_29),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_784),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_839),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_781),
.B(n_32),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_789),
.B(n_35),
.Y(n_996)
);

NAND2x1p5_ASAP7_75t_L g997 ( 
.A(n_866),
.B(n_75),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_810),
.B(n_36),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_808),
.B(n_36),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_818),
.B(n_38),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_791),
.A2(n_40),
.B1(n_46),
.B2(n_47),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_785),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_866),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_841),
.A2(n_46),
.B(n_49),
.C(n_50),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_822),
.B(n_50),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_793),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_776),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_940),
.A2(n_95),
.B(n_56),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_944),
.A2(n_52),
.B(n_84),
.C(n_86),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_845),
.Y(n_1010)
);

AOI22x1_ASAP7_75t_L g1011 ( 
.A1(n_830),
.A2(n_93),
.B1(n_101),
.B2(n_109),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_941),
.B(n_852),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_897),
.A2(n_115),
.B(n_143),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_SL g1014 ( 
.A(n_870),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_786),
.Y(n_1015)
);

INVx6_ASAP7_75t_L g1016 ( 
.A(n_907),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_782),
.B(n_934),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_827),
.B(n_807),
.Y(n_1018)
);

OAI21xp33_ASAP7_75t_SL g1019 ( 
.A1(n_783),
.A2(n_884),
.B(n_873),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_865),
.B(n_874),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_945),
.A2(n_782),
.B(n_801),
.C(n_833),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_796),
.B(n_800),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_829),
.B(n_767),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_803),
.B(n_806),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_816),
.B(n_792),
.Y(n_1025)
);

OR2x6_ASAP7_75t_SL g1026 ( 
.A(n_854),
.B(n_836),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_R g1027 ( 
.A(n_847),
.B(n_767),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_821),
.B(n_824),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_R g1029 ( 
.A(n_907),
.B(n_872),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_858),
.B(n_825),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_845),
.Y(n_1031)
);

NAND2x1p5_ASAP7_75t_L g1032 ( 
.A(n_845),
.B(n_879),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_826),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_798),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_841),
.A2(n_804),
.B(n_812),
.C(n_816),
.Y(n_1035)
);

BUFx12f_ASAP7_75t_L g1036 ( 
.A(n_863),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_858),
.B(n_915),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_769),
.A2(n_809),
.B1(n_843),
.B2(n_869),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_R g1039 ( 
.A(n_952),
.B(n_860),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_875),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_794),
.A2(n_811),
.B(n_814),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_792),
.B(n_823),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_895),
.A2(n_775),
.B(n_797),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_768),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_881),
.Y(n_1045)
);

NAND2xp33_ASAP7_75t_SL g1046 ( 
.A(n_920),
.B(n_802),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_794),
.A2(n_814),
.B(n_811),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_SL g1048 ( 
.A1(n_804),
.A2(n_812),
.B(n_887),
.C(n_901),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_779),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_809),
.B(n_823),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_837),
.A2(n_920),
.B(n_894),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_889),
.A2(n_893),
.B(n_838),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_879),
.B(n_939),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_943),
.A2(n_835),
.B(n_771),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_771),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_798),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_943),
.A2(n_835),
.B(n_890),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_925),
.A2(n_927),
.B(n_928),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_923),
.B(n_805),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_805),
.B(n_883),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_848),
.A2(n_901),
.B(n_887),
.C(n_928),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_925),
.A2(n_930),
.B(n_927),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_805),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_SL g1064 ( 
.A1(n_891),
.A2(n_930),
.B(n_848),
.C(n_912),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_939),
.B(n_885),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_783),
.A2(n_921),
.B1(n_892),
.B2(n_886),
.Y(n_1066)
);

INVx6_ASAP7_75t_L g1067 ( 
.A(n_773),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_900),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_909),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_844),
.A2(n_861),
.B(n_878),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_855),
.A2(n_868),
.B(n_877),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_L g1072 ( 
.A(n_879),
.B(n_856),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_853),
.A2(n_876),
.B(n_951),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_790),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_910),
.B(n_913),
.Y(n_1075)
);

O2A1O1Ixp5_ASAP7_75t_L g1076 ( 
.A1(n_850),
.A2(n_936),
.B(n_853),
.C(n_912),
.Y(n_1076)
);

NOR3xp33_ASAP7_75t_L g1077 ( 
.A(n_850),
.B(n_888),
.C(n_904),
.Y(n_1077)
);

OAI22x1_ASAP7_75t_L g1078 ( 
.A1(n_898),
.A2(n_932),
.B1(n_880),
.B2(n_916),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_900),
.B(n_908),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_908),
.B(n_903),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_919),
.B(n_924),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_931),
.A2(n_949),
.B(n_948),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_879),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_815),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_R g1085 ( 
.A(n_798),
.B(n_864),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_817),
.B(n_882),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_935),
.A2(n_938),
.B(n_831),
.Y(n_1087)
);

NOR3xp33_ASAP7_75t_SL g1088 ( 
.A(n_888),
.B(n_922),
.C(n_946),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_918),
.A2(n_902),
.B(n_919),
.C(n_924),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_917),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_926),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1012),
.B(n_856),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_978),
.A2(n_867),
.B(n_859),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_1027),
.Y(n_1094)
);

NAND2x1_ASAP7_75t_L g1095 ( 
.A(n_989),
.B(n_798),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1012),
.B(n_849),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_991),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_993),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_954),
.A2(n_929),
.B(n_896),
.C(n_906),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1002),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_958),
.A2(n_864),
.B(n_846),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1021),
.B(n_864),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1051),
.A2(n_859),
.B(n_867),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1073),
.A2(n_851),
.B(n_857),
.Y(n_1104)
);

AOI221x1_ASAP7_75t_L g1105 ( 
.A1(n_1038),
.A2(n_924),
.B1(n_919),
.B2(n_862),
.C(n_864),
.Y(n_1105)
);

OR2x6_ASAP7_75t_L g1106 ( 
.A(n_1067),
.B(n_919),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_983),
.B(n_896),
.Y(n_1107)
);

AOI211x1_ASAP7_75t_L g1108 ( 
.A1(n_984),
.A2(n_1022),
.B(n_1028),
.C(n_1024),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1035),
.A2(n_929),
.B1(n_946),
.B2(n_924),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_983),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_1038),
.B(n_906),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1020),
.B(n_946),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1017),
.B(n_946),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_971),
.A2(n_1061),
.A3(n_1052),
.B(n_1062),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_1067),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_967),
.A2(n_914),
.B(n_899),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_1016),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1006),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1001),
.A2(n_1000),
.B1(n_996),
.B2(n_1005),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_967),
.A2(n_957),
.B(n_1058),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1020),
.B(n_969),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1022),
.B(n_1024),
.Y(n_1122)
);

AOI211x1_ASAP7_75t_L g1123 ( 
.A1(n_1028),
.A2(n_995),
.B(n_956),
.C(n_999),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1033),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_1037),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_981),
.B(n_1015),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_957),
.A2(n_1064),
.B(n_1043),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_989),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1043),
.A2(n_955),
.B(n_1071),
.Y(n_1129)
);

NOR2x1_ASAP7_75t_SL g1130 ( 
.A(n_974),
.B(n_976),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1040),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1082),
.A2(n_1054),
.B(n_970),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1070),
.A2(n_961),
.B(n_964),
.Y(n_1133)
);

OA21x2_ASAP7_75t_L g1134 ( 
.A1(n_975),
.A2(n_979),
.B(n_1076),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1023),
.B(n_1065),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1057),
.A2(n_1042),
.B(n_1025),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1045),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1069),
.Y(n_1138)
);

NOR3xp33_ASAP7_75t_L g1139 ( 
.A(n_994),
.B(n_1004),
.C(n_1009),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1090),
.Y(n_1140)
);

AOI221x1_ASAP7_75t_L g1141 ( 
.A1(n_979),
.A2(n_1077),
.B1(n_1078),
.B2(n_972),
.C(n_982),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_996),
.A2(n_1000),
.B(n_1005),
.C(n_1048),
.Y(n_1142)
);

O2A1O1Ixp5_ASAP7_75t_L g1143 ( 
.A1(n_959),
.A2(n_965),
.B(n_966),
.C(n_960),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_SL g1144 ( 
.A1(n_1050),
.A2(n_1089),
.B(n_997),
.Y(n_1144)
);

AOI221xp5_ASAP7_75t_L g1145 ( 
.A1(n_1019),
.A2(n_998),
.B1(n_1018),
.B2(n_1088),
.C(n_1030),
.Y(n_1145)
);

INVxp67_ASAP7_75t_SL g1146 ( 
.A(n_1003),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_962),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1046),
.A2(n_1041),
.B(n_1047),
.Y(n_1148)
);

INVx3_ASAP7_75t_SL g1149 ( 
.A(n_1016),
.Y(n_1149)
);

O2A1O1Ixp5_ASAP7_75t_L g1150 ( 
.A1(n_1008),
.A2(n_1053),
.B(n_1013),
.C(n_987),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_988),
.B(n_992),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1003),
.B(n_980),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1087),
.A2(n_1011),
.B(n_953),
.Y(n_1153)
);

O2A1O1Ixp5_ASAP7_75t_SL g1154 ( 
.A1(n_1063),
.A2(n_1091),
.B(n_968),
.C(n_1075),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_968),
.A2(n_1075),
.B(n_1032),
.Y(n_1155)
);

INVx2_ASAP7_75t_SL g1156 ( 
.A(n_977),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1031),
.Y(n_1157)
);

AOI21xp33_ASAP7_75t_L g1158 ( 
.A1(n_1066),
.A2(n_1055),
.B(n_1060),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1032),
.A2(n_997),
.B(n_1086),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_988),
.B(n_1026),
.Y(n_1160)
);

O2A1O1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1079),
.A2(n_1068),
.B(n_1055),
.C(n_1080),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1081),
.B(n_1084),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_963),
.A2(n_1072),
.B(n_974),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_962),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1044),
.Y(n_1165)
);

NOR4xp25_ASAP7_75t_L g1166 ( 
.A(n_1059),
.B(n_990),
.C(n_1086),
.D(n_1083),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1049),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_L g1168 ( 
.A(n_986),
.B(n_973),
.C(n_1034),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_986),
.B(n_1074),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_973),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1010),
.A2(n_1085),
.B(n_974),
.Y(n_1171)
);

BUFx4_ASAP7_75t_SL g1172 ( 
.A(n_1036),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_974),
.B(n_976),
.Y(n_1173)
);

AND3x2_ASAP7_75t_L g1174 ( 
.A(n_1029),
.B(n_1014),
.C(n_1039),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_976),
.B(n_973),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_985),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_985),
.B(n_1056),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1056),
.B(n_1007),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1007),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1034),
.A2(n_1056),
.B(n_1031),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1010),
.A2(n_978),
.B(n_1051),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1017),
.B(n_452),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_981),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_978),
.A2(n_1051),
.B(n_1073),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1017),
.B(n_452),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_954),
.A2(n_871),
.B(n_780),
.C(n_1058),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_978),
.A2(n_1051),
.B(n_1073),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1012),
.B(n_638),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_969),
.B(n_694),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_971),
.A2(n_905),
.A3(n_895),
.B(n_1061),
.Y(n_1190)
);

INVx1_ASAP7_75t_SL g1191 ( 
.A(n_981),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_958),
.A2(n_905),
.B(n_967),
.Y(n_1192)
);

BUFx8_ASAP7_75t_L g1193 ( 
.A(n_1036),
.Y(n_1193)
);

CKINVDCx11_ASAP7_75t_R g1194 ( 
.A(n_1036),
.Y(n_1194)
);

O2A1O1Ixp5_ASAP7_75t_L g1195 ( 
.A1(n_958),
.A2(n_905),
.B(n_871),
.C(n_780),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_969),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_SL g1197 ( 
.A1(n_1035),
.A2(n_957),
.B(n_1061),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_958),
.A2(n_905),
.B(n_967),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1021),
.B(n_753),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_978),
.A2(n_1051),
.B(n_1073),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_969),
.B(n_519),
.Y(n_1201)
);

AO32x2_ASAP7_75t_L g1202 ( 
.A1(n_1038),
.A2(n_905),
.A3(n_833),
.B1(n_715),
.B2(n_757),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_958),
.A2(n_905),
.B(n_967),
.Y(n_1203)
);

INVx4_ASAP7_75t_L g1204 ( 
.A(n_986),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_969),
.B(n_519),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_991),
.Y(n_1206)
);

AOI221x1_ASAP7_75t_L g1207 ( 
.A1(n_1038),
.A2(n_871),
.B1(n_1004),
.B2(n_994),
.C(n_1058),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_1017),
.B(n_452),
.Y(n_1208)
);

OA21x2_ASAP7_75t_L g1209 ( 
.A1(n_1043),
.A2(n_975),
.B(n_978),
.Y(n_1209)
);

AOI31xp67_ASAP7_75t_L g1210 ( 
.A1(n_953),
.A2(n_940),
.A3(n_1042),
.B(n_1025),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_994),
.A2(n_780),
.B(n_871),
.C(n_638),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_958),
.A2(n_905),
.B(n_967),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_958),
.A2(n_905),
.B(n_967),
.Y(n_1213)
);

AOI21xp33_ASAP7_75t_L g1214 ( 
.A1(n_1038),
.A2(n_905),
.B(n_1019),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_991),
.Y(n_1215)
);

AND2x6_ASAP7_75t_L g1216 ( 
.A(n_1060),
.B(n_1003),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1012),
.B(n_1020),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_969),
.B(n_694),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1027),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_991),
.Y(n_1220)
);

NOR4xp25_ASAP7_75t_L g1221 ( 
.A(n_1001),
.B(n_1004),
.C(n_994),
.D(n_944),
.Y(n_1221)
);

AO21x1_ASAP7_75t_L g1222 ( 
.A1(n_1038),
.A2(n_1062),
.B(n_1058),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1035),
.A2(n_905),
.B(n_1061),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_SL g1224 ( 
.A1(n_979),
.A2(n_1047),
.B(n_1041),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1104),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_1171),
.B(n_1110),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1122),
.B(n_1188),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1184),
.A2(n_1200),
.B(n_1187),
.Y(n_1228)
);

OA21x2_ASAP7_75t_L g1229 ( 
.A1(n_1133),
.A2(n_1129),
.B(n_1105),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1223),
.A2(n_1186),
.B1(n_1199),
.B2(n_1214),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1145),
.A2(n_1182),
.B1(n_1185),
.B2(n_1208),
.Y(n_1231)
);

OAI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1207),
.A2(n_1141),
.B1(n_1109),
.B2(n_1214),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_SL g1233 ( 
.A(n_1193),
.B(n_1174),
.Y(n_1233)
);

NOR2xp33_ASAP7_75t_L g1234 ( 
.A(n_1152),
.B(n_1183),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1098),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1132),
.A2(n_1181),
.B(n_1153),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1189),
.B(n_1218),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1148),
.A2(n_1101),
.B(n_1143),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1103),
.A2(n_1093),
.B(n_1192),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_SL g1240 ( 
.A1(n_1109),
.A2(n_1119),
.B1(n_1223),
.B2(n_1113),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1222),
.B(n_1127),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1119),
.A2(n_1111),
.B1(n_1139),
.B2(n_1217),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1198),
.A2(n_1213),
.B(n_1212),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1211),
.A2(n_1142),
.B(n_1195),
.C(n_1099),
.Y(n_1244)
);

AOI21xp33_ASAP7_75t_L g1245 ( 
.A1(n_1161),
.A2(n_1112),
.B(n_1162),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_SL g1246 ( 
.A(n_1193),
.B(n_1149),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1120),
.A2(n_1203),
.A3(n_1116),
.B(n_1092),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1102),
.A2(n_1221),
.B(n_1197),
.Y(n_1248)
);

CKINVDCx11_ASAP7_75t_R g1249 ( 
.A(n_1194),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1100),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1224),
.A2(n_1136),
.B(n_1150),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1118),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1159),
.A2(n_1163),
.B(n_1155),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_1094),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1209),
.A2(n_1154),
.B(n_1144),
.Y(n_1255)
);

INVx2_ASAP7_75t_SL g1256 ( 
.A(n_1115),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1183),
.B(n_1191),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_SL g1258 ( 
.A1(n_1095),
.A2(n_1092),
.B(n_1217),
.C(n_1177),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1165),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1158),
.A2(n_1201),
.B1(n_1205),
.B2(n_1151),
.Y(n_1260)
);

OAI211xp5_ASAP7_75t_L g1261 ( 
.A1(n_1123),
.A2(n_1166),
.B(n_1221),
.C(n_1108),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1134),
.A2(n_1180),
.B(n_1096),
.Y(n_1262)
);

O2A1O1Ixp33_ASAP7_75t_SL g1263 ( 
.A1(n_1178),
.A2(n_1202),
.B(n_1175),
.C(n_1173),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1219),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1216),
.B(n_1106),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1191),
.A2(n_1126),
.B1(n_1196),
.B2(n_1135),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1124),
.Y(n_1267)
);

AO21x2_ASAP7_75t_L g1268 ( 
.A1(n_1166),
.A2(n_1158),
.B(n_1162),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1115),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1173),
.A2(n_1157),
.B(n_1128),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1168),
.A2(n_1146),
.B(n_1121),
.Y(n_1271)
);

BUFx8_ASAP7_75t_L g1272 ( 
.A(n_1125),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1202),
.A2(n_1220),
.B(n_1215),
.C(n_1206),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1204),
.A2(n_1160),
.B1(n_1107),
.B2(n_1176),
.Y(n_1274)
);

A2O1A1Ixp33_ASAP7_75t_SL g1275 ( 
.A1(n_1128),
.A2(n_1157),
.B(n_1170),
.C(n_1179),
.Y(n_1275)
);

AOI221xp5_ASAP7_75t_L g1276 ( 
.A1(n_1131),
.A2(n_1137),
.B1(n_1138),
.B2(n_1202),
.C(n_1156),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1130),
.A2(n_1168),
.B(n_1169),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_L g1278 ( 
.A(n_1204),
.B(n_1164),
.C(n_1147),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1216),
.B(n_1106),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1117),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1140),
.B(n_1106),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1147),
.A2(n_1164),
.B1(n_1167),
.B2(n_1190),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1114),
.Y(n_1283)
);

OAI211xp5_ASAP7_75t_SL g1284 ( 
.A1(n_1172),
.A2(n_1190),
.B(n_1114),
.C(n_1210),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_R g1285 ( 
.A(n_1216),
.B(n_1147),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1184),
.A2(n_1200),
.B(n_1187),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1097),
.Y(n_1287)
);

AOI221xp5_ASAP7_75t_L g1288 ( 
.A1(n_1119),
.A2(n_540),
.B1(n_668),
.B2(n_1221),
.C(n_871),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_1172),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1184),
.A2(n_1200),
.B(n_1187),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1184),
.A2(n_1200),
.B(n_1187),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1097),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1097),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1097),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1129),
.A2(n_905),
.B(n_1214),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1122),
.B(n_1188),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1189),
.B(n_1218),
.Y(n_1297)
);

OA21x2_ASAP7_75t_L g1298 ( 
.A1(n_1133),
.A2(n_1129),
.B(n_1105),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1176),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1214),
.A2(n_1019),
.B(n_1211),
.C(n_871),
.Y(n_1300)
);

AOI21xp33_ASAP7_75t_L g1301 ( 
.A1(n_1119),
.A2(n_1142),
.B(n_1211),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1122),
.B(n_1188),
.Y(n_1302)
);

AOI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1145),
.A2(n_911),
.B1(n_540),
.B2(n_753),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1184),
.A2(n_1200),
.B(n_1187),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1122),
.B(n_1188),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1223),
.A2(n_780),
.B1(n_1186),
.B2(n_791),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1172),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1176),
.Y(n_1308)
);

BUFx12f_ASAP7_75t_L g1309 ( 
.A(n_1194),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1097),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1184),
.A2(n_1200),
.B(n_1187),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1223),
.A2(n_780),
.B1(n_1186),
.B2(n_791),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1097),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1214),
.A2(n_791),
.B1(n_668),
.B2(n_473),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1196),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1184),
.A2(n_1200),
.B(n_1187),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_1194),
.Y(n_1317)
);

AOI22x1_ASAP7_75t_L g1318 ( 
.A1(n_1223),
.A2(n_452),
.B1(n_1127),
.B2(n_808),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1184),
.A2(n_1200),
.B(n_1187),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1184),
.A2(n_1200),
.B(n_1187),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_SL g1321 ( 
.A1(n_1223),
.A2(n_1186),
.B(n_1214),
.C(n_1035),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1174),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1184),
.A2(n_1200),
.B(n_1187),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1184),
.A2(n_1200),
.B(n_1187),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1097),
.Y(n_1325)
);

AOI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1127),
.A2(n_1148),
.B(n_1102),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1214),
.A2(n_791),
.B1(n_668),
.B2(n_473),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1110),
.Y(n_1328)
);

INVx5_ASAP7_75t_L g1329 ( 
.A(n_1106),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1184),
.A2(n_1200),
.B(n_1187),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1288),
.A2(n_1314),
.B(n_1327),
.C(n_1306),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1231),
.A2(n_1242),
.B1(n_1240),
.B2(n_1314),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_SL g1333 ( 
.A1(n_1312),
.A2(n_1300),
.B(n_1230),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_L g1334 ( 
.A(n_1249),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1227),
.B(n_1296),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1235),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1237),
.B(n_1297),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1250),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1321),
.A2(n_1300),
.B(n_1241),
.Y(n_1339)
);

OA21x2_ASAP7_75t_L g1340 ( 
.A1(n_1243),
.A2(n_1255),
.B(n_1238),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1289),
.Y(n_1341)
);

NOR2xp67_ASAP7_75t_L g1342 ( 
.A(n_1322),
.B(n_1278),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_1289),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1247),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1302),
.B(n_1305),
.Y(n_1345)
);

NOR2xp67_ASAP7_75t_L g1346 ( 
.A(n_1234),
.B(n_1277),
.Y(n_1346)
);

INVxp67_ASAP7_75t_L g1347 ( 
.A(n_1315),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_R g1348 ( 
.A(n_1307),
.B(n_1233),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1242),
.A2(n_1327),
.B1(n_1318),
.B2(n_1248),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1252),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1301),
.A2(n_1244),
.B(n_1261),
.C(n_1284),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1303),
.A2(n_1244),
.B1(n_1232),
.B2(n_1264),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1257),
.B(n_1260),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1267),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1243),
.A2(n_1255),
.B(n_1241),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1269),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1272),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1257),
.B(n_1260),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1287),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1292),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1293),
.Y(n_1361)
);

O2A1O1Ixp5_ASAP7_75t_L g1362 ( 
.A1(n_1326),
.A2(n_1283),
.B(n_1245),
.C(n_1271),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1266),
.B(n_1281),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1247),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1294),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1307),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1254),
.A2(n_1274),
.B1(n_1299),
.B2(n_1308),
.Y(n_1367)
);

AND2x2_ASAP7_75t_SL g1368 ( 
.A(n_1265),
.B(n_1279),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1310),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1321),
.A2(n_1263),
.B(n_1275),
.C(n_1258),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1313),
.B(n_1325),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1273),
.B(n_1259),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1263),
.A2(n_1275),
.B(n_1258),
.C(n_1273),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1276),
.B(n_1269),
.Y(n_1374)
);

AOI21x1_ASAP7_75t_SL g1375 ( 
.A1(n_1251),
.A2(n_1265),
.B(n_1279),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_R g1376 ( 
.A(n_1317),
.B(n_1246),
.Y(n_1376)
);

O2A1O1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1282),
.A2(n_1280),
.B(n_1268),
.C(n_1256),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1228),
.A2(n_1291),
.B(n_1330),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1270),
.Y(n_1379)
);

NAND2xp33_ASAP7_75t_SL g1380 ( 
.A(n_1285),
.B(n_1328),
.Y(n_1380)
);

CKINVDCx6p67_ASAP7_75t_R g1381 ( 
.A(n_1309),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_SL g1382 ( 
.A1(n_1285),
.A2(n_1298),
.B(n_1229),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1283),
.A2(n_1262),
.B(n_1239),
.C(n_1329),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1229),
.A2(n_1298),
.B(n_1226),
.Y(n_1384)
);

CKINVDCx16_ASAP7_75t_R g1385 ( 
.A(n_1309),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1249),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1253),
.B(n_1311),
.Y(n_1387)
);

INVx1_ASAP7_75t_SL g1388 ( 
.A(n_1225),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1236),
.A2(n_1228),
.B(n_1330),
.C(n_1286),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1236),
.A2(n_1304),
.B(n_1286),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_SL g1391 ( 
.A1(n_1290),
.A2(n_1311),
.B(n_1291),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1316),
.B(n_1319),
.Y(n_1392)
);

OR2x2_ASAP7_75t_SL g1393 ( 
.A(n_1320),
.B(n_1323),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1324),
.B(n_1227),
.Y(n_1394)
);

AOI21x1_ASAP7_75t_SL g1395 ( 
.A1(n_1315),
.A2(n_1000),
.B(n_996),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1315),
.B(n_1266),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1237),
.B(n_1297),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1237),
.B(n_1297),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1295),
.A2(n_905),
.B(n_1129),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1376),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1332),
.A2(n_1358),
.B1(n_1353),
.B2(n_1349),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1368),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1344),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1368),
.Y(n_1404)
);

OR2x6_ASAP7_75t_L g1405 ( 
.A(n_1382),
.B(n_1333),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1394),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1347),
.B(n_1346),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1379),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1347),
.B(n_1339),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1364),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1364),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1396),
.B(n_1372),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1336),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1338),
.Y(n_1414)
);

AO21x2_ASAP7_75t_L g1415 ( 
.A1(n_1331),
.A2(n_1399),
.B(n_1383),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1350),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1355),
.B(n_1392),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1354),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1355),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1352),
.B(n_1351),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1340),
.B(n_1371),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1389),
.A2(n_1362),
.B(n_1383),
.Y(n_1422)
);

AO21x2_ASAP7_75t_L g1423 ( 
.A1(n_1331),
.A2(n_1384),
.B(n_1377),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1359),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1360),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1378),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1340),
.B(n_1361),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1378),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1387),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1365),
.B(n_1369),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1378),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1335),
.B(n_1345),
.Y(n_1432)
);

AO21x2_ASAP7_75t_L g1433 ( 
.A1(n_1373),
.A2(n_1374),
.B(n_1390),
.Y(n_1433)
);

OA21x2_ASAP7_75t_L g1434 ( 
.A1(n_1362),
.A2(n_1351),
.B(n_1388),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1363),
.B(n_1397),
.Y(n_1435)
);

OR2x6_ASAP7_75t_L g1436 ( 
.A(n_1370),
.B(n_1391),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1393),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1337),
.B(n_1398),
.Y(n_1438)
);

NOR2x1p5_ASAP7_75t_L g1439 ( 
.A(n_1381),
.B(n_1356),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1426),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1417),
.B(n_1421),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1426),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1427),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1417),
.B(n_1421),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1427),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1406),
.B(n_1367),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1405),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1433),
.Y(n_1448)
);

INVxp67_ASAP7_75t_SL g1449 ( 
.A(n_1419),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1403),
.Y(n_1450)
);

AOI211xp5_ASAP7_75t_L g1451 ( 
.A1(n_1420),
.A2(n_1376),
.B(n_1348),
.C(n_1357),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1420),
.A2(n_1334),
.B1(n_1380),
.B2(n_1342),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1405),
.A2(n_1380),
.B(n_1395),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1408),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1409),
.B(n_1425),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1429),
.B(n_1385),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1403),
.Y(n_1457)
);

NAND2x1p5_ASAP7_75t_L g1458 ( 
.A(n_1422),
.B(n_1434),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1428),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1408),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1429),
.B(n_1375),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1410),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1428),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_L g1464 ( 
.A(n_1448),
.B(n_1401),
.C(n_1409),
.Y(n_1464)
);

AOI33xp33_ASAP7_75t_L g1465 ( 
.A1(n_1441),
.A2(n_1401),
.A3(n_1438),
.B1(n_1437),
.B2(n_1430),
.B3(n_1413),
.Y(n_1465)
);

AOI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1458),
.A2(n_1415),
.B1(n_1423),
.B2(n_1433),
.C(n_1437),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1458),
.A2(n_1448),
.B1(n_1455),
.B2(n_1415),
.C(n_1441),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1454),
.Y(n_1468)
);

AOI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1458),
.A2(n_1415),
.B1(n_1423),
.B2(n_1433),
.C(n_1437),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1455),
.B(n_1407),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1454),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1454),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1441),
.B(n_1438),
.Y(n_1473)
);

NOR4xp25_ASAP7_75t_SL g1474 ( 
.A(n_1449),
.B(n_1400),
.C(n_1410),
.D(n_1411),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1450),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1446),
.B(n_1412),
.Y(n_1476)
);

OAI211xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1446),
.A2(n_1407),
.B(n_1432),
.C(n_1414),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1460),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1461),
.B(n_1447),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1458),
.A2(n_1405),
.B(n_1434),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1446),
.B(n_1438),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1446),
.B(n_1433),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1443),
.B(n_1412),
.Y(n_1483)
);

NOR2x1_ASAP7_75t_L g1484 ( 
.A(n_1453),
.B(n_1405),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1458),
.A2(n_1415),
.B1(n_1423),
.B2(n_1405),
.Y(n_1485)
);

AOI33xp33_ASAP7_75t_L g1486 ( 
.A1(n_1441),
.A2(n_1430),
.A3(n_1416),
.B1(n_1424),
.B2(n_1413),
.B3(n_1418),
.Y(n_1486)
);

AND2x2_ASAP7_75t_SL g1487 ( 
.A(n_1461),
.B(n_1404),
.Y(n_1487)
);

OAI221xp5_ASAP7_75t_L g1488 ( 
.A1(n_1452),
.A2(n_1405),
.B1(n_1434),
.B2(n_1436),
.C(n_1432),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1456),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1440),
.A2(n_1423),
.B(n_1431),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1457),
.Y(n_1491)
);

AO21x2_ASAP7_75t_L g1492 ( 
.A1(n_1442),
.A2(n_1431),
.B(n_1433),
.Y(n_1492)
);

INVx4_ASAP7_75t_L g1493 ( 
.A(n_1456),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1444),
.B(n_1435),
.Y(n_1494)
);

OA21x2_ASAP7_75t_L g1495 ( 
.A1(n_1467),
.A2(n_1442),
.B(n_1463),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1493),
.Y(n_1496)
);

INVx4_ASAP7_75t_SL g1497 ( 
.A(n_1479),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1479),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1493),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1480),
.A2(n_1459),
.B(n_1463),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1468),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1492),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1468),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1473),
.B(n_1444),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1492),
.Y(n_1505)
);

NOR3xp33_ASAP7_75t_L g1506 ( 
.A(n_1464),
.B(n_1453),
.C(n_1451),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1486),
.B(n_1462),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1475),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1471),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1471),
.Y(n_1510)
);

AND2x6_ASAP7_75t_L g1511 ( 
.A(n_1484),
.B(n_1402),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1487),
.B(n_1451),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1472),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1492),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1472),
.Y(n_1515)
);

INVxp67_ASAP7_75t_L g1516 ( 
.A(n_1464),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1478),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1476),
.B(n_1445),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1478),
.Y(n_1519)
);

INVx4_ASAP7_75t_L g1520 ( 
.A(n_1493),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1484),
.A2(n_1459),
.B(n_1463),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1481),
.B(n_1386),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1476),
.Y(n_1523)
);

NAND3xp33_ASAP7_75t_L g1524 ( 
.A(n_1466),
.B(n_1451),
.C(n_1405),
.Y(n_1524)
);

INVx4_ASAP7_75t_SL g1525 ( 
.A(n_1479),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1482),
.B(n_1445),
.Y(n_1526)
);

AND4x1_ASAP7_75t_L g1527 ( 
.A(n_1506),
.B(n_1469),
.C(n_1452),
.D(n_1465),
.Y(n_1527)
);

CKINVDCx20_ASAP7_75t_R g1528 ( 
.A(n_1522),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1497),
.B(n_1525),
.Y(n_1529)
);

NOR3xp33_ASAP7_75t_L g1530 ( 
.A(n_1516),
.B(n_1488),
.C(n_1477),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1501),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1501),
.Y(n_1532)
);

NAND4xp25_ASAP7_75t_L g1533 ( 
.A(n_1506),
.B(n_1485),
.C(n_1493),
.D(n_1461),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1497),
.B(n_1473),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1521),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1516),
.B(n_1470),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1521),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1503),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1497),
.B(n_1494),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1507),
.B(n_1483),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1503),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1507),
.B(n_1523),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1509),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1497),
.B(n_1494),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1508),
.B(n_1444),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1509),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1497),
.B(n_1487),
.Y(n_1547)
);

AOI31xp33_ASAP7_75t_L g1548 ( 
.A1(n_1512),
.A2(n_1524),
.A3(n_1400),
.B(n_1498),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1510),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1525),
.B(n_1487),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1518),
.B(n_1483),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1510),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1525),
.B(n_1479),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1513),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1525),
.B(n_1489),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1513),
.Y(n_1556)
);

INVxp67_ASAP7_75t_L g1557 ( 
.A(n_1496),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1515),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1520),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1515),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1525),
.B(n_1489),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1504),
.B(n_1491),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1504),
.B(n_1491),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1495),
.B(n_1445),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_SL g1565 ( 
.A(n_1524),
.B(n_1456),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1521),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1517),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1535),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1547),
.B(n_1520),
.Y(n_1569)
);

AOI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1548),
.A2(n_1495),
.B(n_1485),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1530),
.B(n_1518),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1531),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1547),
.B(n_1520),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1531),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1529),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1536),
.B(n_1526),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1535),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1550),
.B(n_1520),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1532),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1532),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1538),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1527),
.A2(n_1495),
.B(n_1500),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1538),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1540),
.B(n_1542),
.Y(n_1584)
);

NAND3xp33_ASAP7_75t_L g1585 ( 
.A(n_1527),
.B(n_1495),
.C(n_1499),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1542),
.B(n_1517),
.Y(n_1586)
);

NAND2x1p5_ASAP7_75t_L g1587 ( 
.A(n_1559),
.B(n_1439),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1541),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1557),
.B(n_1519),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1540),
.B(n_1519),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1529),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1537),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1550),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1541),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1543),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1543),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1551),
.B(n_1526),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1546),
.Y(n_1598)
);

NAND2xp33_ASAP7_75t_SL g1599 ( 
.A(n_1528),
.B(n_1496),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1546),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1549),
.Y(n_1601)
);

INVxp33_ASAP7_75t_L g1602 ( 
.A(n_1565),
.Y(n_1602)
);

CKINVDCx16_ASAP7_75t_R g1603 ( 
.A(n_1599),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1571),
.B(n_1551),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1599),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1587),
.B(n_1539),
.Y(n_1606)
);

BUFx3_ASAP7_75t_L g1607 ( 
.A(n_1575),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1593),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1584),
.B(n_1562),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1587),
.B(n_1539),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1600),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1584),
.B(n_1563),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1576),
.B(n_1533),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1593),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1602),
.A2(n_1498),
.B1(n_1544),
.B2(n_1534),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1580),
.Y(n_1616)
);

NOR2x1_ASAP7_75t_L g1617 ( 
.A(n_1585),
.B(n_1559),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1575),
.B(n_1341),
.Y(n_1618)
);

CKINVDCx16_ASAP7_75t_R g1619 ( 
.A(n_1591),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1582),
.A2(n_1415),
.B1(n_1564),
.B2(n_1434),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1580),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1581),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1591),
.Y(n_1623)
);

CKINVDCx14_ASAP7_75t_R g1624 ( 
.A(n_1593),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1587),
.B(n_1544),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1602),
.A2(n_1511),
.B1(n_1490),
.B2(n_1434),
.Y(n_1626)
);

INVxp67_ASAP7_75t_L g1627 ( 
.A(n_1589),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1617),
.A2(n_1570),
.B(n_1586),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1614),
.Y(n_1629)
);

OAI322xp33_ASAP7_75t_L g1630 ( 
.A1(n_1613),
.A2(n_1590),
.A3(n_1576),
.B1(n_1601),
.B2(n_1581),
.C1(n_1597),
.C2(n_1594),
.Y(n_1630)
);

AOI211xp5_ASAP7_75t_L g1631 ( 
.A1(n_1613),
.A2(n_1573),
.B(n_1578),
.C(n_1569),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1604),
.B(n_1597),
.Y(n_1632)
);

OAI21xp33_ASAP7_75t_L g1633 ( 
.A1(n_1605),
.A2(n_1573),
.B(n_1569),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1616),
.Y(n_1634)
);

INVx1_ASAP7_75t_SL g1635 ( 
.A(n_1603),
.Y(n_1635)
);

A2O1A1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1626),
.A2(n_1620),
.B(n_1627),
.C(n_1624),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1619),
.B(n_1603),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1611),
.B(n_1572),
.Y(n_1638)
);

OAI211xp5_ASAP7_75t_SL g1639 ( 
.A1(n_1623),
.A2(n_1559),
.B(n_1601),
.C(n_1596),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1616),
.Y(n_1640)
);

AOI32xp33_ASAP7_75t_L g1641 ( 
.A1(n_1615),
.A2(n_1578),
.A3(n_1566),
.B1(n_1537),
.B2(n_1588),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1621),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1619),
.A2(n_1474),
.B1(n_1436),
.B2(n_1498),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1621),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1606),
.B(n_1553),
.Y(n_1645)
);

OAI22xp5_ASAP7_75t_SL g1646 ( 
.A1(n_1611),
.A2(n_1343),
.B1(n_1366),
.B2(n_1598),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1629),
.Y(n_1647)
);

NAND2x1p5_ASAP7_75t_L g1648 ( 
.A(n_1635),
.B(n_1607),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1634),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1637),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1645),
.B(n_1607),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1632),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1628),
.A2(n_1568),
.B1(n_1577),
.B2(n_1592),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1646),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1631),
.B(n_1606),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1633),
.B(n_1608),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1638),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1630),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1652),
.B(n_1608),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1658),
.A2(n_1636),
.B(n_1639),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1658),
.A2(n_1568),
.B1(n_1592),
.B2(n_1577),
.Y(n_1661)
);

OAI21xp33_ASAP7_75t_L g1662 ( 
.A1(n_1650),
.A2(n_1612),
.B(n_1609),
.Y(n_1662)
);

O2A1O1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1648),
.A2(n_1638),
.B(n_1642),
.C(n_1640),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1652),
.Y(n_1664)
);

NAND2x1_ASAP7_75t_L g1665 ( 
.A(n_1651),
.B(n_1610),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1653),
.B(n_1641),
.C(n_1644),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_SL g1667 ( 
.A1(n_1648),
.A2(n_1625),
.B(n_1610),
.Y(n_1667)
);

AOI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1660),
.A2(n_1657),
.B1(n_1648),
.B2(n_1650),
.C(n_1656),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1659),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1664),
.B(n_1651),
.Y(n_1670)
);

AOI21xp33_ASAP7_75t_L g1671 ( 
.A1(n_1663),
.A2(n_1649),
.B(n_1654),
.Y(n_1671)
);

CKINVDCx11_ASAP7_75t_R g1672 ( 
.A(n_1665),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1670),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1669),
.Y(n_1674)
);

AOI221xp5_ASAP7_75t_L g1675 ( 
.A1(n_1668),
.A2(n_1666),
.B1(n_1661),
.B2(n_1662),
.C(n_1667),
.Y(n_1675)
);

NOR2x1_ASAP7_75t_L g1676 ( 
.A(n_1672),
.B(n_1647),
.Y(n_1676)
);

INVxp67_ASAP7_75t_SL g1677 ( 
.A(n_1671),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1670),
.Y(n_1678)
);

NAND4xp25_ASAP7_75t_L g1679 ( 
.A(n_1675),
.B(n_1676),
.C(n_1673),
.D(n_1678),
.Y(n_1679)
);

OAI211xp5_ASAP7_75t_L g1680 ( 
.A1(n_1677),
.A2(n_1655),
.B(n_1622),
.C(n_1625),
.Y(n_1680)
);

AOI22x1_ASAP7_75t_L g1681 ( 
.A1(n_1674),
.A2(n_1655),
.B1(n_1622),
.B2(n_1559),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1676),
.A2(n_1643),
.B(n_1579),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_R g1683 ( 
.A(n_1673),
.B(n_1618),
.Y(n_1683)
);

NAND5xp2_ASAP7_75t_L g1684 ( 
.A(n_1680),
.B(n_1553),
.C(n_1555),
.D(n_1561),
.E(n_1348),
.Y(n_1684)
);

NOR2xp67_ASAP7_75t_SL g1685 ( 
.A(n_1679),
.B(n_1574),
.Y(n_1685)
);

BUFx12f_ASAP7_75t_L g1686 ( 
.A(n_1683),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1686),
.B(n_1682),
.Y(n_1687)
);

NOR3xp33_ASAP7_75t_L g1688 ( 
.A(n_1687),
.B(n_1684),
.C(n_1686),
.Y(n_1688)
);

XNOR2xp5_ASAP7_75t_L g1689 ( 
.A(n_1688),
.B(n_1681),
.Y(n_1689)
);

XNOR2x1_ASAP7_75t_L g1690 ( 
.A(n_1689),
.B(n_1685),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1690),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1691),
.A2(n_1643),
.B1(n_1566),
.B2(n_1583),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1691),
.Y(n_1693)
);

OAI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1693),
.A2(n_1595),
.B1(n_1567),
.B2(n_1549),
.C(n_1560),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1692),
.B(n_1552),
.Y(n_1695)
);

AOI222xp33_ASAP7_75t_L g1696 ( 
.A1(n_1695),
.A2(n_1555),
.B1(n_1561),
.B2(n_1560),
.C1(n_1558),
.C2(n_1556),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1694),
.A2(n_1567),
.B1(n_1558),
.B2(n_1556),
.Y(n_1697)
);

AOI322xp5_ASAP7_75t_L g1698 ( 
.A1(n_1697),
.A2(n_1534),
.A3(n_1554),
.B1(n_1552),
.B2(n_1505),
.C1(n_1514),
.C2(n_1502),
.Y(n_1698)
);

NOR2x1p5_ASAP7_75t_L g1699 ( 
.A(n_1696),
.B(n_1554),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1699),
.A2(n_1698),
.B1(n_1439),
.B2(n_1545),
.Y(n_1700)
);

AOI211xp5_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_1499),
.B(n_1453),
.C(n_1456),
.Y(n_1701)
);


endmodule