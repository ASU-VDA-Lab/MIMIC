module real_jpeg_5727_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_1),
.Y(n_119)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_1),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_2),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_2),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_2),
.B(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_3),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_4),
.B(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_5),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_5),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_5),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_5),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_5),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_5),
.B(n_245),
.Y(n_244)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_7),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_7),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g245 ( 
.A(n_7),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_8),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_8),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_8),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_8),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_8),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_9),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_9),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_9),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_9),
.B(n_69),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_10),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_10),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_10),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_10),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_10),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_11),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_11),
.B(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_12),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_12),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_13),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_13),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_13),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_13),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_13),
.B(n_48),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_13),
.B(n_225),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_13),
.B(n_156),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_13),
.B(n_273),
.Y(n_272)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_15),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_15),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_15),
.B(n_82),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_15),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_15),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_15),
.B(n_249),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_15),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_16),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_16),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_16),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_16),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_16),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_16),
.B(n_54),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_16),
.B(n_276),
.Y(n_275)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_17),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_17),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g265 ( 
.A(n_17),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_196),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_195),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_166),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_22),
.B(n_166),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_99),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_65),
.C(n_76),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_24),
.B(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_42),
.C(n_51),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_25),
.A2(n_26),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_27),
.B(n_33),
.C(n_41),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_28),
.B(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_31),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_38),
.B2(n_41),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_37),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_37),
.Y(n_243)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_43),
.B(n_52),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_44),
.B(n_47),
.Y(n_292)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_50),
.Y(n_179)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_50),
.Y(n_217)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_57),
.C(n_61),
.Y(n_52)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_53),
.B(n_57),
.CI(n_61),
.CON(n_289),
.SN(n_289)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_59),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_59),
.Y(n_273)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_65),
.B(n_76),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_71),
.C(n_73),
.Y(n_113)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_69),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_86),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_78),
.B(n_81),
.C(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_86),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.C(n_95),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_87),
.B(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_91),
.A2(n_95),
.B1(n_96),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_91),
.Y(n_191)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_93),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_129),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_111),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_125),
.B1(n_126),
.B2(n_128),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_121),
.Y(n_128)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_124),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_150),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_142),
.C(n_149),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_131),
.A2(n_132),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_137),
.C(n_163),
.Y(n_162)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_142),
.A2(n_143),
.B(n_146),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_149),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_153),
.B1(n_164),
.B2(n_165),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_162),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

INVx4_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_161),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.C(n_192),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_168),
.B(n_312),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_170),
.B(n_192),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_187),
.C(n_188),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_171),
.B(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_180),
.C(n_182),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_172),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_173),
.A2(n_174),
.B1(n_177),
.B2(n_178),
.Y(n_266)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_181),
.B(n_183),
.Y(n_286)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_187),
.Y(n_306)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_193),
.Y(n_194)
);

AOI21x1_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_310),
.B(n_314),
.Y(n_196)
);

OAI21x1_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_297),
.B(n_309),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_282),
.B(n_296),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_256),
.B(n_281),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_238),
.B(n_255),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_219),
.B(n_237),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_213),
.B(n_218),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_209),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_208),
.Y(n_220)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_221),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_229),
.B2(n_230),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_232),
.C(n_234),
.Y(n_254)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_227),
.Y(n_246)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_254),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_254),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_247),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_246),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_246),
.C(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_244),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_269),
.C(n_270),
.Y(n_268)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_259),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_268),
.C(n_271),
.Y(n_295)
);

XOR2x2_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_263),
.C(n_266),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.Y(n_262)
);

INVx4_ASAP7_75t_SL g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_277),
.C(n_279),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_274)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_275),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_277),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_295),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_295),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_288),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_287),
.C(n_308),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_288),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_292),
.C(n_293),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g315 ( 
.A(n_289),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_307),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_307),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_304),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_301),
.C(n_304),
.Y(n_313)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_313),
.Y(n_314)
);


endmodule