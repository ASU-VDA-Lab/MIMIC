module fake_jpeg_11846_n_54 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_54);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_54;

wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_18),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_8),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_17),
.B1(n_16),
.B2(n_14),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_20),
.B(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_24),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_23),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_24),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_20),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_30),
.B1(n_23),
.B2(n_26),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_40),
.B1(n_41),
.B2(n_4),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_0),
.C(n_1),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_2),
.C(n_3),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_40)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_47),
.B(n_48),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_42),
.B1(n_39),
.B2(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_44),
.B(n_50),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_46),
.C(n_5),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_52),
.A2(n_4),
.B(n_6),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_7),
.C(n_8),
.Y(n_54)
);


endmodule