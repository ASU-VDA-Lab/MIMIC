module fake_netlist_6_4358_n_3243 (n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_853, n_440, n_587, n_695, n_507, n_909, n_580, n_762, n_881, n_875, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_828, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_933, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_820, n_783, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_805, n_396, n_495, n_815, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_840, n_442, n_480, n_142, n_874, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_883, n_557, n_823, n_349, n_643, n_233, n_617, n_698, n_898, n_845, n_255, n_807, n_739, n_284, n_400, n_140, n_337, n_865, n_893, n_214, n_925, n_485, n_67, n_15, n_443, n_246, n_892, n_768, n_38, n_471, n_289, n_935, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_727, n_894, n_369, n_597, n_685, n_280, n_287, n_832, n_353, n_610, n_555, n_389, n_814, n_415, n_830, n_65, n_230, n_605, n_461, n_873, n_141, n_383, n_826, n_669, n_200, n_447, n_176, n_872, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_852, n_667, n_71, n_74, n_229, n_542, n_847, n_644, n_682, n_851, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_901, n_111, n_504, n_923, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_837, n_836, n_79, n_863, n_375, n_601, n_338, n_522, n_948, n_466, n_704, n_918, n_748, n_506, n_56, n_763, n_360, n_945, n_603, n_119, n_235, n_536, n_895, n_866, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_946, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_641, n_822, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_842, n_611, n_943, n_156, n_491, n_878, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_843, n_797, n_666, n_371, n_795, n_770, n_940, n_567, n_899, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_838, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_844, n_448, n_886, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_930, n_888, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_910, n_37, n_486, n_911, n_381, n_82, n_947, n_27, n_236, n_653, n_887, n_752, n_908, n_112, n_172, n_944, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_490, n_803, n_290, n_220, n_809, n_118, n_224, n_48, n_926, n_927, n_25, n_93, n_839, n_80, n_734, n_708, n_196, n_919, n_402, n_352, n_917, n_668, n_478, n_626, n_574, n_779, n_9, n_800, n_929, n_460, n_107, n_907, n_854, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_870, n_366, n_904, n_777, n_407, n_913, n_450, n_103, n_808, n_867, n_272, n_526, n_921, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_937, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_924, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_824, n_279, n_686, n_796, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_936, n_184, n_552, n_619, n_885, n_216, n_455, n_896, n_83, n_521, n_363, n_572, n_912, n_395, n_813, n_592, n_745, n_654, n_323, n_829, n_606, n_393, n_818, n_411, n_503, n_716, n_152, n_623, n_92, n_884, n_599, n_513, n_855, n_776, n_321, n_645, n_331, n_105, n_916, n_227, n_132, n_868, n_570, n_731, n_859, n_406, n_483, n_735, n_102, n_204, n_482, n_934, n_755, n_931, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_942, n_792, n_880, n_476, n_714, n_2, n_291, n_219, n_543, n_889, n_357, n_150, n_264, n_263, n_589, n_860, n_481, n_788, n_819, n_939, n_821, n_325, n_938, n_767, n_804, n_329, n_464, n_600, n_831, n_802, n_561, n_33, n_477, n_549, n_533, n_408, n_932, n_806, n_864, n_879, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_905, n_94, n_282, n_436, n_833, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_941, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_849, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_811, n_882, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_861, n_674, n_857, n_871, n_775, n_922, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_902, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_914, n_759, n_355, n_426, n_317, n_149, n_915, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_903, n_85, n_99, n_257, n_920, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_834, n_242, n_835, n_928, n_19, n_47, n_690, n_29, n_850, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_463, n_545, n_489, n_877, n_205, n_604, n_848, n_120, n_251, n_301, n_274, n_636, n_825, n_728, n_681, n_729, n_110, n_151, n_876, n_774, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_906, n_688, n_722, n_862, n_135, n_165, n_351, n_869, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_890, n_637, n_295, n_385, n_701, n_817, n_629, n_388, n_190, n_858, n_262, n_484, n_613, n_736, n_187, n_897, n_900, n_846, n_501, n_841, n_531, n_827, n_60, n_361, n_508, n_663, n_856, n_379, n_170, n_778, n_332, n_891, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_3243);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_853;
input n_440;
input n_587;
input n_695;
input n_507;
input n_909;
input n_580;
input n_762;
input n_881;
input n_875;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_828;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_933;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_820;
input n_783;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_805;
input n_396;
input n_495;
input n_815;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_840;
input n_442;
input n_480;
input n_142;
input n_874;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_883;
input n_557;
input n_823;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_898;
input n_845;
input n_255;
input n_807;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_865;
input n_893;
input n_214;
input n_925;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_892;
input n_768;
input n_38;
input n_471;
input n_289;
input n_935;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_727;
input n_894;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_832;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_830;
input n_65;
input n_230;
input n_605;
input n_461;
input n_873;
input n_141;
input n_383;
input n_826;
input n_669;
input n_200;
input n_447;
input n_176;
input n_872;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_852;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_847;
input n_644;
input n_682;
input n_851;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_901;
input n_111;
input n_504;
input n_923;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_837;
input n_836;
input n_79;
input n_863;
input n_375;
input n_601;
input n_338;
input n_522;
input n_948;
input n_466;
input n_704;
input n_918;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_945;
input n_603;
input n_119;
input n_235;
input n_536;
input n_895;
input n_866;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_946;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_822;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_842;
input n_611;
input n_943;
input n_156;
input n_491;
input n_878;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_843;
input n_797;
input n_666;
input n_371;
input n_795;
input n_770;
input n_940;
input n_567;
input n_899;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_838;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_844;
input n_448;
input n_886;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_930;
input n_888;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_910;
input n_37;
input n_486;
input n_911;
input n_381;
input n_82;
input n_947;
input n_27;
input n_236;
input n_653;
input n_887;
input n_752;
input n_908;
input n_112;
input n_172;
input n_944;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_118;
input n_224;
input n_48;
input n_926;
input n_927;
input n_25;
input n_93;
input n_839;
input n_80;
input n_734;
input n_708;
input n_196;
input n_919;
input n_402;
input n_352;
input n_917;
input n_668;
input n_478;
input n_626;
input n_574;
input n_779;
input n_9;
input n_800;
input n_929;
input n_460;
input n_107;
input n_907;
input n_854;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_870;
input n_366;
input n_904;
input n_777;
input n_407;
input n_913;
input n_450;
input n_103;
input n_808;
input n_867;
input n_272;
input n_526;
input n_921;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_937;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_924;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_824;
input n_279;
input n_686;
input n_796;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_936;
input n_184;
input n_552;
input n_619;
input n_885;
input n_216;
input n_455;
input n_896;
input n_83;
input n_521;
input n_363;
input n_572;
input n_912;
input n_395;
input n_813;
input n_592;
input n_745;
input n_654;
input n_323;
input n_829;
input n_606;
input n_393;
input n_818;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_884;
input n_599;
input n_513;
input n_855;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_916;
input n_227;
input n_132;
input n_868;
input n_570;
input n_731;
input n_859;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_934;
input n_755;
input n_931;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_942;
input n_792;
input n_880;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_889;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_860;
input n_481;
input n_788;
input n_819;
input n_939;
input n_821;
input n_325;
input n_938;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_831;
input n_802;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_932;
input n_806;
input n_864;
input n_879;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_905;
input n_94;
input n_282;
input n_436;
input n_833;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_941;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_849;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_882;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_861;
input n_674;
input n_857;
input n_871;
input n_775;
input n_922;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_902;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_914;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_915;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_903;
input n_85;
input n_99;
input n_257;
input n_920;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_834;
input n_242;
input n_835;
input n_928;
input n_19;
input n_47;
input n_690;
input n_29;
input n_850;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_877;
input n_205;
input n_604;
input n_848;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_825;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_876;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_906;
input n_688;
input n_722;
input n_862;
input n_135;
input n_165;
input n_351;
input n_869;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_890;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_629;
input n_388;
input n_190;
input n_858;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_897;
input n_900;
input n_846;
input n_501;
input n_841;
input n_531;
input n_827;
input n_60;
input n_361;
input n_508;
input n_663;
input n_856;
input n_379;
input n_170;
input n_778;
input n_332;
input n_891;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_3243;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1674;
wire n_1199;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_3152;
wire n_1212;
wire n_2157;
wire n_2332;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_1357;
wire n_1853;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_2299;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_1172;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_3232;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_1591;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3077;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3107;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_2843;
wire n_1467;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_2370;
wire n_2612;
wire n_1446;
wire n_2591;
wire n_1815;
wire n_2214;
wire n_1658;
wire n_2593;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_2397;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_1530;
wire n_1543;
wire n_2811;
wire n_1302;
wire n_1599;
wire n_1068;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_2831;
wire n_2998;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_966;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3055;
wire n_3092;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3069;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_1165;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_2624;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_1214;
wire n_1801;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_1157;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3153;
wire n_1188;
wire n_1752;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1624;
wire n_1124;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_2476;
wire n_1515;
wire n_961;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_2377;
wire n_2178;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_2657;
wire n_1792;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_1369;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_2078;
wire n_1634;
wire n_2932;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_3209;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_2750;
wire n_1164;
wire n_1627;
wire n_1295;
wire n_2954;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_2913;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1565;
wire n_1067;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_1952;
wire n_2573;
wire n_2646;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_963;
wire n_2767;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_2707;
wire n_3240;
wire n_1514;
wire n_1863;
wire n_3037;
wire n_1646;
wire n_1139;
wire n_1714;
wire n_3179;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_2897;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_3171;
wire n_1913;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_2517;
wire n_2713;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_1432;
wire n_2208;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_3119;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_1049;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_2610;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_2868;
wire n_1698;
wire n_2231;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_998;
wire n_3200;
wire n_1665;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_1195;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3006;
wire n_2481;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_1048;
wire n_1398;
wire n_1201;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_1021;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_3142;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_1314;
wire n_1837;
wire n_964;
wire n_2218;
wire n_2788;
wire n_3196;
wire n_2435;
wire n_954;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3211;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_2990;
wire n_1773;
wire n_1775;
wire n_1286;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_2920;
wire n_1901;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_3109;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_1077;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_2803;
wire n_2100;
wire n_2993;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_1129;
wire n_2829;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_1593;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_2420;
wire n_2984;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_1037;
wire n_1397;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_2755;
wire n_3141;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3108;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_1108;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3010;
wire n_2499;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_2486;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_1043;
wire n_3040;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_3134;
wire n_1569;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_1846;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_1548;
wire n_3044;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_1758;
wire n_3221;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1914;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_1706;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_3156;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_1045;
wire n_1794;
wire n_1650;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_3091;
wire n_2695;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_2671;
wire n_2885;
wire n_2888;
wire n_2793;
wire n_2715;
wire n_2761;
wire n_1804;
wire n_2923;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_2054;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_1154;
wire n_1600;
wire n_1113;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_1098;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_2978;
wire n_2066;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_1150;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_978;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_3027;
wire n_1554;
wire n_3231;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_1120;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_2935;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_2649;
wire n_2721;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_2437;
wire n_2743;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3035;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3204;
wire n_1104;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_2934;
wire n_1109;
wire n_2222;
wire n_1276;
wire n_3176;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_1584;
wire n_2425;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_2592;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_3123;
wire n_2600;
wire n_984;
wire n_1829;
wire n_2035;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3038;
wire n_3086;
wire n_2033;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_1133;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_2795;
wire n_2471;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_2879;
wire n_967;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_1170;
wire n_1629;
wire n_2221;
wire n_1819;
wire n_1260;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3001;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_3039;
wire n_1226;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_3070;
wire n_2223;
wire n_2091;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_1449;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g949 ( 
.A(n_775),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_838),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_618),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_863),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_1),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_356),
.Y(n_954)
);

BUFx10_ASAP7_75t_L g955 ( 
.A(n_870),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_833),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_799),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_844),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_543),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_657),
.Y(n_960)
);

CKINVDCx20_ASAP7_75t_R g961 ( 
.A(n_379),
.Y(n_961)
);

INVxp67_ASAP7_75t_L g962 ( 
.A(n_825),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_92),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_149),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_899),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_798),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_150),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_908),
.Y(n_968)
);

BUFx10_ASAP7_75t_L g969 ( 
.A(n_820),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_650),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_823),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_750),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_930),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_816),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_194),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_651),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_821),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_720),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_745),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_890),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_357),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_36),
.Y(n_982)
);

CKINVDCx16_ASAP7_75t_R g983 ( 
.A(n_190),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_738),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_848),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_132),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_893),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_850),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_875),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_463),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_649),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_694),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_873),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_628),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_603),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_336),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_941),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_897),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_562),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_306),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_906),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_834),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_867),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_887),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_668),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_491),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_381),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_662),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_202),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_354),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_794),
.Y(n_1011)
);

CKINVDCx20_ASAP7_75t_R g1012 ( 
.A(n_858),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_818),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_349),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_914),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_853),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_166),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_842),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_502),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_885),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_910),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_603),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_284),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_916),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_445),
.Y(n_1025)
);

CKINVDCx16_ASAP7_75t_R g1026 ( 
.A(n_656),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_835),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_761),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_918),
.Y(n_1029)
);

CKINVDCx16_ASAP7_75t_R g1030 ( 
.A(n_549),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_119),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_929),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_658),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_936),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_928),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_901),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_877),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_470),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_876),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_198),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_164),
.Y(n_1041)
);

BUFx10_ASAP7_75t_L g1042 ( 
.A(n_840),
.Y(n_1042)
);

INVxp33_ASAP7_75t_L g1043 ( 
.A(n_605),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_444),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_41),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_247),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_558),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_477),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_200),
.Y(n_1049)
);

BUFx5_ASAP7_75t_L g1050 ( 
.A(n_634),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_826),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_384),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_712),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_347),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_637),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_513),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_684),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_646),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_889),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_896),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_423),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_836),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_679),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_382),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_776),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_473),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_604),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_246),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_813),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_596),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_903),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_674),
.Y(n_1072)
);

BUFx2_ASAP7_75t_SL g1073 ( 
.A(n_565),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_280),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_376),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_822),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_318),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_329),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_232),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_696),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_801),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_421),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_841),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_865),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_401),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_907),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_514),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_805),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_291),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_795),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_375),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_117),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_107),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_547),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_886),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_874),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_617),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_831),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_222),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_120),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_426),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_849),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_748),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_869),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_294),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_645),
.Y(n_1106)
);

CKINVDCx20_ASAP7_75t_R g1107 ( 
.A(n_880),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_318),
.Y(n_1108)
);

BUFx10_ASAP7_75t_L g1109 ( 
.A(n_692),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_648),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_576),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_97),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_915),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_882),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_878),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_920),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_183),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_372),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_425),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_827),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_864),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_341),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_487),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_797),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_832),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_75),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_859),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_82),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_488),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_70),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_156),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_385),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_824),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_922),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_872),
.Y(n_1135)
);

INVxp67_ASAP7_75t_SL g1136 ( 
.A(n_169),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_919),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_455),
.Y(n_1138)
);

BUFx10_ASAP7_75t_L g1139 ( 
.A(n_180),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_366),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_812),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_524),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_527),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_948),
.Y(n_1144)
);

BUFx5_ASAP7_75t_L g1145 ( 
.A(n_361),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_172),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_94),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_19),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_883),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_200),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_75),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_667),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_855),
.Y(n_1153)
);

BUFx10_ASAP7_75t_L g1154 ( 
.A(n_647),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_135),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_693),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_687),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_754),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_489),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_512),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_549),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_636),
.Y(n_1162)
);

BUFx5_ASAP7_75t_L g1163 ( 
.A(n_423),
.Y(n_1163)
);

INVxp67_ASAP7_75t_L g1164 ( 
.A(n_360),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_117),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_810),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_846),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_404),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_868),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_909),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_806),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_358),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_796),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_830),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_269),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_193),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_443),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_448),
.Y(n_1178)
);

CKINVDCx20_ASAP7_75t_R g1179 ( 
.A(n_325),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_42),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_465),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_226),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_852),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_811),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_735),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_246),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_190),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_829),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_898),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_879),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_121),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_309),
.Y(n_1192)
);

BUFx5_ASAP7_75t_L g1193 ( 
.A(n_415),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_946),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_837),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_894),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_800),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_118),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_296),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_845),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_891),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_847),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_856),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_132),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_809),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_33),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_697),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_802),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_814),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_347),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_41),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_725),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_718),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_707),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_467),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_25),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_751),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_804),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_843),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_925),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_888),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_71),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_911),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_649),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_917),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_871),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_471),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_786),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_286),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_653),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_817),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_476),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_652),
.Y(n_1233)
);

CKINVDCx16_ASAP7_75t_R g1234 ( 
.A(n_451),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_211),
.Y(n_1235)
);

BUFx8_ASAP7_75t_SL g1236 ( 
.A(n_14),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_927),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_146),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_654),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_866),
.Y(n_1240)
);

CKINVDCx14_ASAP7_75t_R g1241 ( 
.A(n_257),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_426),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_325),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_857),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_187),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_456),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_860),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_862),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_389),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_904),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_431),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_905),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_884),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_416),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_881),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_188),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_565),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_501),
.Y(n_1258)
);

CKINVDCx14_ASAP7_75t_R g1259 ( 
.A(n_515),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_210),
.Y(n_1260)
);

BUFx10_ASAP7_75t_L g1261 ( 
.A(n_358),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_202),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_839),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_643),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_209),
.Y(n_1265)
);

INVxp67_ASAP7_75t_L g1266 ( 
.A(n_815),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_517),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_545),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_396),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_497),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_194),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_819),
.Y(n_1272)
);

CKINVDCx16_ASAP7_75t_R g1273 ( 
.A(n_205),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_316),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_516),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_321),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_851),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_22),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_807),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_660),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_233),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_278),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_8),
.Y(n_1283)
);

BUFx10_ASAP7_75t_L g1284 ( 
.A(n_640),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_322),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_628),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_644),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_892),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_217),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_434),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_828),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_655),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_921),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_129),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_192),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_803),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_13),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_373),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_482),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_717),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_895),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_861),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_601),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_642),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_252),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_115),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_93),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_900),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_576),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_74),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_592),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_140),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_69),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_13),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_364),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_421),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_854),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_476),
.Y(n_1318)
);

INVx2_ASAP7_75t_SL g1319 ( 
.A(n_902),
.Y(n_1319)
);

CKINVDCx16_ASAP7_75t_R g1320 ( 
.A(n_808),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_940),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_274),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_419),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1050),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1050),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1070),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1050),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1050),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_983),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1050),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1145),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1145),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1145),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1145),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1145),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1163),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_955),
.Y(n_1337)
);

CKINVDCx16_ASAP7_75t_R g1338 ( 
.A(n_1026),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1163),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1236),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_950),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_952),
.Y(n_1342)
);

INVxp67_ASAP7_75t_L g1343 ( 
.A(n_1100),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1163),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_956),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1163),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_979),
.Y(n_1347)
);

INVxp67_ASAP7_75t_SL g1348 ( 
.A(n_1212),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1163),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1193),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1193),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1117),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_1004),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1193),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1193),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_957),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_1008),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1030),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1193),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_981),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_981),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_981),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_965),
.Y(n_1363)
);

INVxp67_ASAP7_75t_L g1364 ( 
.A(n_1181),
.Y(n_1364)
);

INVxp33_ASAP7_75t_SL g1365 ( 
.A(n_1017),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1094),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1094),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_1012),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_966),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1094),
.Y(n_1370)
);

INVxp67_ASAP7_75t_SL g1371 ( 
.A(n_1308),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1187),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1187),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_973),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1187),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_974),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1282),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_977),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1282),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1282),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1303),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1234),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1303),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1303),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_978),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_1307),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_980),
.Y(n_1387)
);

INVxp67_ASAP7_75t_SL g1388 ( 
.A(n_1114),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_991),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1309),
.Y(n_1390)
);

INVxp33_ASAP7_75t_L g1391 ( 
.A(n_1043),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1309),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1309),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1380),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1362),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1391),
.B(n_1241),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1367),
.Y(n_1397)
);

OA21x2_ASAP7_75t_L g1398 ( 
.A1(n_1324),
.A2(n_962),
.B(n_958),
.Y(n_1398)
);

INVx5_ASAP7_75t_L g1399 ( 
.A(n_1380),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1337),
.B(n_1223),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1375),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1325),
.A2(n_1266),
.B(n_1248),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1379),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1341),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1392),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1360),
.Y(n_1406)
);

AND2x6_ASAP7_75t_L g1407 ( 
.A(n_1389),
.B(n_1114),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1361),
.Y(n_1408)
);

AOI22x1_ASAP7_75t_SL g1409 ( 
.A1(n_1347),
.A2(n_951),
.B1(n_961),
.B2(n_960),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1366),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1348),
.B(n_1259),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1370),
.Y(n_1412)
);

INVx4_ASAP7_75t_L g1413 ( 
.A(n_1342),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1371),
.B(n_1018),
.Y(n_1414)
);

XNOR2xp5_ASAP7_75t_L g1415 ( 
.A(n_1353),
.B(n_1087),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1345),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1357),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1372),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1327),
.A2(n_971),
.B(n_949),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1373),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_SL g1421 ( 
.A(n_1389),
.B(n_1320),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1377),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1356),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1381),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1383),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1363),
.Y(n_1426)
);

INVx4_ASAP7_75t_L g1427 ( 
.A(n_1369),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1374),
.B(n_1319),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1384),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1338),
.B(n_1273),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1376),
.B(n_1314),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1390),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1328),
.A2(n_984),
.B(n_972),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1365),
.A2(n_1164),
.B1(n_970),
.B2(n_975),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1393),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1331),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1378),
.B(n_968),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1349),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1330),
.Y(n_1439)
);

INVxp67_ASAP7_75t_SL g1440 ( 
.A(n_1388),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1332),
.A2(n_1057),
.B(n_998),
.Y(n_1441)
);

BUFx8_ASAP7_75t_SL g1442 ( 
.A(n_1340),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1333),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1423),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1438),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1426),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1438),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1417),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1442),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_R g1450 ( 
.A(n_1421),
.B(n_1385),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1439),
.Y(n_1451)
);

AND3x2_ASAP7_75t_L g1452 ( 
.A(n_1396),
.B(n_1358),
.C(n_1329),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1443),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1415),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1404),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1436),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1416),
.Y(n_1457)
);

AOI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1428),
.A2(n_1335),
.B(n_1334),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1411),
.B(n_1382),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1413),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1394),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1406),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1427),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1431),
.Y(n_1464)
);

CKINVDCx20_ASAP7_75t_R g1465 ( 
.A(n_1430),
.Y(n_1465)
);

XNOR2xp5_ASAP7_75t_L g1466 ( 
.A(n_1409),
.B(n_1368),
.Y(n_1466)
);

AND3x2_ASAP7_75t_L g1467 ( 
.A(n_1400),
.B(n_1352),
.C(n_1136),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1440),
.B(n_1387),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1422),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1437),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1414),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1434),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1398),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1407),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1395),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1407),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1422),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_1424),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1424),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_R g1480 ( 
.A(n_1408),
.B(n_1015),
.Y(n_1480)
);

CKINVDCx20_ASAP7_75t_R g1481 ( 
.A(n_1402),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1410),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1425),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1420),
.Y(n_1484)
);

AO21x2_ASAP7_75t_L g1485 ( 
.A1(n_1441),
.A2(n_988),
.B(n_987),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1425),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1435),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1419),
.B(n_1336),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1435),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1412),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1433),
.Y(n_1491)
);

INVxp67_ASAP7_75t_SL g1492 ( 
.A(n_1418),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1429),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1432),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1399),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1399),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1397),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1401),
.B(n_1326),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1403),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1405),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_R g1501 ( 
.A(n_1423),
.B(n_1021),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1423),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1438),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1438),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1423),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1417),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1423),
.Y(n_1507)
);

NAND2xp33_ASAP7_75t_R g1508 ( 
.A(n_1423),
.B(n_959),
.Y(n_1508)
);

CKINVDCx20_ASAP7_75t_R g1509 ( 
.A(n_1417),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1423),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1438),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1423),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1438),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1423),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1438),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1423),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1423),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1511),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1459),
.B(n_1343),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1475),
.Y(n_1520)
);

AND2x6_ASAP7_75t_L g1521 ( 
.A(n_1498),
.B(n_1049),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1489),
.B(n_1364),
.Y(n_1522)
);

INVx4_ASAP7_75t_L g1523 ( 
.A(n_1478),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1462),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1506),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1482),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1484),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1456),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1515),
.Y(n_1529)
);

INVx4_ASAP7_75t_L g1530 ( 
.A(n_1483),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1493),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1469),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1471),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1480),
.Y(n_1534)
);

INVxp67_ASAP7_75t_SL g1535 ( 
.A(n_1515),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1499),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1500),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1451),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1470),
.B(n_1386),
.Y(n_1539)
);

OR2x6_ASAP7_75t_L g1540 ( 
.A(n_1468),
.B(n_1073),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1494),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1492),
.B(n_1039),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1515),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1486),
.B(n_1126),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1469),
.Y(n_1545)
);

INVxp33_ASAP7_75t_SL g1546 ( 
.A(n_1501),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1461),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1469),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1453),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1503),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1503),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1477),
.B(n_1256),
.Y(n_1552)
);

NAND3x1_ASAP7_75t_L g1553 ( 
.A(n_1466),
.B(n_1251),
.C(n_1242),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1487),
.Y(n_1554)
);

BUFx4f_ASAP7_75t_L g1555 ( 
.A(n_1479),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1464),
.B(n_1028),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1479),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1445),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1488),
.B(n_1104),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1491),
.B(n_1121),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1447),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_1479),
.Y(n_1562)
);

INVx4_ASAP7_75t_L g1563 ( 
.A(n_1455),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1504),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1474),
.B(n_995),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1513),
.B(n_953),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1490),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1450),
.B(n_1033),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1460),
.B(n_1107),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1497),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1458),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1457),
.B(n_1139),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1463),
.B(n_1339),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1473),
.A2(n_1069),
.B1(n_1157),
.B2(n_1065),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1476),
.B(n_1207),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_1508),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1485),
.Y(n_1577)
);

INVx4_ASAP7_75t_SL g1578 ( 
.A(n_1509),
.Y(n_1578)
);

INVxp67_ASAP7_75t_SL g1579 ( 
.A(n_1481),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1485),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1495),
.Y(n_1581)
);

INVx4_ASAP7_75t_L g1582 ( 
.A(n_1444),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1467),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_1472),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1452),
.Y(n_1585)
);

AND2x6_ASAP7_75t_L g1586 ( 
.A(n_1446),
.B(n_954),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1448),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1465),
.A2(n_1280),
.B1(n_1170),
.B2(n_992),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1496),
.B(n_963),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1502),
.B(n_1344),
.Y(n_1590)
);

INVx4_ASAP7_75t_L g1591 ( 
.A(n_1505),
.Y(n_1591)
);

INVx3_ASAP7_75t_L g1592 ( 
.A(n_1507),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1510),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1512),
.B(n_1346),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1517),
.B(n_1350),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1514),
.B(n_1516),
.Y(n_1596)
);

BUFx10_ASAP7_75t_L g1597 ( 
.A(n_1449),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1454),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1462),
.Y(n_1599)
);

INVx4_ASAP7_75t_L g1600 ( 
.A(n_1478),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1511),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1470),
.B(n_1034),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1444),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1470),
.B(n_1351),
.Y(n_1604)
);

AND2x6_ASAP7_75t_L g1605 ( 
.A(n_1459),
.B(n_1007),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1475),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1470),
.B(n_1354),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1444),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_1469),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1470),
.B(n_1355),
.Y(n_1610)
);

BUFx10_ASAP7_75t_L g1611 ( 
.A(n_1449),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1462),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1506),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1491),
.A2(n_1002),
.B1(n_1013),
.B2(n_997),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1489),
.B(n_1014),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1475),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1470),
.B(n_1359),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1470),
.B(n_1016),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1470),
.B(n_1020),
.Y(n_1619)
);

AND2x6_ASAP7_75t_L g1620 ( 
.A(n_1459),
.B(n_1025),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1506),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1470),
.B(n_1209),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1462),
.Y(n_1623)
);

NAND2xp33_ASAP7_75t_L g1624 ( 
.A(n_1470),
.B(n_985),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1475),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1470),
.B(n_1291),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1475),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1511),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1506),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1462),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1470),
.B(n_1024),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1506),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_L g1633 ( 
.A(n_1459),
.B(n_982),
.C(n_976),
.Y(n_1633)
);

INVx4_ASAP7_75t_L g1634 ( 
.A(n_1478),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1475),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1567),
.B(n_989),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1602),
.A2(n_1051),
.B1(n_1053),
.B2(n_1027),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1520),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1626),
.B(n_1062),
.Y(n_1639)
);

INVx2_ASAP7_75t_SL g1640 ( 
.A(n_1544),
.Y(n_1640)
);

A2O1A1Ixp33_ASAP7_75t_L g1641 ( 
.A1(n_1614),
.A2(n_1071),
.B(n_1086),
.C(n_1084),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1565),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1524),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1574),
.A2(n_1560),
.B1(n_1580),
.B2(n_1559),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1539),
.B(n_964),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1526),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1576),
.B(n_1052),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1606),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1577),
.A2(n_1125),
.B1(n_1144),
.B2(n_1120),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1527),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1604),
.B(n_1152),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1607),
.B(n_1156),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1531),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1525),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1519),
.B(n_1099),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1610),
.B(n_1158),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1617),
.B(n_993),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1599),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1570),
.B(n_1289),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1569),
.B(n_1055),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_SL g1661 ( 
.A(n_1596),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1584),
.B(n_1068),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1618),
.B(n_1167),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1616),
.Y(n_1664)
);

AND2x4_ASAP7_75t_SL g1665 ( 
.A(n_1523),
.B(n_955),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1625),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1556),
.B(n_1148),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1572),
.B(n_1530),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1627),
.Y(n_1669)
);

BUFx6f_ASAP7_75t_L g1670 ( 
.A(n_1529),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1619),
.B(n_1631),
.Y(n_1671)
);

AND2x6_ASAP7_75t_SL g1672 ( 
.A(n_1598),
.B(n_1310),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1612),
.A2(n_1169),
.B1(n_1174),
.B2(n_1171),
.Y(n_1673)
);

AND2x4_ASAP7_75t_SL g1674 ( 
.A(n_1600),
.B(n_969),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1623),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1573),
.B(n_1188),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1630),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1536),
.B(n_1201),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1635),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1622),
.B(n_1168),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1537),
.B(n_1208),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1590),
.B(n_1217),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1594),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_SL g1684 ( 
.A(n_1595),
.B(n_1001),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1528),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1546),
.B(n_1179),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1538),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1563),
.B(n_1003),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1549),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1542),
.B(n_1541),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1568),
.B(n_1224),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1615),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1571),
.B(n_1220),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1588),
.A2(n_1252),
.B1(n_1255),
.B2(n_1225),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1547),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1535),
.B(n_1277),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1634),
.B(n_1139),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1558),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1555),
.A2(n_1296),
.B(n_1288),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1561),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1564),
.Y(n_1701)
);

INVx8_ASAP7_75t_L g1702 ( 
.A(n_1521),
.Y(n_1702)
);

INVx4_ASAP7_75t_L g1703 ( 
.A(n_1593),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1575),
.B(n_1304),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1534),
.B(n_986),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1624),
.B(n_1301),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1566),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1592),
.B(n_1154),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1605),
.B(n_1321),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1550),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1582),
.B(n_1005),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1591),
.B(n_1011),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1551),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1545),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1579),
.A2(n_1036),
.B1(n_1037),
.B2(n_1032),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1605),
.B(n_1059),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1562),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1529),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1620),
.B(n_1060),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1554),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1620),
.B(n_1063),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1533),
.B(n_1154),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1548),
.B(n_1072),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1587),
.B(n_990),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1548),
.B(n_1076),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1543),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1518),
.B(n_1601),
.Y(n_1727)
);

NAND2x1_ASAP7_75t_L g1728 ( 
.A(n_1557),
.B(n_1029),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1543),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1613),
.B(n_967),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1557),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1628),
.B(n_1540),
.Y(n_1732)
);

CKINVDCx20_ASAP7_75t_R g1733 ( 
.A(n_1603),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1522),
.B(n_1081),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1633),
.B(n_1608),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1532),
.B(n_1083),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1521),
.B(n_1088),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1621),
.B(n_994),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1609),
.B(n_1552),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1589),
.B(n_1090),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1586),
.B(n_1095),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1581),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1585),
.A2(n_1192),
.B(n_1292),
.C(n_1160),
.Y(n_1743)
);

AOI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1586),
.A2(n_1583),
.B1(n_1098),
.B2(n_1102),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1583),
.B(n_1578),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1629),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_SL g1747 ( 
.A(n_1597),
.B(n_1611),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1632),
.B(n_1044),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1553),
.B(n_1096),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1602),
.B(n_996),
.Y(n_1750)
);

INVx5_ASAP7_75t_L g1751 ( 
.A(n_1523),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_SL g1752 ( 
.A(n_1582),
.B(n_969),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1520),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1614),
.A2(n_1035),
.B1(n_1080),
.B2(n_1029),
.Y(n_1754)
);

NOR2xp67_ASAP7_75t_L g1755 ( 
.A(n_1582),
.B(n_1103),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1602),
.B(n_1113),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1567),
.B(n_1115),
.Y(n_1757)
);

AO221x1_ASAP7_75t_L g1758 ( 
.A1(n_1576),
.A2(n_1045),
.B1(n_1085),
.B2(n_1074),
.C(n_1056),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1602),
.B(n_1116),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1614),
.A2(n_1035),
.B1(n_1080),
.B2(n_1029),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1602),
.B(n_1124),
.Y(n_1761)
);

AO22x1_ASAP7_75t_L g1762 ( 
.A1(n_1602),
.A2(n_1000),
.B1(n_1006),
.B2(n_999),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1602),
.B(n_1261),
.Y(n_1763)
);

INVxp67_ASAP7_75t_SL g1764 ( 
.A(n_1529),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1524),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1567),
.B(n_1127),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1602),
.B(n_1133),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1602),
.B(n_1009),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1602),
.B(n_1010),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1520),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1602),
.B(n_1134),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1602),
.B(n_1135),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1602),
.B(n_1137),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1520),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1602),
.B(n_1141),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1602),
.B(n_1149),
.Y(n_1776)
);

INVxp67_ASAP7_75t_SL g1777 ( 
.A(n_1529),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1524),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1567),
.B(n_1153),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1520),
.Y(n_1780)
);

INVxp67_ASAP7_75t_L g1781 ( 
.A(n_1565),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1614),
.A2(n_1080),
.B1(n_1197),
.B2(n_1035),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1524),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1602),
.B(n_1166),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1602),
.B(n_1173),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1602),
.B(n_1019),
.Y(n_1786)
);

INVx3_ASAP7_75t_L g1787 ( 
.A(n_1532),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1567),
.B(n_1183),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1567),
.B(n_1184),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1520),
.Y(n_1790)
);

AND2x4_ASAP7_75t_SL g1791 ( 
.A(n_1523),
.B(n_1042),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1559),
.A2(n_1197),
.B(n_1189),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1567),
.B(n_1185),
.Y(n_1793)
);

AOI22x1_ASAP7_75t_L g1794 ( 
.A1(n_1580),
.A2(n_1194),
.B1(n_1195),
.B2(n_1190),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1520),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1602),
.B(n_1196),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1602),
.B(n_1200),
.Y(n_1797)
);

AOI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1671),
.A2(n_1690),
.B(n_1644),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1683),
.B(n_1202),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1748),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1693),
.A2(n_1197),
.B(n_1203),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1689),
.Y(n_1802)
);

INVx2_ASAP7_75t_SL g1803 ( 
.A(n_1640),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1727),
.A2(n_1302),
.B(n_1300),
.Y(n_1804)
);

AOI21x1_ASAP7_75t_L g1805 ( 
.A1(n_1706),
.A2(n_1093),
.B(n_1092),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1696),
.A2(n_1317),
.B(n_1213),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1750),
.B(n_1205),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1768),
.B(n_1214),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1756),
.A2(n_1219),
.B(n_1218),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1638),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1759),
.A2(n_1226),
.B(n_1221),
.Y(n_1811)
);

INVx3_ASAP7_75t_L g1812 ( 
.A(n_1670),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1769),
.B(n_1786),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1648),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1643),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1639),
.B(n_1228),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1761),
.B(n_1231),
.Y(n_1817)
);

O2A1O1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1645),
.A2(n_1106),
.B(n_1108),
.C(n_1101),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1767),
.B(n_1771),
.Y(n_1819)
);

O2A1O1Ixp33_ASAP7_75t_L g1820 ( 
.A1(n_1641),
.A2(n_1123),
.B(n_1130),
.C(n_1118),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1667),
.B(n_1660),
.Y(n_1821)
);

INVx3_ASAP7_75t_L g1822 ( 
.A(n_1670),
.Y(n_1822)
);

O2A1O1Ixp33_ASAP7_75t_L g1823 ( 
.A1(n_1743),
.A2(n_1155),
.B(n_1165),
.C(n_1146),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1646),
.A2(n_1240),
.B1(n_1244),
.B2(n_1237),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1650),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1772),
.B(n_1247),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1653),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1773),
.A2(n_1253),
.B(n_1250),
.Y(n_1828)
);

AOI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1775),
.A2(n_1272),
.B(n_1263),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1682),
.A2(n_1293),
.B(n_1279),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1776),
.A2(n_1177),
.B(n_1175),
.Y(n_1831)
);

INVx1_ASAP7_75t_SL g1832 ( 
.A(n_1730),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1784),
.B(n_1022),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1785),
.B(n_1023),
.Y(n_1834)
);

INVx3_ASAP7_75t_L g1835 ( 
.A(n_1703),
.Y(n_1835)
);

A2O1A1Ixp33_ASAP7_75t_L g1836 ( 
.A1(n_1691),
.A2(n_1204),
.B(n_1233),
.C(n_1198),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1658),
.A2(n_1038),
.B1(n_1040),
.B2(n_1031),
.Y(n_1837)
);

NOR2xp67_ASAP7_75t_L g1838 ( 
.A(n_1751),
.B(n_659),
.Y(n_1838)
);

O2A1O1Ixp5_ASAP7_75t_L g1839 ( 
.A1(n_1651),
.A2(n_1268),
.B(n_1269),
.C(n_1267),
.Y(n_1839)
);

BUFx4f_ASAP7_75t_L g1840 ( 
.A(n_1702),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1796),
.B(n_1041),
.Y(n_1841)
);

OAI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1652),
.A2(n_1271),
.B(n_1270),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1647),
.B(n_1704),
.Y(n_1843)
);

AOI21x1_ASAP7_75t_L g1844 ( 
.A1(n_1792),
.A2(n_1285),
.B(n_1275),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1797),
.A2(n_1657),
.B(n_1684),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1733),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1751),
.B(n_1042),
.Y(n_1847)
);

BUFx3_ASAP7_75t_L g1848 ( 
.A(n_1654),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1656),
.B(n_1046),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1675),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1680),
.A2(n_1109),
.B1(n_1089),
.B2(n_1075),
.Y(n_1851)
);

BUFx4f_ASAP7_75t_L g1852 ( 
.A(n_1702),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1677),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1664),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1763),
.B(n_1047),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1765),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1642),
.B(n_1048),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1781),
.B(n_1054),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1676),
.A2(n_1313),
.B(n_1297),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1778),
.B(n_1058),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1732),
.A2(n_1315),
.B(n_1128),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1666),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1669),
.A2(n_1140),
.B(n_1119),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1662),
.B(n_1686),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1783),
.B(n_1061),
.Y(n_1865)
);

BUFx6f_ASAP7_75t_L g1866 ( 
.A(n_1751),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1663),
.B(n_1064),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1720),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1655),
.B(n_1066),
.Y(n_1869)
);

BUFx12f_ASAP7_75t_L g1870 ( 
.A(n_1672),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1695),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1679),
.A2(n_1211),
.B(n_1186),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1649),
.A2(n_1681),
.B(n_1678),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1659),
.B(n_1261),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1742),
.B(n_1109),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1668),
.B(n_1067),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1685),
.B(n_1077),
.Y(n_1877)
);

AOI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1753),
.A2(n_1278),
.B(n_1276),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1770),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1746),
.B(n_1305),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1687),
.B(n_1774),
.Y(n_1881)
);

AOI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1780),
.A2(n_1316),
.B(n_663),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1790),
.B(n_1078),
.Y(n_1883)
);

NAND2x1p5_ASAP7_75t_L g1884 ( 
.A(n_1787),
.B(n_661),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1724),
.B(n_1705),
.Y(n_1885)
);

BUFx4f_ASAP7_75t_L g1886 ( 
.A(n_1726),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1735),
.B(n_1079),
.Y(n_1887)
);

NOR2x1_ASAP7_75t_L g1888 ( 
.A(n_1755),
.B(n_1284),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1795),
.A2(n_665),
.B(n_664),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1698),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1700),
.B(n_1082),
.Y(n_1891)
);

INVxp67_ASAP7_75t_L g1892 ( 
.A(n_1738),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1701),
.B(n_1091),
.Y(n_1893)
);

BUFx2_ASAP7_75t_L g1894 ( 
.A(n_1718),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1723),
.A2(n_669),
.B(n_666),
.Y(n_1895)
);

O2A1O1Ixp33_ASAP7_75t_L g1896 ( 
.A1(n_1749),
.A2(n_1673),
.B(n_1709),
.C(n_1741),
.Y(n_1896)
);

OAI21xp33_ASAP7_75t_L g1897 ( 
.A1(n_1637),
.A2(n_1105),
.B(n_1097),
.Y(n_1897)
);

O2A1O1Ixp33_ASAP7_75t_L g1898 ( 
.A1(n_1716),
.A2(n_1284),
.B(n_1111),
.C(n_1112),
.Y(n_1898)
);

BUFx6f_ASAP7_75t_L g1899 ( 
.A(n_1731),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_SL g1900 ( 
.A(n_1708),
.B(n_1110),
.Y(n_1900)
);

O2A1O1Ixp33_ASAP7_75t_L g1901 ( 
.A1(n_1719),
.A2(n_1721),
.B(n_1715),
.C(n_1737),
.Y(n_1901)
);

A2O1A1Ixp33_ASAP7_75t_L g1902 ( 
.A1(n_1754),
.A2(n_1760),
.B(n_1782),
.C(n_1710),
.Y(n_1902)
);

BUFx8_ASAP7_75t_L g1903 ( 
.A(n_1661),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1713),
.B(n_1122),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1762),
.B(n_1129),
.Y(n_1905)
);

AOI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1725),
.A2(n_1757),
.B(n_1636),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1752),
.B(n_1131),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1745),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1747),
.B(n_1132),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1714),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1766),
.A2(n_671),
.B(n_670),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1739),
.B(n_1138),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1779),
.A2(n_673),
.B(n_672),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1764),
.B(n_1777),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_SL g1915 ( 
.A(n_1722),
.B(n_1697),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1813),
.B(n_1734),
.Y(n_1916)
);

O2A1O1Ixp33_ASAP7_75t_L g1917 ( 
.A1(n_1821),
.A2(n_1885),
.B(n_1843),
.C(n_1864),
.Y(n_1917)
);

A2O1A1Ixp33_ASAP7_75t_L g1918 ( 
.A1(n_1798),
.A2(n_1699),
.B(n_1694),
.C(n_1692),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_R g1919 ( 
.A(n_1908),
.B(n_1729),
.Y(n_1919)
);

OAI21xp33_ASAP7_75t_L g1920 ( 
.A1(n_1851),
.A2(n_1674),
.B(n_1665),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1868),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1819),
.B(n_1788),
.Y(n_1922)
);

INVx1_ASAP7_75t_SL g1923 ( 
.A(n_1832),
.Y(n_1923)
);

AO32x2_ASAP7_75t_L g1924 ( 
.A1(n_1837),
.A2(n_1758),
.A3(n_1794),
.B1(n_1744),
.B2(n_1736),
.Y(n_1924)
);

AOI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1892),
.A2(n_1791),
.B1(n_1789),
.B2(n_1793),
.Y(n_1925)
);

AOI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1873),
.A2(n_1688),
.B(n_1740),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1835),
.B(n_1707),
.Y(n_1927)
);

AOI21xp5_ASAP7_75t_L g1928 ( 
.A1(n_1845),
.A2(n_1712),
.B(n_1711),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1815),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_L g1930 ( 
.A(n_1848),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1833),
.B(n_1834),
.Y(n_1931)
);

CKINVDCx14_ASAP7_75t_R g1932 ( 
.A(n_1840),
.Y(n_1932)
);

INVx1_ASAP7_75t_SL g1933 ( 
.A(n_1846),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1886),
.B(n_1717),
.Y(n_1934)
);

BUFx3_ASAP7_75t_L g1935 ( 
.A(n_1903),
.Y(n_1935)
);

BUFx6f_ASAP7_75t_L g1936 ( 
.A(n_1866),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1825),
.Y(n_1937)
);

NAND3xp33_ASAP7_75t_L g1938 ( 
.A(n_1818),
.B(n_1143),
.C(n_1142),
.Y(n_1938)
);

AO22x2_ASAP7_75t_L g1939 ( 
.A1(n_1887),
.A2(n_1728),
.B1(n_2),
.B2(n_0),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1827),
.Y(n_1940)
);

AOI21x1_ASAP7_75t_L g1941 ( 
.A1(n_1906),
.A2(n_676),
.B(n_675),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1894),
.Y(n_1942)
);

BUFx3_ASAP7_75t_L g1943 ( 
.A(n_1812),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1897),
.A2(n_1150),
.B1(n_1151),
.B2(n_1147),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1850),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1841),
.B(n_1159),
.Y(n_1946)
);

OAI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1807),
.A2(n_1162),
.B1(n_1172),
.B2(n_1161),
.Y(n_1947)
);

OAI221xp5_ASAP7_75t_L g1948 ( 
.A1(n_1855),
.A2(n_1180),
.B1(n_1182),
.B2(n_1178),
.C(n_1176),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1800),
.Y(n_1949)
);

OAI21xp33_ASAP7_75t_L g1950 ( 
.A1(n_1874),
.A2(n_1199),
.B(n_1191),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1808),
.B(n_1206),
.Y(n_1951)
);

INVx3_ASAP7_75t_L g1952 ( 
.A(n_1866),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1853),
.Y(n_1953)
);

AO21x1_ASAP7_75t_L g1954 ( 
.A1(n_1896),
.A2(n_2),
.B(n_1),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1856),
.A2(n_1215),
.B1(n_1216),
.B2(n_1210),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1802),
.Y(n_1956)
);

INVx4_ASAP7_75t_L g1957 ( 
.A(n_1866),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1822),
.B(n_677),
.Y(n_1958)
);

A2O1A1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1901),
.A2(n_1227),
.B(n_1229),
.C(n_1222),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1817),
.A2(n_680),
.B(n_678),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1871),
.Y(n_1961)
);

AOI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1826),
.A2(n_682),
.B(n_681),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_R g1963 ( 
.A(n_1852),
.B(n_683),
.Y(n_1963)
);

INVx2_ASAP7_75t_SL g1964 ( 
.A(n_1803),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1890),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1849),
.B(n_1230),
.Y(n_1966)
);

AOI21xp5_ASAP7_75t_L g1967 ( 
.A1(n_1816),
.A2(n_686),
.B(n_685),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_SL g1968 ( 
.A1(n_1870),
.A2(n_1235),
.B1(n_1238),
.B2(n_1232),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1867),
.B(n_1239),
.Y(n_1969)
);

INVx5_ASAP7_75t_L g1970 ( 
.A(n_1899),
.Y(n_1970)
);

BUFx12f_ASAP7_75t_L g1971 ( 
.A(n_1880),
.Y(n_1971)
);

BUFx3_ASAP7_75t_L g1972 ( 
.A(n_1899),
.Y(n_1972)
);

OAI21x1_ASAP7_75t_L g1973 ( 
.A1(n_1844),
.A2(n_689),
.B(n_688),
.Y(n_1973)
);

A2O1A1Ixp33_ASAP7_75t_L g1974 ( 
.A1(n_1842),
.A2(n_1245),
.B(n_1246),
.C(n_1243),
.Y(n_1974)
);

OAI21x1_ASAP7_75t_L g1975 ( 
.A1(n_1889),
.A2(n_691),
.B(n_690),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1799),
.B(n_1249),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_SL g1977 ( 
.A(n_1838),
.B(n_1298),
.Y(n_1977)
);

AOI21xp5_ASAP7_75t_L g1978 ( 
.A1(n_1902),
.A2(n_698),
.B(n_695),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1810),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1914),
.A2(n_1257),
.B1(n_1258),
.B2(n_1254),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1814),
.Y(n_1981)
);

OAI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1801),
.A2(n_1262),
.B(n_1260),
.Y(n_1982)
);

BUFx6f_ASAP7_75t_L g1983 ( 
.A(n_1899),
.Y(n_1983)
);

AOI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1882),
.A2(n_700),
.B(n_699),
.Y(n_1984)
);

AOI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1915),
.A2(n_1900),
.B1(n_1876),
.B2(n_1858),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1881),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1869),
.B(n_1264),
.Y(n_1987)
);

HB1xp67_ASAP7_75t_L g1988 ( 
.A(n_1910),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1860),
.B(n_1265),
.Y(n_1989)
);

INVx3_ASAP7_75t_L g1990 ( 
.A(n_1854),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1857),
.B(n_1274),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1865),
.B(n_1281),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1909),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1862),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1912),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_L g1996 ( 
.A(n_1905),
.B(n_1283),
.Y(n_1996)
);

BUFx6f_ASAP7_75t_L g1997 ( 
.A(n_1884),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1879),
.B(n_701),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1883),
.Y(n_1999)
);

BUFx2_ASAP7_75t_L g2000 ( 
.A(n_1904),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1877),
.B(n_1286),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1805),
.Y(n_2002)
);

AOI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1830),
.A2(n_1290),
.B1(n_1294),
.B2(n_1287),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1911),
.A2(n_703),
.B(n_702),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1891),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1875),
.B(n_1295),
.Y(n_2006)
);

OAI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1893),
.A2(n_1306),
.B1(n_1311),
.B2(n_1299),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1831),
.B(n_1312),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1888),
.B(n_704),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1839),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1847),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1824),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_L g2013 ( 
.A(n_1907),
.B(n_1318),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_L g2014 ( 
.A(n_1836),
.B(n_1322),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1863),
.Y(n_2015)
);

A2O1A1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1898),
.A2(n_1323),
.B(n_4),
.C(n_0),
.Y(n_2016)
);

BUFx3_ASAP7_75t_L g2017 ( 
.A(n_1861),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1872),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1820),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1878),
.Y(n_2020)
);

INVx1_ASAP7_75t_SL g2021 ( 
.A(n_1859),
.Y(n_2021)
);

O2A1O1Ixp33_ASAP7_75t_L g2022 ( 
.A1(n_1823),
.A2(n_1809),
.B(n_1828),
.C(n_1811),
.Y(n_2022)
);

CKINVDCx20_ASAP7_75t_R g2023 ( 
.A(n_1913),
.Y(n_2023)
);

BUFx3_ASAP7_75t_L g2024 ( 
.A(n_1895),
.Y(n_2024)
);

AOI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1829),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_2025)
);

NOR2xp33_ASAP7_75t_L g2026 ( 
.A(n_1804),
.B(n_3),
.Y(n_2026)
);

A2O1A1Ixp33_ASAP7_75t_L g2027 ( 
.A1(n_1806),
.A2(n_7),
.B(n_5),
.C(n_6),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1815),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1813),
.B(n_6),
.Y(n_2029)
);

INVx3_ASAP7_75t_SL g2030 ( 
.A(n_1908),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1813),
.B(n_7),
.Y(n_2031)
);

NAND3xp33_ASAP7_75t_L g2032 ( 
.A(n_1813),
.B(n_8),
.C(n_9),
.Y(n_2032)
);

A2O1A1Ixp33_ASAP7_75t_L g2033 ( 
.A1(n_1813),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_2033)
);

OAI21x1_ASAP7_75t_L g2034 ( 
.A1(n_1798),
.A2(n_706),
.B(n_705),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1813),
.B(n_10),
.Y(n_2035)
);

BUFx6f_ASAP7_75t_L g2036 ( 
.A(n_1848),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1813),
.B(n_11),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1813),
.B(n_12),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_L g2039 ( 
.A(n_1813),
.B(n_12),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1815),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_SL g2041 ( 
.A(n_1885),
.B(n_708),
.Y(n_2041)
);

O2A1O1Ixp33_ASAP7_75t_L g2042 ( 
.A1(n_1813),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_2042)
);

AOI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_1813),
.A2(n_710),
.B(n_709),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1874),
.B(n_15),
.Y(n_2044)
);

AOI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_2029),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_2045)
);

BUFx2_ASAP7_75t_R g2046 ( 
.A(n_1935),
.Y(n_2046)
);

BUFx2_ASAP7_75t_L g2047 ( 
.A(n_1923),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1929),
.Y(n_2048)
);

AOI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_1926),
.A2(n_943),
.B(n_942),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_1917),
.B(n_17),
.Y(n_2050)
);

AOI21x1_ASAP7_75t_L g2051 ( 
.A1(n_1928),
.A2(n_713),
.B(n_711),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1940),
.Y(n_2052)
);

AOI21xp5_ASAP7_75t_SL g2053 ( 
.A1(n_1918),
.A2(n_715),
.B(n_714),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1953),
.Y(n_2054)
);

OR2x6_ASAP7_75t_L g2055 ( 
.A(n_1930),
.B(n_716),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_L g2056 ( 
.A(n_1916),
.B(n_719),
.Y(n_2056)
);

NAND3xp33_ASAP7_75t_L g2057 ( 
.A(n_2037),
.B(n_18),
.C(n_19),
.Y(n_2057)
);

OAI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_2039),
.A2(n_20),
.B(n_21),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_2000),
.B(n_20),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1931),
.B(n_21),
.Y(n_2060)
);

NAND3xp33_ASAP7_75t_L g2061 ( 
.A(n_2014),
.B(n_22),
.C(n_23),
.Y(n_2061)
);

OAI21xp5_ASAP7_75t_L g2062 ( 
.A1(n_1959),
.A2(n_23),
.B(n_24),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_1933),
.B(n_24),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_2022),
.A2(n_939),
.B(n_938),
.Y(n_2064)
);

INVxp67_ASAP7_75t_L g2065 ( 
.A(n_1949),
.Y(n_2065)
);

OAI21x1_ASAP7_75t_L g2066 ( 
.A1(n_2034),
.A2(n_722),
.B(n_721),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1987),
.B(n_25),
.Y(n_2067)
);

AOI221x1_ASAP7_75t_L g2068 ( 
.A1(n_1939),
.A2(n_2016),
.B1(n_2033),
.B2(n_2032),
.C(n_2027),
.Y(n_2068)
);

OAI21x1_ASAP7_75t_L g2069 ( 
.A1(n_1941),
.A2(n_724),
.B(n_723),
.Y(n_2069)
);

OAI21x1_ASAP7_75t_L g2070 ( 
.A1(n_1973),
.A2(n_727),
.B(n_726),
.Y(n_2070)
);

AOI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_1922),
.A2(n_931),
.B(n_926),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2044),
.B(n_26),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1919),
.Y(n_2073)
);

OAI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_1996),
.A2(n_26),
.B(n_27),
.Y(n_2074)
);

BUFx6f_ASAP7_75t_L g2075 ( 
.A(n_1930),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2040),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1999),
.B(n_27),
.Y(n_2077)
);

OAI21x1_ASAP7_75t_L g2078 ( 
.A1(n_1975),
.A2(n_729),
.B(n_728),
.Y(n_2078)
);

AOI21x1_ASAP7_75t_L g2079 ( 
.A1(n_1978),
.A2(n_731),
.B(n_730),
.Y(n_2079)
);

AO31x2_ASAP7_75t_L g2080 ( 
.A1(n_1954),
.A2(n_733),
.A3(n_734),
.B(n_732),
.Y(n_2080)
);

AOI21xp5_ASAP7_75t_L g2081 ( 
.A1(n_2024),
.A2(n_947),
.B(n_945),
.Y(n_2081)
);

AOI31xp67_ASAP7_75t_L g2082 ( 
.A1(n_2002),
.A2(n_737),
.A3(n_739),
.B(n_736),
.Y(n_2082)
);

INVx1_ASAP7_75t_SL g2083 ( 
.A(n_1942),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1961),
.Y(n_2084)
);

INVx2_ASAP7_75t_SL g2085 ( 
.A(n_2036),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_SL g2086 ( 
.A(n_1985),
.B(n_28),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1956),
.Y(n_2087)
);

AO31x2_ASAP7_75t_L g2088 ( 
.A1(n_2010),
.A2(n_741),
.A3(n_742),
.B(n_740),
.Y(n_2088)
);

AOI21xp5_ASAP7_75t_L g2089 ( 
.A1(n_2041),
.A2(n_932),
.B(n_924),
.Y(n_2089)
);

OAI21x1_ASAP7_75t_SL g2090 ( 
.A1(n_2042),
.A2(n_28),
.B(n_29),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_2036),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1986),
.B(n_29),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2005),
.B(n_30),
.Y(n_2093)
);

NOR2xp67_ASAP7_75t_L g2094 ( 
.A(n_1964),
.B(n_1925),
.Y(n_2094)
);

INVx3_ASAP7_75t_L g2095 ( 
.A(n_1943),
.Y(n_2095)
);

AO21x1_ASAP7_75t_L g2096 ( 
.A1(n_2026),
.A2(n_30),
.B(n_31),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_1988),
.B(n_31),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_SL g2098 ( 
.A(n_2030),
.B(n_743),
.Y(n_2098)
);

CKINVDCx8_ASAP7_75t_R g2099 ( 
.A(n_1970),
.Y(n_2099)
);

OR2x2_ASAP7_75t_L g2100 ( 
.A(n_2031),
.B(n_2035),
.Y(n_2100)
);

OAI21x1_ASAP7_75t_L g2101 ( 
.A1(n_2015),
.A2(n_746),
.B(n_744),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1937),
.Y(n_2102)
);

INVx2_ASAP7_75t_SL g2103 ( 
.A(n_1936),
.Y(n_2103)
);

BUFx3_ASAP7_75t_L g2104 ( 
.A(n_1971),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1945),
.Y(n_2105)
);

OAI21x1_ASAP7_75t_L g2106 ( 
.A1(n_2018),
.A2(n_749),
.B(n_747),
.Y(n_2106)
);

AOI21x1_ASAP7_75t_L g2107 ( 
.A1(n_2019),
.A2(n_753),
.B(n_752),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1991),
.B(n_32),
.Y(n_2108)
);

CKINVDCx14_ASAP7_75t_R g2109 ( 
.A(n_1932),
.Y(n_2109)
);

OA21x2_ASAP7_75t_L g2110 ( 
.A1(n_2020),
.A2(n_756),
.B(n_755),
.Y(n_2110)
);

O2A1O1Ixp5_ASAP7_75t_SL g2111 ( 
.A1(n_2038),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_2111)
);

AOI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_1984),
.A2(n_933),
.B(n_923),
.Y(n_2112)
);

AOI21xp5_ASAP7_75t_L g2113 ( 
.A1(n_2021),
.A2(n_935),
.B(n_934),
.Y(n_2113)
);

NAND3xp33_ASAP7_75t_L g2114 ( 
.A(n_2003),
.B(n_2025),
.C(n_2013),
.Y(n_2114)
);

AOI21xp5_ASAP7_75t_SL g2115 ( 
.A1(n_1920),
.A2(n_758),
.B(n_757),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1951),
.B(n_1921),
.Y(n_2116)
);

AOI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_2023),
.A2(n_944),
.B(n_937),
.Y(n_2117)
);

A2O1A1Ixp33_ASAP7_75t_L g2118 ( 
.A1(n_1948),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_2118)
);

AOI21xp5_ASAP7_75t_L g2119 ( 
.A1(n_2004),
.A2(n_913),
.B(n_912),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_1972),
.B(n_759),
.Y(n_2120)
);

OAI21x1_ASAP7_75t_L g2121 ( 
.A1(n_1960),
.A2(n_762),
.B(n_760),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1946),
.B(n_35),
.Y(n_2122)
);

OAI22xp5_ASAP7_75t_L g2123 ( 
.A1(n_1995),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_2123)
);

OAI21x1_ASAP7_75t_L g2124 ( 
.A1(n_1962),
.A2(n_764),
.B(n_763),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1966),
.B(n_37),
.Y(n_2125)
);

BUFx3_ASAP7_75t_L g2126 ( 
.A(n_1936),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2102),
.Y(n_2127)
);

OAI21x1_ASAP7_75t_L g2128 ( 
.A1(n_2051),
.A2(n_2043),
.B(n_1967),
.Y(n_2128)
);

AOI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_2114),
.A2(n_1993),
.B1(n_2006),
.B2(n_2009),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2105),
.Y(n_2130)
);

AO21x2_ASAP7_75t_L g2131 ( 
.A1(n_2064),
.A2(n_1982),
.B(n_2008),
.Y(n_2131)
);

OAI21x1_ASAP7_75t_L g2132 ( 
.A1(n_2069),
.A2(n_2028),
.B(n_2012),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2048),
.Y(n_2133)
);

HB1xp67_ASAP7_75t_L g2134 ( 
.A(n_2065),
.Y(n_2134)
);

OAI21x1_ASAP7_75t_L g2135 ( 
.A1(n_2066),
.A2(n_1979),
.B(n_1965),
.Y(n_2135)
);

INVx1_ASAP7_75t_SL g2136 ( 
.A(n_2047),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2052),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2054),
.Y(n_2138)
);

CKINVDCx11_ASAP7_75t_R g2139 ( 
.A(n_2099),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2076),
.Y(n_2140)
);

AO32x2_ASAP7_75t_L g2141 ( 
.A1(n_2123),
.A2(n_1980),
.A3(n_1947),
.B1(n_2007),
.B2(n_2096),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2084),
.Y(n_2142)
);

AOI21xp33_ASAP7_75t_L g2143 ( 
.A1(n_2100),
.A2(n_2017),
.B(n_1938),
.Y(n_2143)
);

AND2x4_ASAP7_75t_L g2144 ( 
.A(n_2083),
.B(n_1970),
.Y(n_2144)
);

CKINVDCx5p33_ASAP7_75t_R g2145 ( 
.A(n_2073),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2087),
.Y(n_2146)
);

INVx2_ASAP7_75t_SL g2147 ( 
.A(n_2075),
.Y(n_2147)
);

BUFx3_ASAP7_75t_L g2148 ( 
.A(n_2075),
.Y(n_2148)
);

INVx3_ASAP7_75t_L g2149 ( 
.A(n_2095),
.Y(n_2149)
);

BUFx2_ASAP7_75t_L g2150 ( 
.A(n_2088),
.Y(n_2150)
);

OAI21x1_ASAP7_75t_L g2151 ( 
.A1(n_2070),
.A2(n_1994),
.B(n_1981),
.Y(n_2151)
);

AO21x1_ASAP7_75t_L g2152 ( 
.A1(n_2050),
.A2(n_1977),
.B(n_1976),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2092),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2116),
.B(n_2060),
.Y(n_2154)
);

OAI22xp5_ASAP7_75t_L g2155 ( 
.A1(n_2094),
.A2(n_2011),
.B1(n_1974),
.B2(n_1944),
.Y(n_2155)
);

OAI22xp5_ASAP7_75t_L g2156 ( 
.A1(n_2108),
.A2(n_1989),
.B1(n_1992),
.B2(n_1934),
.Y(n_2156)
);

OAI21x1_ASAP7_75t_L g2157 ( 
.A1(n_2078),
.A2(n_1990),
.B(n_1927),
.Y(n_2157)
);

AOI22xp33_ASAP7_75t_L g2158 ( 
.A1(n_2074),
.A2(n_1939),
.B1(n_1950),
.B2(n_1969),
.Y(n_2158)
);

AOI22xp33_ASAP7_75t_SL g2159 ( 
.A1(n_2058),
.A2(n_2062),
.B1(n_2061),
.B2(n_2057),
.Y(n_2159)
);

CKINVDCx5p33_ASAP7_75t_R g2160 ( 
.A(n_2109),
.Y(n_2160)
);

OAI22xp33_ASAP7_75t_L g2161 ( 
.A1(n_2045),
.A2(n_1997),
.B1(n_2001),
.B2(n_1957),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_2077),
.Y(n_2162)
);

AO21x2_ASAP7_75t_L g2163 ( 
.A1(n_2053),
.A2(n_1963),
.B(n_1955),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2120),
.Y(n_2164)
);

AO21x2_ASAP7_75t_L g2165 ( 
.A1(n_2079),
.A2(n_1998),
.B(n_1924),
.Y(n_2165)
);

O2A1O1Ixp33_ASAP7_75t_SL g2166 ( 
.A1(n_2118),
.A2(n_1952),
.B(n_1924),
.C(n_1997),
.Y(n_2166)
);

BUFx12f_ASAP7_75t_L g2167 ( 
.A(n_2085),
.Y(n_2167)
);

CKINVDCx20_ASAP7_75t_R g2168 ( 
.A(n_2104),
.Y(n_2168)
);

O2A1O1Ixp33_ASAP7_75t_SL g2169 ( 
.A1(n_2086),
.A2(n_40),
.B(n_42),
.C(n_39),
.Y(n_2169)
);

HB1xp67_ASAP7_75t_L g2170 ( 
.A(n_2097),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2088),
.Y(n_2171)
);

OAI22xp5_ASAP7_75t_L g2172 ( 
.A1(n_2056),
.A2(n_1958),
.B1(n_1983),
.B2(n_1968),
.Y(n_2172)
);

OAI21x1_ASAP7_75t_L g2173 ( 
.A1(n_2101),
.A2(n_1983),
.B(n_766),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2154),
.B(n_2093),
.Y(n_2174)
);

AO21x2_ASAP7_75t_L g2175 ( 
.A1(n_2171),
.A2(n_2128),
.B(n_2152),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2127),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2153),
.B(n_2122),
.Y(n_2177)
);

INVxp67_ASAP7_75t_SL g2178 ( 
.A(n_2132),
.Y(n_2178)
);

OAI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_2159),
.A2(n_2068),
.B(n_2117),
.Y(n_2179)
);

AOI21xp5_ASAP7_75t_L g2180 ( 
.A1(n_2131),
.A2(n_2115),
.B(n_2049),
.Y(n_2180)
);

AND2x4_ASAP7_75t_L g2181 ( 
.A(n_2136),
.B(n_2091),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2130),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2170),
.B(n_2072),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2162),
.B(n_2125),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2134),
.B(n_2067),
.Y(n_2185)
);

OAI21x1_ASAP7_75t_L g2186 ( 
.A1(n_2173),
.A2(n_2107),
.B(n_2121),
.Y(n_2186)
);

OAI21xp5_ASAP7_75t_L g2187 ( 
.A1(n_2129),
.A2(n_2071),
.B(n_2089),
.Y(n_2187)
);

OAI21x1_ASAP7_75t_L g2188 ( 
.A1(n_2157),
.A2(n_2124),
.B(n_2106),
.Y(n_2188)
);

AOI22x1_ASAP7_75t_L g2189 ( 
.A1(n_2149),
.A2(n_2090),
.B1(n_2081),
.B2(n_2113),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2133),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2137),
.B(n_2063),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2138),
.Y(n_2192)
);

BUFx8_ASAP7_75t_L g2193 ( 
.A(n_2167),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2140),
.B(n_2059),
.Y(n_2194)
);

OAI21x1_ASAP7_75t_L g2195 ( 
.A1(n_2135),
.A2(n_2112),
.B(n_2119),
.Y(n_2195)
);

OAI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_2158),
.A2(n_2055),
.B1(n_2046),
.B2(n_2103),
.Y(n_2196)
);

AOI22xp33_ASAP7_75t_L g2197 ( 
.A1(n_2143),
.A2(n_2055),
.B1(n_2098),
.B2(n_2110),
.Y(n_2197)
);

OAI21x1_ASAP7_75t_SL g2198 ( 
.A1(n_2155),
.A2(n_2111),
.B(n_2082),
.Y(n_2198)
);

AO21x2_ASAP7_75t_L g2199 ( 
.A1(n_2165),
.A2(n_2080),
.B(n_2126),
.Y(n_2199)
);

OAI21x1_ASAP7_75t_L g2200 ( 
.A1(n_2151),
.A2(n_2080),
.B(n_767),
.Y(n_2200)
);

INVx6_ASAP7_75t_L g2201 ( 
.A(n_2148),
.Y(n_2201)
);

OAI21x1_ASAP7_75t_L g2202 ( 
.A1(n_2146),
.A2(n_768),
.B(n_765),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2142),
.Y(n_2203)
);

AOI21xp5_ASAP7_75t_L g2204 ( 
.A1(n_2163),
.A2(n_770),
.B(n_769),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2156),
.B(n_38),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_2150),
.Y(n_2206)
);

AO31x2_ASAP7_75t_L g2207 ( 
.A1(n_2150),
.A2(n_44),
.A3(n_40),
.B(n_43),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2141),
.Y(n_2208)
);

AO31x2_ASAP7_75t_L g2209 ( 
.A1(n_2172),
.A2(n_45),
.A3(n_43),
.B(n_44),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2164),
.B(n_45),
.Y(n_2210)
);

BUFx6f_ASAP7_75t_L g2211 ( 
.A(n_2139),
.Y(n_2211)
);

AOI21xp5_ASAP7_75t_L g2212 ( 
.A1(n_2166),
.A2(n_772),
.B(n_771),
.Y(n_2212)
);

BUFx2_ASAP7_75t_L g2213 ( 
.A(n_2144),
.Y(n_2213)
);

OAI21xp5_ASAP7_75t_L g2214 ( 
.A1(n_2161),
.A2(n_774),
.B(n_773),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_2141),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_2147),
.B(n_777),
.Y(n_2216)
);

OAI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_2168),
.A2(n_2160),
.B1(n_2145),
.B2(n_2169),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2127),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2127),
.Y(n_2219)
);

AO31x2_ASAP7_75t_L g2220 ( 
.A1(n_2150),
.A2(n_48),
.A3(n_46),
.B(n_47),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2133),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2133),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2154),
.B(n_46),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2176),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2182),
.Y(n_2225)
);

AO21x2_ASAP7_75t_L g2226 ( 
.A1(n_2198),
.A2(n_47),
.B(n_48),
.Y(n_2226)
);

INVx3_ASAP7_75t_L g2227 ( 
.A(n_2181),
.Y(n_2227)
);

NAND2x1_ASAP7_75t_L g2228 ( 
.A(n_2206),
.B(n_49),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2221),
.Y(n_2229)
);

INVxp33_ASAP7_75t_SL g2230 ( 
.A(n_2185),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2222),
.B(n_50),
.Y(n_2231)
);

INVx3_ASAP7_75t_L g2232 ( 
.A(n_2201),
.Y(n_2232)
);

OR2x6_ASAP7_75t_L g2233 ( 
.A(n_2179),
.B(n_778),
.Y(n_2233)
);

OAI21x1_ASAP7_75t_L g2234 ( 
.A1(n_2180),
.A2(n_780),
.B(n_779),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2218),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2213),
.B(n_50),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2219),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2190),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2174),
.B(n_51),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2192),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2203),
.Y(n_2241)
);

INVx1_ASAP7_75t_SL g2242 ( 
.A(n_2183),
.Y(n_2242)
);

AND2x4_ASAP7_75t_L g2243 ( 
.A(n_2191),
.B(n_781),
.Y(n_2243)
);

OR2x2_ASAP7_75t_L g2244 ( 
.A(n_2215),
.B(n_51),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2175),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2208),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2207),
.Y(n_2247)
);

INVx2_ASAP7_75t_SL g2248 ( 
.A(n_2211),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2207),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2177),
.B(n_52),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_L g2251 ( 
.A(n_2184),
.B(n_52),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2220),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2199),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2220),
.Y(n_2254)
);

HB1xp67_ASAP7_75t_L g2255 ( 
.A(n_2194),
.Y(n_2255)
);

BUFx2_ASAP7_75t_L g2256 ( 
.A(n_2193),
.Y(n_2256)
);

BUFx3_ASAP7_75t_L g2257 ( 
.A(n_2211),
.Y(n_2257)
);

CKINVDCx8_ASAP7_75t_R g2258 ( 
.A(n_2216),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2178),
.Y(n_2259)
);

OAI21x1_ASAP7_75t_L g2260 ( 
.A1(n_2195),
.A2(n_783),
.B(n_782),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2210),
.B(n_2223),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2188),
.Y(n_2262)
);

INVx3_ASAP7_75t_L g2263 ( 
.A(n_2202),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2200),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2209),
.B(n_53),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2186),
.Y(n_2266)
);

BUFx12f_ASAP7_75t_L g2267 ( 
.A(n_2214),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2205),
.Y(n_2268)
);

HB1xp67_ASAP7_75t_L g2269 ( 
.A(n_2209),
.Y(n_2269)
);

OAI21xp5_ASAP7_75t_L g2270 ( 
.A1(n_2187),
.A2(n_53),
.B(n_54),
.Y(n_2270)
);

INVx2_ASAP7_75t_SL g2271 ( 
.A(n_2189),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2197),
.B(n_54),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2217),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2196),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2212),
.Y(n_2275)
);

HB1xp67_ASAP7_75t_L g2276 ( 
.A(n_2204),
.Y(n_2276)
);

OA21x2_ASAP7_75t_L g2277 ( 
.A1(n_2208),
.A2(n_55),
.B(n_56),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2176),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2176),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2176),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_2213),
.B(n_55),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2221),
.Y(n_2282)
);

AND2x4_ASAP7_75t_L g2283 ( 
.A(n_2213),
.B(n_784),
.Y(n_2283)
);

INVxp67_ASAP7_75t_L g2284 ( 
.A(n_2185),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2176),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2176),
.Y(n_2286)
);

BUFx2_ASAP7_75t_L g2287 ( 
.A(n_2213),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2176),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2213),
.B(n_56),
.Y(n_2289)
);

INVx3_ASAP7_75t_L g2290 ( 
.A(n_2181),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2221),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2221),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2213),
.B(n_57),
.Y(n_2293)
);

AOI22xp5_ASAP7_75t_L g2294 ( 
.A1(n_2179),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_2294)
);

OR2x2_ASAP7_75t_L g2295 ( 
.A(n_2206),
.B(n_58),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_2206),
.B(n_59),
.Y(n_2296)
);

OAI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_2233),
.A2(n_2294),
.B1(n_2267),
.B2(n_2270),
.Y(n_2297)
);

NAND3xp33_ASAP7_75t_L g2298 ( 
.A(n_2276),
.B(n_60),
.C(n_61),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2224),
.Y(n_2299)
);

AOI22xp33_ASAP7_75t_L g2300 ( 
.A1(n_2233),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_2300)
);

AOI21xp33_ASAP7_75t_SL g2301 ( 
.A1(n_2273),
.A2(n_62),
.B(n_63),
.Y(n_2301)
);

AOI21xp5_ASAP7_75t_L g2302 ( 
.A1(n_2271),
.A2(n_787),
.B(n_785),
.Y(n_2302)
);

OAI211xp5_ASAP7_75t_SL g2303 ( 
.A1(n_2268),
.A2(n_2272),
.B(n_2239),
.C(n_2284),
.Y(n_2303)
);

OR2x6_ASAP7_75t_L g2304 ( 
.A(n_2287),
.B(n_63),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2225),
.Y(n_2305)
);

AOI222xp33_ASAP7_75t_L g2306 ( 
.A1(n_2265),
.A2(n_66),
.B1(n_68),
.B2(n_64),
.C1(n_65),
.C2(n_67),
.Y(n_2306)
);

OR2x2_ASAP7_75t_L g2307 ( 
.A(n_2242),
.B(n_64),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2235),
.Y(n_2308)
);

AOI22xp33_ASAP7_75t_SL g2309 ( 
.A1(n_2275),
.A2(n_67),
.B1(n_68),
.B2(n_66),
.Y(n_2309)
);

INVx2_ASAP7_75t_SL g2310 ( 
.A(n_2257),
.Y(n_2310)
);

OAI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_2274),
.A2(n_70),
.B1(n_65),
.B2(n_69),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_2255),
.B(n_71),
.Y(n_2312)
);

OA21x2_ASAP7_75t_L g2313 ( 
.A1(n_2245),
.A2(n_72),
.B(n_73),
.Y(n_2313)
);

AOI21xp5_ASAP7_75t_L g2314 ( 
.A1(n_2234),
.A2(n_789),
.B(n_788),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_L g2315 ( 
.A(n_2230),
.B(n_72),
.Y(n_2315)
);

AOI22xp33_ASAP7_75t_SL g2316 ( 
.A1(n_2269),
.A2(n_76),
.B1(n_77),
.B2(n_74),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2237),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2238),
.Y(n_2318)
);

AOI22xp33_ASAP7_75t_L g2319 ( 
.A1(n_2226),
.A2(n_77),
.B1(n_73),
.B2(n_76),
.Y(n_2319)
);

OAI22xp33_ASAP7_75t_L g2320 ( 
.A1(n_2228),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_2320)
);

AOI21xp5_ASAP7_75t_L g2321 ( 
.A1(n_2264),
.A2(n_791),
.B(n_790),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2240),
.Y(n_2322)
);

AOI22xp33_ASAP7_75t_L g2323 ( 
.A1(n_2261),
.A2(n_2290),
.B1(n_2227),
.B2(n_2251),
.Y(n_2323)
);

AOI33xp33_ASAP7_75t_L g2324 ( 
.A1(n_2250),
.A2(n_80),
.A3(n_82),
.B1(n_78),
.B2(n_79),
.B3(n_81),
.Y(n_2324)
);

INVx3_ASAP7_75t_L g2325 ( 
.A(n_2232),
.Y(n_2325)
);

INVx1_ASAP7_75t_SL g2326 ( 
.A(n_2256),
.Y(n_2326)
);

OAI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_2258),
.A2(n_84),
.B1(n_81),
.B2(n_83),
.Y(n_2327)
);

OAI211xp5_ASAP7_75t_L g2328 ( 
.A1(n_2277),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_2328)
);

AOI22xp33_ASAP7_75t_L g2329 ( 
.A1(n_2263),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_2329)
);

AOI22xp33_ASAP7_75t_L g2330 ( 
.A1(n_2243),
.A2(n_2283),
.B1(n_2277),
.B2(n_2249),
.Y(n_2330)
);

OA21x2_ASAP7_75t_L g2331 ( 
.A1(n_2253),
.A2(n_86),
.B(n_87),
.Y(n_2331)
);

OR2x2_ASAP7_75t_L g2332 ( 
.A(n_2229),
.B(n_88),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2278),
.Y(n_2333)
);

OAI22xp33_ASAP7_75t_L g2334 ( 
.A1(n_2244),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_2334)
);

AOI22xp33_ASAP7_75t_L g2335 ( 
.A1(n_2247),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_2335)
);

OAI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_2231),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_2336)
);

AOI221xp5_ASAP7_75t_L g2337 ( 
.A1(n_2252),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.C(n_97),
.Y(n_2337)
);

AND2x4_ASAP7_75t_L g2338 ( 
.A(n_2282),
.B(n_95),
.Y(n_2338)
);

INVxp67_ASAP7_75t_L g2339 ( 
.A(n_2279),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2241),
.B(n_96),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2280),
.Y(n_2341)
);

AOI22xp33_ASAP7_75t_SL g2342 ( 
.A1(n_2254),
.A2(n_100),
.B1(n_101),
.B2(n_99),
.Y(n_2342)
);

AOI22xp33_ASAP7_75t_L g2343 ( 
.A1(n_2236),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_2343)
);

AOI22xp33_ASAP7_75t_L g2344 ( 
.A1(n_2281),
.A2(n_102),
.B1(n_98),
.B2(n_101),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2285),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2286),
.Y(n_2346)
);

AOI22xp33_ASAP7_75t_L g2347 ( 
.A1(n_2289),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2291),
.B(n_103),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2292),
.B(n_104),
.Y(n_2349)
);

CKINVDCx5p33_ASAP7_75t_R g2350 ( 
.A(n_2248),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2288),
.Y(n_2351)
);

OR2x2_ASAP7_75t_L g2352 ( 
.A(n_2259),
.B(n_105),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2295),
.B(n_105),
.Y(n_2353)
);

AOI22xp33_ASAP7_75t_L g2354 ( 
.A1(n_2293),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_2354)
);

NAND2x1_ASAP7_75t_L g2355 ( 
.A(n_2266),
.B(n_106),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2246),
.Y(n_2356)
);

BUFx6f_ASAP7_75t_L g2357 ( 
.A(n_2296),
.Y(n_2357)
);

AOI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_2260),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2262),
.B(n_109),
.Y(n_2359)
);

AOI22xp33_ASAP7_75t_L g2360 ( 
.A1(n_2267),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_2360)
);

OR2x2_ASAP7_75t_L g2361 ( 
.A(n_2242),
.B(n_113),
.Y(n_2361)
);

INVx5_ASAP7_75t_L g2362 ( 
.A(n_2233),
.Y(n_2362)
);

OR2x2_ASAP7_75t_L g2363 ( 
.A(n_2242),
.B(n_114),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2255),
.B(n_114),
.Y(n_2364)
);

AOI22xp33_ASAP7_75t_L g2365 ( 
.A1(n_2267),
.A2(n_118),
.B1(n_115),
.B2(n_116),
.Y(n_2365)
);

OAI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2270),
.A2(n_116),
.B(n_119),
.Y(n_2366)
);

OAI21x1_ASAP7_75t_L g2367 ( 
.A1(n_2245),
.A2(n_120),
.B(n_121),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2224),
.Y(n_2368)
);

OAI22xp5_ASAP7_75t_L g2369 ( 
.A1(n_2233),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_2369)
);

OAI221xp5_ASAP7_75t_L g2370 ( 
.A1(n_2270),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.C(n_128),
.Y(n_2370)
);

OAI221xp5_ASAP7_75t_L g2371 ( 
.A1(n_2270),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.C(n_128),
.Y(n_2371)
);

NAND4xp25_ASAP7_75t_L g2372 ( 
.A(n_2294),
.B(n_131),
.C(n_129),
.D(n_130),
.Y(n_2372)
);

AOI22xp5_ASAP7_75t_L g2373 ( 
.A1(n_2267),
.A2(n_133),
.B1(n_130),
.B2(n_131),
.Y(n_2373)
);

AOI21xp5_ASAP7_75t_L g2374 ( 
.A1(n_2271),
.A2(n_793),
.B(n_792),
.Y(n_2374)
);

BUFx4f_ASAP7_75t_L g2375 ( 
.A(n_2256),
.Y(n_2375)
);

OAI22xp5_ASAP7_75t_L g2376 ( 
.A1(n_2233),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_2376)
);

AOI22xp33_ASAP7_75t_L g2377 ( 
.A1(n_2267),
.A2(n_137),
.B1(n_134),
.B2(n_136),
.Y(n_2377)
);

A2O1A1Ixp33_ASAP7_75t_L g2378 ( 
.A1(n_2270),
.A2(n_138),
.B(n_139),
.C(n_137),
.Y(n_2378)
);

AOI211xp5_ASAP7_75t_L g2379 ( 
.A1(n_2270),
.A2(n_139),
.B(n_136),
.C(n_138),
.Y(n_2379)
);

OAI21x1_ASAP7_75t_L g2380 ( 
.A1(n_2245),
.A2(n_140),
.B(n_141),
.Y(n_2380)
);

OR2x2_ASAP7_75t_L g2381 ( 
.A(n_2242),
.B(n_141),
.Y(n_2381)
);

OR2x2_ASAP7_75t_L g2382 ( 
.A(n_2242),
.B(n_142),
.Y(n_2382)
);

AOI33xp33_ASAP7_75t_L g2383 ( 
.A1(n_2265),
.A2(n_145),
.A3(n_147),
.B1(n_143),
.B2(n_144),
.B3(n_146),
.Y(n_2383)
);

AND2x4_ASAP7_75t_L g2384 ( 
.A(n_2287),
.B(n_147),
.Y(n_2384)
);

OAI22xp5_ASAP7_75t_L g2385 ( 
.A1(n_2233),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_2385)
);

AOI22xp33_ASAP7_75t_L g2386 ( 
.A1(n_2267),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_2386)
);

AOI22xp33_ASAP7_75t_L g2387 ( 
.A1(n_2267),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_2387)
);

OAI22xp33_ASAP7_75t_L g2388 ( 
.A1(n_2233),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2357),
.B(n_2323),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2356),
.Y(n_2390)
);

OR2x2_ASAP7_75t_L g2391 ( 
.A(n_2339),
.B(n_157),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2308),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2299),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2318),
.Y(n_2394)
);

NOR2x1_ASAP7_75t_L g2395 ( 
.A(n_2325),
.B(n_157),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2305),
.B(n_158),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2317),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2322),
.Y(n_2398)
);

HB1xp67_ASAP7_75t_L g2399 ( 
.A(n_2346),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2333),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2341),
.Y(n_2401)
);

OR2x2_ASAP7_75t_L g2402 ( 
.A(n_2351),
.B(n_158),
.Y(n_2402)
);

BUFx2_ASAP7_75t_L g2403 ( 
.A(n_2375),
.Y(n_2403)
);

INVx3_ASAP7_75t_L g2404 ( 
.A(n_2326),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2345),
.B(n_159),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2368),
.B(n_159),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2352),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2332),
.Y(n_2408)
);

HB1xp67_ASAP7_75t_L g2409 ( 
.A(n_2359),
.Y(n_2409)
);

AOI22xp33_ASAP7_75t_L g2410 ( 
.A1(n_2297),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2348),
.Y(n_2411)
);

AND2x2_ASAP7_75t_L g2412 ( 
.A(n_2310),
.B(n_161),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_2312),
.B(n_162),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2313),
.Y(n_2414)
);

OAI221xp5_ASAP7_75t_SL g2415 ( 
.A1(n_2373),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.C(n_166),
.Y(n_2415)
);

AND2x4_ASAP7_75t_L g2416 ( 
.A(n_2330),
.B(n_163),
.Y(n_2416)
);

NOR2xp67_ASAP7_75t_L g2417 ( 
.A(n_2362),
.B(n_165),
.Y(n_2417)
);

NOR2xp67_ASAP7_75t_L g2418 ( 
.A(n_2362),
.B(n_167),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2364),
.B(n_167),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2384),
.B(n_168),
.Y(n_2420)
);

INVxp67_ASAP7_75t_SL g2421 ( 
.A(n_2313),
.Y(n_2421)
);

AND2x4_ASAP7_75t_L g2422 ( 
.A(n_2362),
.B(n_168),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2340),
.Y(n_2423)
);

INVxp67_ASAP7_75t_L g2424 ( 
.A(n_2353),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_2350),
.B(n_169),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2331),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2304),
.B(n_170),
.Y(n_2427)
);

HB1xp67_ASAP7_75t_L g2428 ( 
.A(n_2331),
.Y(n_2428)
);

OAI211xp5_ASAP7_75t_L g2429 ( 
.A1(n_2306),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_2429)
);

INVx3_ASAP7_75t_L g2430 ( 
.A(n_2338),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2304),
.B(n_171),
.Y(n_2431)
);

AND2x2_ASAP7_75t_L g2432 ( 
.A(n_2307),
.B(n_173),
.Y(n_2432)
);

AND2x4_ASAP7_75t_L g2433 ( 
.A(n_2361),
.B(n_173),
.Y(n_2433)
);

BUFx3_ASAP7_75t_L g2434 ( 
.A(n_2363),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_2381),
.B(n_174),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2382),
.B(n_174),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2349),
.B(n_175),
.Y(n_2437)
);

AND2x4_ASAP7_75t_SL g2438 ( 
.A(n_2315),
.B(n_2300),
.Y(n_2438)
);

INVx3_ASAP7_75t_L g2439 ( 
.A(n_2355),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2367),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2380),
.B(n_175),
.Y(n_2441)
);

NOR2xp33_ASAP7_75t_L g2442 ( 
.A(n_2303),
.B(n_176),
.Y(n_2442)
);

HB1xp67_ASAP7_75t_L g2443 ( 
.A(n_2298),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2358),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2301),
.B(n_2319),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2336),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2369),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2314),
.B(n_176),
.Y(n_2448)
);

AND2x2_ASAP7_75t_L g2449 ( 
.A(n_2327),
.B(n_2316),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2383),
.B(n_177),
.Y(n_2450)
);

BUFx2_ASAP7_75t_L g2451 ( 
.A(n_2366),
.Y(n_2451)
);

BUFx3_ASAP7_75t_L g2452 ( 
.A(n_2376),
.Y(n_2452)
);

INVxp67_ASAP7_75t_L g2453 ( 
.A(n_2328),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2385),
.Y(n_2454)
);

BUFx2_ASAP7_75t_L g2455 ( 
.A(n_2334),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2370),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2371),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2324),
.Y(n_2458)
);

OAI22xp5_ASAP7_75t_L g2459 ( 
.A1(n_2379),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2311),
.Y(n_2460)
);

OR2x2_ASAP7_75t_L g2461 ( 
.A(n_2372),
.B(n_179),
.Y(n_2461)
);

HB1xp67_ASAP7_75t_L g2462 ( 
.A(n_2320),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2342),
.Y(n_2463)
);

HB1xp67_ASAP7_75t_L g2464 ( 
.A(n_2337),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_2343),
.B(n_181),
.Y(n_2465)
);

OR2x2_ASAP7_75t_L g2466 ( 
.A(n_2344),
.B(n_181),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2378),
.B(n_182),
.Y(n_2467)
);

BUFx2_ASAP7_75t_L g2468 ( 
.A(n_2388),
.Y(n_2468)
);

INVx1_ASAP7_75t_SL g2469 ( 
.A(n_2309),
.Y(n_2469)
);

HB1xp67_ASAP7_75t_L g2470 ( 
.A(n_2321),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_SL g2471 ( 
.A(n_2360),
.B(n_184),
.Y(n_2471)
);

AND2x2_ASAP7_75t_L g2472 ( 
.A(n_2347),
.B(n_185),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2354),
.B(n_185),
.Y(n_2473)
);

NOR2xp33_ASAP7_75t_L g2474 ( 
.A(n_2365),
.B(n_186),
.Y(n_2474)
);

OR2x2_ASAP7_75t_L g2475 ( 
.A(n_2329),
.B(n_186),
.Y(n_2475)
);

INVxp67_ASAP7_75t_SL g2476 ( 
.A(n_2302),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2335),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2377),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2386),
.Y(n_2479)
);

NOR2xp33_ASAP7_75t_L g2480 ( 
.A(n_2387),
.B(n_187),
.Y(n_2480)
);

INVxp67_ASAP7_75t_SL g2481 ( 
.A(n_2374),
.Y(n_2481)
);

NAND2xp33_ASAP7_75t_L g2482 ( 
.A(n_2362),
.B(n_188),
.Y(n_2482)
);

AND2x2_ASAP7_75t_L g2483 ( 
.A(n_2357),
.B(n_189),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2356),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2356),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2356),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2356),
.Y(n_2487)
);

AND2x2_ASAP7_75t_L g2488 ( 
.A(n_2357),
.B(n_191),
.Y(n_2488)
);

INVx5_ASAP7_75t_L g2489 ( 
.A(n_2304),
.Y(n_2489)
);

AND2x4_ASAP7_75t_L g2490 ( 
.A(n_2326),
.B(n_191),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2339),
.B(n_192),
.Y(n_2491)
);

AND2x4_ASAP7_75t_L g2492 ( 
.A(n_2326),
.B(n_193),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2356),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2356),
.Y(n_2494)
);

AND2x4_ASAP7_75t_L g2495 ( 
.A(n_2326),
.B(n_195),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2357),
.B(n_195),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2356),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_2357),
.B(n_196),
.Y(n_2498)
);

HB1xp67_ASAP7_75t_L g2499 ( 
.A(n_2339),
.Y(n_2499)
);

OR2x2_ASAP7_75t_L g2500 ( 
.A(n_2339),
.B(n_196),
.Y(n_2500)
);

HB1xp67_ASAP7_75t_L g2501 ( 
.A(n_2339),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2357),
.B(n_197),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2356),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2356),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2356),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2356),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2390),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2443),
.B(n_197),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2393),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2397),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2392),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2400),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2499),
.B(n_198),
.Y(n_2513)
);

AND2x2_ASAP7_75t_L g2514 ( 
.A(n_2389),
.B(n_199),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2401),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2484),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2486),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2487),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2501),
.B(n_201),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2440),
.B(n_2423),
.Y(n_2520)
);

AND2x4_ASAP7_75t_L g2521 ( 
.A(n_2404),
.B(n_203),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2494),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2409),
.B(n_203),
.Y(n_2523)
);

NAND2x1_ASAP7_75t_L g2524 ( 
.A(n_2414),
.B(n_205),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2497),
.Y(n_2525)
);

NAND3xp33_ASAP7_75t_L g2526 ( 
.A(n_2464),
.B(n_2451),
.C(n_2453),
.Y(n_2526)
);

OR2x2_ASAP7_75t_L g2527 ( 
.A(n_2408),
.B(n_204),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2394),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2424),
.B(n_206),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2398),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2485),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2434),
.B(n_206),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2493),
.Y(n_2533)
);

AND2x4_ASAP7_75t_L g2534 ( 
.A(n_2403),
.B(n_207),
.Y(n_2534)
);

OR2x2_ASAP7_75t_L g2535 ( 
.A(n_2407),
.B(n_207),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2411),
.B(n_208),
.Y(n_2536)
);

AND2x2_ASAP7_75t_L g2537 ( 
.A(n_2430),
.B(n_208),
.Y(n_2537)
);

INVxp67_ASAP7_75t_SL g2538 ( 
.A(n_2417),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2503),
.Y(n_2539)
);

NAND2x1_ASAP7_75t_L g2540 ( 
.A(n_2426),
.B(n_210),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2506),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2399),
.B(n_209),
.Y(n_2542)
);

HB1xp67_ASAP7_75t_L g2543 ( 
.A(n_2428),
.Y(n_2543)
);

OR2x2_ASAP7_75t_L g2544 ( 
.A(n_2421),
.B(n_211),
.Y(n_2544)
);

AND2x4_ASAP7_75t_L g2545 ( 
.A(n_2489),
.B(n_212),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2489),
.B(n_212),
.Y(n_2546)
);

AND2x4_ASAP7_75t_L g2547 ( 
.A(n_2489),
.B(n_213),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2444),
.B(n_213),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2504),
.Y(n_2549)
);

AND2x4_ASAP7_75t_L g2550 ( 
.A(n_2422),
.B(n_214),
.Y(n_2550)
);

AND2x2_ASAP7_75t_L g2551 ( 
.A(n_2462),
.B(n_214),
.Y(n_2551)
);

NAND2xp33_ASAP7_75t_L g2552 ( 
.A(n_2395),
.B(n_215),
.Y(n_2552)
);

AND2x4_ASAP7_75t_L g2553 ( 
.A(n_2418),
.B(n_215),
.Y(n_2553)
);

INVx3_ASAP7_75t_L g2554 ( 
.A(n_2490),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2446),
.B(n_216),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2505),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2402),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2391),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2406),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2468),
.B(n_216),
.Y(n_2560)
);

OR2x2_ASAP7_75t_L g2561 ( 
.A(n_2500),
.B(n_217),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2483),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2416),
.B(n_218),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2447),
.B(n_218),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2454),
.B(n_219),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2455),
.B(n_219),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2488),
.Y(n_2567)
);

HB1xp67_ASAP7_75t_L g2568 ( 
.A(n_2470),
.Y(n_2568)
);

AND2x2_ASAP7_75t_L g2569 ( 
.A(n_2452),
.B(n_220),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2491),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2396),
.B(n_220),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2405),
.B(n_221),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2496),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2460),
.B(n_221),
.Y(n_2574)
);

OR2x2_ASAP7_75t_L g2575 ( 
.A(n_2477),
.B(n_222),
.Y(n_2575)
);

BUFx2_ASAP7_75t_L g2576 ( 
.A(n_2476),
.Y(n_2576)
);

AND2x4_ASAP7_75t_L g2577 ( 
.A(n_2498),
.B(n_223),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2502),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2432),
.B(n_223),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2442),
.B(n_224),
.Y(n_2580)
);

HB1xp67_ASAP7_75t_L g2581 ( 
.A(n_2441),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_2435),
.B(n_224),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2437),
.Y(n_2583)
);

NOR2xp67_ASAP7_75t_L g2584 ( 
.A(n_2492),
.B(n_225),
.Y(n_2584)
);

INVxp67_ASAP7_75t_SL g2585 ( 
.A(n_2482),
.Y(n_2585)
);

NAND3xp33_ASAP7_75t_L g2586 ( 
.A(n_2459),
.B(n_2457),
.C(n_2456),
.Y(n_2586)
);

HB1xp67_ASAP7_75t_L g2587 ( 
.A(n_2433),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_SL g2588 ( 
.A(n_2481),
.B(n_225),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2463),
.B(n_226),
.Y(n_2589)
);

NOR3xp33_ASAP7_75t_SL g2590 ( 
.A(n_2429),
.B(n_227),
.C(n_228),
.Y(n_2590)
);

OR2x2_ASAP7_75t_L g2591 ( 
.A(n_2419),
.B(n_227),
.Y(n_2591)
);

OR2x2_ASAP7_75t_L g2592 ( 
.A(n_2479),
.B(n_228),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2412),
.Y(n_2593)
);

INVxp67_ASAP7_75t_L g2594 ( 
.A(n_2427),
.Y(n_2594)
);

NAND2x1_ASAP7_75t_SL g2595 ( 
.A(n_2495),
.B(n_229),
.Y(n_2595)
);

AND2x2_ASAP7_75t_L g2596 ( 
.A(n_2436),
.B(n_2413),
.Y(n_2596)
);

NOR2xp33_ASAP7_75t_L g2597 ( 
.A(n_2458),
.B(n_229),
.Y(n_2597)
);

OR2x2_ASAP7_75t_L g2598 ( 
.A(n_2469),
.B(n_230),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2445),
.B(n_230),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2431),
.Y(n_2600)
);

OAI22xp5_ASAP7_75t_L g2601 ( 
.A1(n_2410),
.A2(n_2415),
.B1(n_2449),
.B2(n_2467),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2478),
.Y(n_2602)
);

AND2x4_ASAP7_75t_SL g2603 ( 
.A(n_2425),
.B(n_2420),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2448),
.B(n_231),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2438),
.B(n_231),
.Y(n_2605)
);

INVx3_ASAP7_75t_L g2606 ( 
.A(n_2461),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2466),
.Y(n_2607)
);

OR2x2_ASAP7_75t_L g2608 ( 
.A(n_2450),
.B(n_234),
.Y(n_2608)
);

OAI21xp5_ASAP7_75t_SL g2609 ( 
.A1(n_2474),
.A2(n_234),
.B(n_235),
.Y(n_2609)
);

HB1xp67_ASAP7_75t_L g2610 ( 
.A(n_2465),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2472),
.B(n_235),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2475),
.Y(n_2612)
);

OR2x2_ASAP7_75t_L g2613 ( 
.A(n_2473),
.B(n_236),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2480),
.B(n_236),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_L g2615 ( 
.A(n_2471),
.B(n_237),
.Y(n_2615)
);

INVxp67_ASAP7_75t_L g2616 ( 
.A(n_2443),
.Y(n_2616)
);

BUFx2_ASAP7_75t_L g2617 ( 
.A(n_2428),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2443),
.B(n_237),
.Y(n_2618)
);

HB1xp67_ASAP7_75t_L g2619 ( 
.A(n_2428),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2439),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2389),
.B(n_238),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2439),
.Y(n_2622)
);

OR2x2_ASAP7_75t_L g2623 ( 
.A(n_2408),
.B(n_238),
.Y(n_2623)
);

BUFx3_ASAP7_75t_L g2624 ( 
.A(n_2403),
.Y(n_2624)
);

OR2x2_ASAP7_75t_L g2625 ( 
.A(n_2408),
.B(n_239),
.Y(n_2625)
);

AND2x4_ASAP7_75t_L g2626 ( 
.A(n_2404),
.B(n_239),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2389),
.B(n_240),
.Y(n_2627)
);

OR2x2_ASAP7_75t_L g2628 ( 
.A(n_2408),
.B(n_240),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2390),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2443),
.B(n_241),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2389),
.B(n_241),
.Y(n_2631)
);

AND2x2_ASAP7_75t_L g2632 ( 
.A(n_2389),
.B(n_242),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2439),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2443),
.B(n_242),
.Y(n_2634)
);

OR2x2_ASAP7_75t_L g2635 ( 
.A(n_2408),
.B(n_243),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2390),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2443),
.B(n_243),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2390),
.Y(n_2638)
);

AND2x4_ASAP7_75t_SL g2639 ( 
.A(n_2404),
.B(n_244),
.Y(n_2639)
);

OR2x2_ASAP7_75t_L g2640 ( 
.A(n_2408),
.B(n_244),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2390),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2389),
.B(n_245),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2389),
.B(n_245),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2390),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2390),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2443),
.B(n_247),
.Y(n_2646)
);

OR2x2_ASAP7_75t_L g2647 ( 
.A(n_2408),
.B(n_248),
.Y(n_2647)
);

NOR2xp33_ASAP7_75t_L g2648 ( 
.A(n_2403),
.B(n_248),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2389),
.B(n_249),
.Y(n_2649)
);

INVxp33_ASAP7_75t_SL g2650 ( 
.A(n_2403),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2390),
.Y(n_2651)
);

OR2x2_ASAP7_75t_L g2652 ( 
.A(n_2408),
.B(n_249),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2443),
.B(n_250),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2389),
.B(n_250),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2390),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2439),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2439),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2389),
.B(n_251),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2389),
.B(n_251),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2390),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2389),
.B(n_252),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2443),
.B(n_253),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2390),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2390),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2390),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2389),
.B(n_253),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2390),
.Y(n_2667)
);

OR2x2_ASAP7_75t_L g2668 ( 
.A(n_2616),
.B(n_254),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2606),
.B(n_2538),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2624),
.B(n_254),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2581),
.B(n_255),
.Y(n_2671)
);

AOI21xp5_ASAP7_75t_SL g2672 ( 
.A1(n_2585),
.A2(n_255),
.B(n_256),
.Y(n_2672)
);

INVx2_ASAP7_75t_SL g2673 ( 
.A(n_2545),
.Y(n_2673)
);

OAI21xp5_ASAP7_75t_L g2674 ( 
.A1(n_2526),
.A2(n_257),
.B(n_258),
.Y(n_2674)
);

OAI321xp33_ASAP7_75t_L g2675 ( 
.A1(n_2601),
.A2(n_261),
.A3(n_263),
.B1(n_259),
.B2(n_260),
.C(n_262),
.Y(n_2675)
);

OR2x2_ASAP7_75t_L g2676 ( 
.A(n_2602),
.B(n_263),
.Y(n_2676)
);

OAI221xp5_ASAP7_75t_L g2677 ( 
.A1(n_2609),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.C(n_267),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2617),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2617),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2557),
.B(n_264),
.Y(n_2680)
);

OAI22xp5_ASAP7_75t_L g2681 ( 
.A1(n_2590),
.A2(n_2650),
.B1(n_2586),
.B2(n_2576),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2620),
.Y(n_2682)
);

AOI33xp33_ASAP7_75t_L g2683 ( 
.A1(n_2566),
.A2(n_267),
.A3(n_269),
.B1(n_265),
.B2(n_266),
.B3(n_268),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2507),
.Y(n_2684)
);

INVxp67_ASAP7_75t_SL g2685 ( 
.A(n_2568),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2509),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2622),
.B(n_268),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2510),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2633),
.B(n_270),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2656),
.Y(n_2690)
);

INVxp67_ASAP7_75t_SL g2691 ( 
.A(n_2595),
.Y(n_2691)
);

OAI33xp33_ASAP7_75t_L g2692 ( 
.A1(n_2560),
.A2(n_272),
.A3(n_274),
.B1(n_270),
.B2(n_271),
.B3(n_273),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2512),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2594),
.B(n_2558),
.Y(n_2694)
);

OAI22xp5_ASAP7_75t_L g2695 ( 
.A1(n_2576),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.Y(n_2695)
);

OR2x2_ASAP7_75t_L g2696 ( 
.A(n_2520),
.B(n_275),
.Y(n_2696)
);

OAI33xp33_ASAP7_75t_L g2697 ( 
.A1(n_2580),
.A2(n_278),
.A3(n_280),
.B1(n_276),
.B2(n_277),
.B3(n_279),
.Y(n_2697)
);

BUFx3_ASAP7_75t_L g2698 ( 
.A(n_2639),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2657),
.B(n_2607),
.Y(n_2699)
);

AOI221xp5_ASAP7_75t_L g2700 ( 
.A1(n_2588),
.A2(n_282),
.B1(n_279),
.B2(n_281),
.C(n_283),
.Y(n_2700)
);

NOR2xp33_ASAP7_75t_SL g2701 ( 
.A(n_2584),
.B(n_281),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2600),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2562),
.Y(n_2703)
);

OR2x2_ASAP7_75t_L g2704 ( 
.A(n_2583),
.B(n_282),
.Y(n_2704)
);

AOI21xp5_ASAP7_75t_SL g2705 ( 
.A1(n_2553),
.A2(n_283),
.B(n_284),
.Y(n_2705)
);

NAND5xp2_ASAP7_75t_L g2706 ( 
.A(n_2648),
.B(n_287),
.C(n_285),
.D(n_286),
.E(n_288),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2515),
.Y(n_2707)
);

INVx2_ASAP7_75t_SL g2708 ( 
.A(n_2547),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2567),
.Y(n_2709)
);

BUFx2_ASAP7_75t_L g2710 ( 
.A(n_2587),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2516),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2573),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2610),
.B(n_285),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2570),
.B(n_287),
.Y(n_2714)
);

OAI31xp33_ASAP7_75t_SL g2715 ( 
.A1(n_2551),
.A2(n_291),
.A3(n_292),
.B(n_290),
.Y(n_2715)
);

INVx5_ASAP7_75t_L g2716 ( 
.A(n_2546),
.Y(n_2716)
);

HB1xp67_ASAP7_75t_L g2717 ( 
.A(n_2543),
.Y(n_2717)
);

NAND4xp25_ASAP7_75t_L g2718 ( 
.A(n_2597),
.B(n_292),
.C(n_293),
.D(n_290),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2514),
.B(n_289),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2517),
.Y(n_2720)
);

OR2x2_ASAP7_75t_L g2721 ( 
.A(n_2612),
.B(n_289),
.Y(n_2721)
);

AND2x2_ASAP7_75t_L g2722 ( 
.A(n_2578),
.B(n_293),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2518),
.Y(n_2723)
);

AND2x2_ASAP7_75t_L g2724 ( 
.A(n_2559),
.B(n_294),
.Y(n_2724)
);

NAND2x1_ASAP7_75t_L g2725 ( 
.A(n_2531),
.B(n_2533),
.Y(n_2725)
);

BUFx2_ASAP7_75t_L g2726 ( 
.A(n_2619),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2522),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2593),
.Y(n_2728)
);

OAI221xp5_ASAP7_75t_L g2729 ( 
.A1(n_2552),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.C(n_298),
.Y(n_2729)
);

NOR2xp33_ASAP7_75t_L g2730 ( 
.A(n_2508),
.B(n_295),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2596),
.B(n_297),
.Y(n_2731)
);

NAND3xp33_ASAP7_75t_L g2732 ( 
.A(n_2618),
.B(n_298),
.C(n_299),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2525),
.Y(n_2733)
);

INVx3_ASAP7_75t_L g2734 ( 
.A(n_2554),
.Y(n_2734)
);

INVxp67_ASAP7_75t_L g2735 ( 
.A(n_2544),
.Y(n_2735)
);

AOI33xp33_ASAP7_75t_L g2736 ( 
.A1(n_2614),
.A2(n_301),
.A3(n_303),
.B1(n_299),
.B2(n_300),
.B3(n_302),
.Y(n_2736)
);

NOR2xp67_ASAP7_75t_L g2737 ( 
.A(n_2541),
.B(n_303),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2511),
.Y(n_2738)
);

NOR2x1_ASAP7_75t_L g2739 ( 
.A(n_2524),
.B(n_304),
.Y(n_2739)
);

NAND4xp25_ASAP7_75t_L g2740 ( 
.A(n_2599),
.B(n_2634),
.C(n_2637),
.D(n_2630),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2539),
.Y(n_2741)
);

INVxp67_ASAP7_75t_SL g2742 ( 
.A(n_2540),
.Y(n_2742)
);

NOR3xp33_ASAP7_75t_L g2743 ( 
.A(n_2646),
.B(n_304),
.C(n_305),
.Y(n_2743)
);

NOR2xp67_ASAP7_75t_L g2744 ( 
.A(n_2549),
.B(n_305),
.Y(n_2744)
);

OAI221xp5_ASAP7_75t_SL g2745 ( 
.A1(n_2653),
.A2(n_2662),
.B1(n_2615),
.B2(n_2598),
.C(n_2608),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2621),
.B(n_306),
.Y(n_2746)
);

AND2x4_ASAP7_75t_L g2747 ( 
.A(n_2603),
.B(n_307),
.Y(n_2747)
);

AOI221xp5_ASAP7_75t_L g2748 ( 
.A1(n_2589),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.C(n_310),
.Y(n_2748)
);

AOI22xp5_ASAP7_75t_L g2749 ( 
.A1(n_2627),
.A2(n_311),
.B1(n_308),
.B2(n_310),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2556),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2528),
.Y(n_2751)
);

OR2x2_ASAP7_75t_L g2752 ( 
.A(n_2530),
.B(n_311),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2631),
.B(n_2666),
.Y(n_2753)
);

OR2x2_ASAP7_75t_L g2754 ( 
.A(n_2629),
.B(n_312),
.Y(n_2754)
);

HB1xp67_ASAP7_75t_L g2755 ( 
.A(n_2636),
.Y(n_2755)
);

INVx3_ASAP7_75t_L g2756 ( 
.A(n_2534),
.Y(n_2756)
);

INVx2_ASAP7_75t_SL g2757 ( 
.A(n_2521),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2632),
.B(n_313),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2638),
.Y(n_2759)
);

BUFx2_ASAP7_75t_L g2760 ( 
.A(n_2626),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2641),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2642),
.B(n_313),
.Y(n_2762)
);

AND2x4_ASAP7_75t_L g2763 ( 
.A(n_2537),
.B(n_314),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2643),
.B(n_314),
.Y(n_2764)
);

AND2x2_ASAP7_75t_L g2765 ( 
.A(n_2649),
.B(n_315),
.Y(n_2765)
);

AOI21xp5_ASAP7_75t_L g2766 ( 
.A1(n_2605),
.A2(n_315),
.B(n_316),
.Y(n_2766)
);

OAI221xp5_ASAP7_75t_L g2767 ( 
.A1(n_2548),
.A2(n_320),
.B1(n_317),
.B2(n_319),
.C(n_321),
.Y(n_2767)
);

AO21x2_ASAP7_75t_L g2768 ( 
.A1(n_2513),
.A2(n_2519),
.B(n_2542),
.Y(n_2768)
);

AND2x2_ASAP7_75t_L g2769 ( 
.A(n_2654),
.B(n_317),
.Y(n_2769)
);

OAI21x1_ASAP7_75t_L g2770 ( 
.A1(n_2644),
.A2(n_2651),
.B(n_2645),
.Y(n_2770)
);

OAI22xp5_ASAP7_75t_L g2771 ( 
.A1(n_2555),
.A2(n_2592),
.B1(n_2613),
.B2(n_2575),
.Y(n_2771)
);

AOI221xp5_ASAP7_75t_L g2772 ( 
.A1(n_2604),
.A2(n_322),
.B1(n_319),
.B2(n_320),
.C(n_323),
.Y(n_2772)
);

NOR2x1_ASAP7_75t_L g2773 ( 
.A(n_2658),
.B(n_323),
.Y(n_2773)
);

AOI221xp5_ASAP7_75t_L g2774 ( 
.A1(n_2569),
.A2(n_327),
.B1(n_324),
.B2(n_326),
.C(n_328),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2655),
.Y(n_2775)
);

NAND3xp33_ASAP7_75t_L g2776 ( 
.A(n_2571),
.B(n_324),
.C(n_326),
.Y(n_2776)
);

BUFx2_ASAP7_75t_L g2777 ( 
.A(n_2659),
.Y(n_2777)
);

OR2x2_ASAP7_75t_L g2778 ( 
.A(n_2660),
.B(n_327),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2661),
.B(n_328),
.Y(n_2779)
);

AOI22xp5_ASAP7_75t_L g2780 ( 
.A1(n_2574),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_2780)
);

OR2x2_ASAP7_75t_L g2781 ( 
.A(n_2663),
.B(n_330),
.Y(n_2781)
);

NOR2xp33_ASAP7_75t_L g2782 ( 
.A(n_2673),
.B(n_2591),
.Y(n_2782)
);

NOR2x1_ASAP7_75t_L g2783 ( 
.A(n_2672),
.B(n_2535),
.Y(n_2783)
);

AND2x2_ASAP7_75t_L g2784 ( 
.A(n_2716),
.B(n_2564),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2756),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2691),
.B(n_2565),
.Y(n_2786)
);

NOR2xp33_ASAP7_75t_L g2787 ( 
.A(n_2708),
.B(n_2572),
.Y(n_2787)
);

INVx1_ASAP7_75t_SL g2788 ( 
.A(n_2698),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2716),
.B(n_2523),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2716),
.B(n_2529),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2717),
.Y(n_2791)
);

OAI21xp5_ASAP7_75t_L g2792 ( 
.A1(n_2681),
.A2(n_2611),
.B(n_2563),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2710),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2777),
.B(n_2579),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2760),
.Y(n_2795)
);

AND2x2_ASAP7_75t_L g2796 ( 
.A(n_2734),
.B(n_2582),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2742),
.B(n_2532),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2757),
.Y(n_2798)
);

NAND3xp33_ASAP7_75t_SL g2799 ( 
.A(n_2674),
.B(n_2623),
.C(n_2527),
.Y(n_2799)
);

AND2x2_ASAP7_75t_L g2800 ( 
.A(n_2699),
.B(n_2536),
.Y(n_2800)
);

INVx1_ASAP7_75t_SL g2801 ( 
.A(n_2747),
.Y(n_2801)
);

OR2x2_ASAP7_75t_L g2802 ( 
.A(n_2669),
.B(n_2625),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2715),
.B(n_2628),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2726),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2735),
.B(n_2635),
.Y(n_2805)
);

AND2x2_ASAP7_75t_L g2806 ( 
.A(n_2768),
.B(n_2664),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2703),
.B(n_2665),
.Y(n_2807)
);

AND2x4_ASAP7_75t_L g2808 ( 
.A(n_2685),
.B(n_2667),
.Y(n_2808)
);

OR2x2_ASAP7_75t_L g2809 ( 
.A(n_2694),
.B(n_2709),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2771),
.B(n_2640),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2712),
.B(n_2577),
.Y(n_2811)
);

AOI22xp33_ASAP7_75t_L g2812 ( 
.A1(n_2743),
.A2(n_2647),
.B1(n_2652),
.B2(n_2550),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2755),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2744),
.B(n_2561),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2678),
.Y(n_2815)
);

OR2x2_ASAP7_75t_L g2816 ( 
.A(n_2702),
.B(n_332),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2679),
.Y(n_2817)
);

INVxp67_ASAP7_75t_L g2818 ( 
.A(n_2701),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2684),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2753),
.B(n_332),
.Y(n_2820)
);

INVx1_ASAP7_75t_SL g2821 ( 
.A(n_2773),
.Y(n_2821)
);

OAI21xp33_ASAP7_75t_L g2822 ( 
.A1(n_2706),
.A2(n_333),
.B(n_334),
.Y(n_2822)
);

AND2x4_ASAP7_75t_L g2823 ( 
.A(n_2687),
.B(n_333),
.Y(n_2823)
);

INVx2_ASAP7_75t_SL g2824 ( 
.A(n_2725),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2686),
.Y(n_2825)
);

O2A1O1Ixp33_ASAP7_75t_L g2826 ( 
.A1(n_2675),
.A2(n_336),
.B(n_334),
.C(n_335),
.Y(n_2826)
);

OR2x2_ASAP7_75t_L g2827 ( 
.A(n_2728),
.B(n_2740),
.Y(n_2827)
);

AND2x2_ASAP7_75t_L g2828 ( 
.A(n_2682),
.B(n_2690),
.Y(n_2828)
);

INVxp67_ASAP7_75t_SL g2829 ( 
.A(n_2737),
.Y(n_2829)
);

OR2x2_ASAP7_75t_L g2830 ( 
.A(n_2696),
.B(n_337),
.Y(n_2830)
);

INVx1_ASAP7_75t_SL g2831 ( 
.A(n_2739),
.Y(n_2831)
);

INVx1_ASAP7_75t_SL g2832 ( 
.A(n_2670),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2752),
.Y(n_2833)
);

AND2x4_ASAP7_75t_L g2834 ( 
.A(n_2689),
.B(n_337),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_SL g2835 ( 
.A(n_2683),
.B(n_338),
.Y(n_2835)
);

OR2x2_ASAP7_75t_L g2836 ( 
.A(n_2738),
.B(n_338),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2688),
.Y(n_2837)
);

OR2x2_ASAP7_75t_L g2838 ( 
.A(n_2751),
.B(n_339),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2831),
.B(n_2766),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2821),
.B(n_2671),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2788),
.B(n_2731),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2791),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2829),
.B(n_2713),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2789),
.B(n_2746),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2795),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2824),
.Y(n_2846)
);

OR2x2_ASAP7_75t_L g2847 ( 
.A(n_2793),
.B(n_2745),
.Y(n_2847)
);

AND2x2_ASAP7_75t_L g2848 ( 
.A(n_2797),
.B(n_2758),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2801),
.B(n_2794),
.Y(n_2849)
);

INVx3_ASAP7_75t_SL g2850 ( 
.A(n_2823),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2836),
.Y(n_2851)
);

NOR2x1_ASAP7_75t_L g2852 ( 
.A(n_2783),
.B(n_2705),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2838),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2816),
.Y(n_2854)
);

AND2x2_ASAP7_75t_L g2855 ( 
.A(n_2784),
.B(n_2765),
.Y(n_2855)
);

INVx2_ASAP7_75t_SL g2856 ( 
.A(n_2804),
.Y(n_2856)
);

AND2x2_ASAP7_75t_L g2857 ( 
.A(n_2796),
.B(n_2769),
.Y(n_2857)
);

AND2x2_ASAP7_75t_L g2858 ( 
.A(n_2800),
.B(n_2779),
.Y(n_2858)
);

INVx1_ASAP7_75t_SL g2859 ( 
.A(n_2832),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2815),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2817),
.Y(n_2861)
);

OR2x2_ASAP7_75t_L g2862 ( 
.A(n_2827),
.B(n_2721),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2818),
.B(n_2798),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2785),
.B(n_2680),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2811),
.Y(n_2865)
);

OR2x2_ASAP7_75t_L g2866 ( 
.A(n_2810),
.B(n_2668),
.Y(n_2866)
);

AND2x2_ASAP7_75t_L g2867 ( 
.A(n_2833),
.B(n_2762),
.Y(n_2867)
);

AND2x2_ASAP7_75t_L g2868 ( 
.A(n_2782),
.B(n_2764),
.Y(n_2868)
);

INVxp67_ASAP7_75t_L g2869 ( 
.A(n_2814),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2813),
.Y(n_2870)
);

NOR2xp33_ASAP7_75t_L g2871 ( 
.A(n_2850),
.B(n_2803),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2841),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2867),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2849),
.Y(n_2874)
);

A2O1A1Ixp33_ASAP7_75t_L g2875 ( 
.A1(n_2852),
.A2(n_2826),
.B(n_2822),
.C(n_2792),
.Y(n_2875)
);

AND2x4_ASAP7_75t_L g2876 ( 
.A(n_2855),
.B(n_2790),
.Y(n_2876)
);

OAI21xp5_ASAP7_75t_L g2877 ( 
.A1(n_2839),
.A2(n_2835),
.B(n_2806),
.Y(n_2877)
);

INVx2_ASAP7_75t_SL g2878 ( 
.A(n_2844),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2846),
.Y(n_2879)
);

OAI22xp5_ASAP7_75t_L g2880 ( 
.A1(n_2847),
.A2(n_2677),
.B1(n_2786),
.B2(n_2812),
.Y(n_2880)
);

OAI22xp33_ASAP7_75t_L g2881 ( 
.A1(n_2859),
.A2(n_2718),
.B1(n_2767),
.B2(n_2729),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2851),
.Y(n_2882)
);

INVxp67_ASAP7_75t_L g2883 ( 
.A(n_2848),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2857),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2858),
.B(n_2856),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2845),
.B(n_2787),
.Y(n_2886)
);

AOI22xp33_ASAP7_75t_SL g2887 ( 
.A1(n_2843),
.A2(n_2732),
.B1(n_2776),
.B2(n_2695),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2869),
.B(n_2808),
.Y(n_2888)
);

AND2x2_ASAP7_75t_L g2889 ( 
.A(n_2868),
.B(n_2828),
.Y(n_2889)
);

INVx1_ASAP7_75t_SL g2890 ( 
.A(n_2840),
.Y(n_2890)
);

OAI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2875),
.A2(n_2863),
.B(n_2864),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2873),
.Y(n_2892)
);

OAI22xp5_ASAP7_75t_L g2893 ( 
.A1(n_2887),
.A2(n_2866),
.B1(n_2862),
.B2(n_2802),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2878),
.B(n_2865),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2872),
.Y(n_2895)
);

AOI322xp5_ASAP7_75t_L g2896 ( 
.A1(n_2881),
.A2(n_2842),
.A3(n_2799),
.B1(n_2870),
.B2(n_2860),
.C1(n_2861),
.C2(n_2730),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2876),
.Y(n_2897)
);

NOR2x1_ASAP7_75t_SL g2898 ( 
.A(n_2889),
.B(n_2853),
.Y(n_2898)
);

OAI211xp5_ASAP7_75t_L g2899 ( 
.A1(n_2877),
.A2(n_2772),
.B(n_2748),
.C(n_2774),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2883),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2898),
.B(n_2871),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2894),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2897),
.B(n_2890),
.Y(n_2903)
);

OR2x2_ASAP7_75t_L g2904 ( 
.A(n_2893),
.B(n_2884),
.Y(n_2904)
);

AOI22xp5_ASAP7_75t_L g2905 ( 
.A1(n_2899),
.A2(n_2880),
.B1(n_2874),
.B2(n_2885),
.Y(n_2905)
);

AOI22xp33_ASAP7_75t_L g2906 ( 
.A1(n_2891),
.A2(n_2879),
.B1(n_2886),
.B2(n_2854),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2895),
.Y(n_2907)
);

AOI22xp33_ASAP7_75t_SL g2908 ( 
.A1(n_2900),
.A2(n_2888),
.B1(n_2882),
.B2(n_2870),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2892),
.Y(n_2909)
);

NOR2xp33_ASAP7_75t_L g2910 ( 
.A(n_2901),
.B(n_2905),
.Y(n_2910)
);

OAI211xp5_ASAP7_75t_SL g2911 ( 
.A1(n_2906),
.A2(n_2896),
.B(n_2820),
.C(n_2805),
.Y(n_2911)
);

NAND4xp25_ASAP7_75t_L g2912 ( 
.A(n_2904),
.B(n_2809),
.C(n_2700),
.D(n_2736),
.Y(n_2912)
);

OAI33xp33_ASAP7_75t_L g2913 ( 
.A1(n_2909),
.A2(n_2819),
.A3(n_2837),
.B1(n_2825),
.B2(n_2830),
.B3(n_2714),
.Y(n_2913)
);

AOI22xp33_ASAP7_75t_SL g2914 ( 
.A1(n_2902),
.A2(n_2903),
.B1(n_2907),
.B2(n_2808),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2908),
.B(n_2834),
.Y(n_2915)
);

OAI321xp33_ASAP7_75t_L g2916 ( 
.A1(n_2905),
.A2(n_2780),
.A3(n_2749),
.B1(n_2676),
.B2(n_2704),
.C(n_2807),
.Y(n_2916)
);

NOR4xp75_ASAP7_75t_SL g2917 ( 
.A(n_2901),
.B(n_2719),
.C(n_2692),
.D(n_2697),
.Y(n_2917)
);

CKINVDCx16_ASAP7_75t_R g2918 ( 
.A(n_2904),
.Y(n_2918)
);

AOI211x1_ASAP7_75t_L g2919 ( 
.A1(n_2901),
.A2(n_2707),
.B(n_2711),
.C(n_2693),
.Y(n_2919)
);

NOR2xp33_ASAP7_75t_L g2920 ( 
.A(n_2901),
.B(n_2778),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2908),
.B(n_2720),
.Y(n_2921)
);

AOI211xp5_ASAP7_75t_L g2922 ( 
.A1(n_2901),
.A2(n_2754),
.B(n_2781),
.C(n_2722),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2903),
.Y(n_2923)
);

OAI221xp5_ASAP7_75t_SL g2924 ( 
.A1(n_2905),
.A2(n_2727),
.B1(n_2741),
.B2(n_2733),
.C(n_2723),
.Y(n_2924)
);

AOI221xp5_ASAP7_75t_L g2925 ( 
.A1(n_2916),
.A2(n_2761),
.B1(n_2775),
.B2(n_2759),
.C(n_2750),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2918),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2915),
.Y(n_2927)
);

NOR2x1_ASAP7_75t_L g2928 ( 
.A(n_2910),
.B(n_2724),
.Y(n_2928)
);

AOI211xp5_ASAP7_75t_SL g2929 ( 
.A1(n_2920),
.A2(n_2763),
.B(n_2770),
.C(n_342),
.Y(n_2929)
);

NAND3xp33_ASAP7_75t_L g2930 ( 
.A(n_2914),
.B(n_340),
.C(n_341),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2921),
.Y(n_2931)
);

AOI22xp5_ASAP7_75t_L g2932 ( 
.A1(n_2911),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_2932)
);

OAI322xp33_ASAP7_75t_L g2933 ( 
.A1(n_2923),
.A2(n_352),
.A3(n_351),
.B1(n_349),
.B2(n_346),
.C1(n_348),
.C2(n_350),
.Y(n_2933)
);

A2O1A1Ixp33_ASAP7_75t_L g2934 ( 
.A1(n_2912),
.A2(n_352),
.B(n_353),
.C(n_351),
.Y(n_2934)
);

AOI221xp5_ASAP7_75t_L g2935 ( 
.A1(n_2924),
.A2(n_354),
.B1(n_356),
.B2(n_353),
.C(n_355),
.Y(n_2935)
);

INVxp67_ASAP7_75t_SL g2936 ( 
.A(n_2922),
.Y(n_2936)
);

NAND4xp75_ASAP7_75t_L g2937 ( 
.A(n_2919),
.B(n_357),
.C(n_350),
.D(n_355),
.Y(n_2937)
);

AOI22xp5_ASAP7_75t_L g2938 ( 
.A1(n_2913),
.A2(n_2917),
.B1(n_361),
.B2(n_359),
.Y(n_2938)
);

OAI211xp5_ASAP7_75t_SL g2939 ( 
.A1(n_2915),
.A2(n_362),
.B(n_359),
.C(n_360),
.Y(n_2939)
);

OAI22xp5_ASAP7_75t_SL g2940 ( 
.A1(n_2918),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2918),
.Y(n_2941)
);

AOI221xp5_ASAP7_75t_L g2942 ( 
.A1(n_2930),
.A2(n_366),
.B1(n_363),
.B2(n_365),
.C(n_367),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2941),
.B(n_2926),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2940),
.Y(n_2944)
);

OAI22xp5_ASAP7_75t_L g2945 ( 
.A1(n_2932),
.A2(n_368),
.B1(n_365),
.B2(n_367),
.Y(n_2945)
);

NAND5xp2_ASAP7_75t_L g2946 ( 
.A(n_2936),
.B(n_384),
.C(n_392),
.D(n_376),
.E(n_368),
.Y(n_2946)
);

OAI21xp33_ASAP7_75t_SL g2947 ( 
.A1(n_2938),
.A2(n_369),
.B(n_370),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2928),
.Y(n_2948)
);

AOI221xp5_ASAP7_75t_L g2949 ( 
.A1(n_2925),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.C(n_374),
.Y(n_2949)
);

INVxp67_ASAP7_75t_L g2950 ( 
.A(n_2937),
.Y(n_2950)
);

AOI21xp5_ASAP7_75t_L g2951 ( 
.A1(n_2929),
.A2(n_371),
.B(n_374),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2927),
.Y(n_2952)
);

OAI211xp5_ASAP7_75t_L g2953 ( 
.A1(n_2935),
.A2(n_385),
.B(n_393),
.C(n_375),
.Y(n_2953)
);

INVxp67_ASAP7_75t_L g2954 ( 
.A(n_2931),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2934),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2933),
.Y(n_2956)
);

AOI211xp5_ASAP7_75t_L g2957 ( 
.A1(n_2939),
.A2(n_380),
.B(n_377),
.C(n_378),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2941),
.Y(n_2958)
);

A2O1A1Ixp33_ASAP7_75t_L g2959 ( 
.A1(n_2951),
.A2(n_2947),
.B(n_2948),
.C(n_2950),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2944),
.Y(n_2960)
);

NOR3xp33_ASAP7_75t_L g2961 ( 
.A(n_2943),
.B(n_387),
.C(n_386),
.Y(n_2961)
);

AOI221x1_ASAP7_75t_SL g2962 ( 
.A1(n_2956),
.A2(n_387),
.B1(n_383),
.B2(n_386),
.C(n_388),
.Y(n_2962)
);

OAI21xp33_ASAP7_75t_SL g2963 ( 
.A1(n_2949),
.A2(n_388),
.B(n_389),
.Y(n_2963)
);

NOR3x1_ASAP7_75t_L g2964 ( 
.A(n_2953),
.B(n_390),
.C(n_391),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2958),
.Y(n_2965)
);

NOR2xp67_ASAP7_75t_L g2966 ( 
.A(n_2946),
.B(n_395),
.Y(n_2966)
);

INVx2_ASAP7_75t_L g2967 ( 
.A(n_2952),
.Y(n_2967)
);

OAI211xp5_ASAP7_75t_SL g2968 ( 
.A1(n_2954),
.A2(n_396),
.B(n_394),
.C(n_395),
.Y(n_2968)
);

AOI22xp5_ASAP7_75t_L g2969 ( 
.A1(n_2955),
.A2(n_398),
.B1(n_394),
.B2(n_397),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2945),
.Y(n_2970)
);

NOR2xp33_ASAP7_75t_L g2971 ( 
.A(n_2942),
.B(n_399),
.Y(n_2971)
);

AOI21xp33_ASAP7_75t_SL g2972 ( 
.A1(n_2948),
.A2(n_400),
.B(n_401),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2950),
.B(n_400),
.Y(n_2973)
);

NOR2x1_ASAP7_75t_L g2974 ( 
.A(n_2948),
.B(n_402),
.Y(n_2974)
);

OAI21xp5_ASAP7_75t_L g2975 ( 
.A1(n_2947),
.A2(n_404),
.B(n_403),
.Y(n_2975)
);

XNOR2x1_ASAP7_75t_L g2976 ( 
.A(n_2958),
.B(n_402),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2943),
.Y(n_2977)
);

AOI22xp33_ASAP7_75t_SL g2978 ( 
.A1(n_2948),
.A2(n_406),
.B1(n_403),
.B2(n_405),
.Y(n_2978)
);

HB1xp67_ASAP7_75t_L g2979 ( 
.A(n_2948),
.Y(n_2979)
);

AND2x2_ASAP7_75t_L g2980 ( 
.A(n_2950),
.B(n_405),
.Y(n_2980)
);

BUFx12f_ASAP7_75t_L g2981 ( 
.A(n_2943),
.Y(n_2981)
);

AOI211xp5_ASAP7_75t_SL g2982 ( 
.A1(n_2950),
.A2(n_409),
.B(n_407),
.C(n_408),
.Y(n_2982)
);

XNOR2x1_ASAP7_75t_L g2983 ( 
.A(n_2958),
.B(n_409),
.Y(n_2983)
);

XNOR2xp5_ASAP7_75t_L g2984 ( 
.A(n_2957),
.B(n_410),
.Y(n_2984)
);

NOR2xp33_ASAP7_75t_L g2985 ( 
.A(n_2950),
.B(n_410),
.Y(n_2985)
);

AO22x1_ASAP7_75t_SL g2986 ( 
.A1(n_2948),
.A2(n_413),
.B1(n_411),
.B2(n_412),
.Y(n_2986)
);

NOR2xp33_ASAP7_75t_L g2987 ( 
.A(n_2950),
.B(n_411),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2943),
.Y(n_2988)
);

INVx1_ASAP7_75t_SL g2989 ( 
.A(n_2948),
.Y(n_2989)
);

O2A1O1Ixp33_ASAP7_75t_L g2990 ( 
.A1(n_2950),
.A2(n_414),
.B(n_412),
.C(n_413),
.Y(n_2990)
);

OR2x2_ASAP7_75t_L g2991 ( 
.A(n_2986),
.B(n_414),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2976),
.Y(n_2992)
);

NAND2x1p5_ASAP7_75t_L g2993 ( 
.A(n_2974),
.B(n_416),
.Y(n_2993)
);

NOR2x1_ASAP7_75t_L g2994 ( 
.A(n_2983),
.B(n_415),
.Y(n_2994)
);

NOR3xp33_ASAP7_75t_L g2995 ( 
.A(n_2959),
.B(n_417),
.C(n_418),
.Y(n_2995)
);

HB1xp67_ASAP7_75t_L g2996 ( 
.A(n_2966),
.Y(n_2996)
);

NOR2x1_ASAP7_75t_L g2997 ( 
.A(n_2968),
.B(n_417),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2980),
.Y(n_2998)
);

HB1xp67_ASAP7_75t_L g2999 ( 
.A(n_2979),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2962),
.B(n_418),
.Y(n_3000)
);

INVx2_ASAP7_75t_SL g3001 ( 
.A(n_2981),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2984),
.Y(n_3002)
);

AND2x2_ASAP7_75t_L g3003 ( 
.A(n_2960),
.B(n_419),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2973),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2985),
.Y(n_3005)
);

NOR2x1_ASAP7_75t_L g3006 ( 
.A(n_2990),
.B(n_2965),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_SL g3007 ( 
.A(n_2978),
.B(n_420),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2967),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2987),
.Y(n_3009)
);

AND3x4_ASAP7_75t_L g3010 ( 
.A(n_2961),
.B(n_420),
.C(n_422),
.Y(n_3010)
);

HB1xp67_ASAP7_75t_L g3011 ( 
.A(n_2964),
.Y(n_3011)
);

AO211x2_ASAP7_75t_L g3012 ( 
.A1(n_2975),
.A2(n_425),
.B(n_422),
.C(n_424),
.Y(n_3012)
);

OAI22xp5_ASAP7_75t_SL g3013 ( 
.A1(n_2989),
.A2(n_428),
.B1(n_424),
.B2(n_427),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2977),
.Y(n_3014)
);

NOR2x1_ASAP7_75t_L g3015 ( 
.A(n_2988),
.B(n_427),
.Y(n_3015)
);

AO22x2_ASAP7_75t_L g3016 ( 
.A1(n_2970),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2982),
.B(n_2972),
.Y(n_3017)
);

INVxp67_ASAP7_75t_SL g3018 ( 
.A(n_2969),
.Y(n_3018)
);

OAI211xp5_ASAP7_75t_SL g3019 ( 
.A1(n_2963),
.A2(n_434),
.B(n_432),
.C(n_433),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2971),
.Y(n_3020)
);

AOI22xp5_ASAP7_75t_L g3021 ( 
.A1(n_2981),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.Y(n_3021)
);

NOR2x1_ASAP7_75t_L g3022 ( 
.A(n_2974),
.B(n_437),
.Y(n_3022)
);

INVx1_ASAP7_75t_SL g3023 ( 
.A(n_2976),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2986),
.Y(n_3024)
);

AOI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_2981),
.A2(n_440),
.B1(n_438),
.B2(n_439),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2986),
.Y(n_3026)
);

XNOR2xp5_ASAP7_75t_L g3027 ( 
.A(n_3012),
.B(n_441),
.Y(n_3027)
);

AND2x2_ASAP7_75t_L g3028 ( 
.A(n_3024),
.B(n_441),
.Y(n_3028)
);

NOR2xp33_ASAP7_75t_L g3029 ( 
.A(n_3019),
.B(n_442),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_3026),
.B(n_442),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2991),
.Y(n_3031)
);

NOR2xp33_ASAP7_75t_L g3032 ( 
.A(n_2996),
.B(n_446),
.Y(n_3032)
);

XNOR2xp5_ASAP7_75t_L g3033 ( 
.A(n_3010),
.B(n_446),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_3011),
.B(n_447),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2993),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_3022),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2999),
.B(n_449),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_3016),
.Y(n_3038)
);

NAND4xp75_ASAP7_75t_L g3039 ( 
.A(n_2994),
.B(n_452),
.C(n_450),
.D(n_451),
.Y(n_3039)
);

HB1xp67_ASAP7_75t_L g3040 ( 
.A(n_3015),
.Y(n_3040)
);

NAND4xp75_ASAP7_75t_L g3041 ( 
.A(n_3006),
.B(n_454),
.C(n_452),
.D(n_453),
.Y(n_3041)
);

HB1xp67_ASAP7_75t_L g3042 ( 
.A(n_3016),
.Y(n_3042)
);

NAND2x1_ASAP7_75t_SL g3043 ( 
.A(n_2997),
.B(n_453),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_3003),
.Y(n_3044)
);

INVx3_ASAP7_75t_L g3045 ( 
.A(n_2998),
.Y(n_3045)
);

NOR2xp67_ASAP7_75t_L g3046 ( 
.A(n_3017),
.B(n_455),
.Y(n_3046)
);

AND2x4_ASAP7_75t_L g3047 ( 
.A(n_3008),
.B(n_454),
.Y(n_3047)
);

XOR2xp5_ASAP7_75t_L g3048 ( 
.A(n_2992),
.B(n_456),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_3013),
.Y(n_3049)
);

XNOR2xp5_ASAP7_75t_L g3050 ( 
.A(n_3023),
.B(n_457),
.Y(n_3050)
);

INVx2_ASAP7_75t_L g3051 ( 
.A(n_3005),
.Y(n_3051)
);

NAND4xp75_ASAP7_75t_L g3052 ( 
.A(n_3000),
.B(n_460),
.C(n_458),
.D(n_459),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_3021),
.Y(n_3053)
);

XNOR2xp5_ASAP7_75t_L g3054 ( 
.A(n_3025),
.B(n_461),
.Y(n_3054)
);

AND2x4_ASAP7_75t_L g3055 ( 
.A(n_3009),
.B(n_462),
.Y(n_3055)
);

NOR2xp67_ASAP7_75t_L g3056 ( 
.A(n_3007),
.B(n_3014),
.Y(n_3056)
);

NOR3xp33_ASAP7_75t_L g3057 ( 
.A(n_3002),
.B(n_472),
.C(n_464),
.Y(n_3057)
);

NOR2x1_ASAP7_75t_L g3058 ( 
.A(n_3004),
.B(n_464),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2995),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_3018),
.Y(n_3060)
);

NOR2xp33_ASAP7_75t_L g3061 ( 
.A(n_3020),
.B(n_466),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_2993),
.Y(n_3062)
);

NAND2x1_ASAP7_75t_L g3063 ( 
.A(n_3022),
.B(n_466),
.Y(n_3063)
);

NOR2xp67_ASAP7_75t_L g3064 ( 
.A(n_2991),
.B(n_469),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2991),
.Y(n_3065)
);

NOR3xp33_ASAP7_75t_L g3066 ( 
.A(n_3001),
.B(n_478),
.C(n_468),
.Y(n_3066)
);

AOI22xp5_ASAP7_75t_L g3067 ( 
.A1(n_3001),
.A2(n_475),
.B1(n_473),
.B2(n_474),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2991),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2991),
.Y(n_3069)
);

NOR2x1_ASAP7_75t_L g3070 ( 
.A(n_3022),
.B(n_475),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2993),
.Y(n_3071)
);

BUFx3_ASAP7_75t_L g3072 ( 
.A(n_2993),
.Y(n_3072)
);

AOI211xp5_ASAP7_75t_L g3073 ( 
.A1(n_3032),
.A2(n_479),
.B(n_477),
.C(n_478),
.Y(n_3073)
);

NOR3xp33_ASAP7_75t_L g3074 ( 
.A(n_3045),
.B(n_481),
.C(n_480),
.Y(n_3074)
);

OAI22x1_ASAP7_75t_L g3075 ( 
.A1(n_3027),
.A2(n_481),
.B1(n_479),
.B2(n_480),
.Y(n_3075)
);

OAI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_3064),
.A2(n_3046),
.B(n_3030),
.Y(n_3076)
);

AOI21xp5_ASAP7_75t_L g3077 ( 
.A1(n_3063),
.A2(n_3070),
.B(n_3036),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_3042),
.B(n_483),
.Y(n_3078)
);

OAI22xp5_ASAP7_75t_L g3079 ( 
.A1(n_3060),
.A2(n_485),
.B1(n_482),
.B2(n_484),
.Y(n_3079)
);

CKINVDCx20_ASAP7_75t_R g3080 ( 
.A(n_3072),
.Y(n_3080)
);

OAI211xp5_ASAP7_75t_L g3081 ( 
.A1(n_3043),
.A2(n_486),
.B(n_484),
.C(n_485),
.Y(n_3081)
);

XNOR2x1_ASAP7_75t_L g3082 ( 
.A(n_3033),
.B(n_486),
.Y(n_3082)
);

O2A1O1Ixp33_ASAP7_75t_L g3083 ( 
.A1(n_3040),
.A2(n_489),
.B(n_487),
.C(n_488),
.Y(n_3083)
);

OAI211xp5_ASAP7_75t_SL g3084 ( 
.A1(n_3031),
.A2(n_492),
.B(n_490),
.C(n_491),
.Y(n_3084)
);

OAI211xp5_ASAP7_75t_SL g3085 ( 
.A1(n_3065),
.A2(n_493),
.B(n_490),
.C(n_492),
.Y(n_3085)
);

XOR2xp5_ASAP7_75t_L g3086 ( 
.A(n_3050),
.B(n_493),
.Y(n_3086)
);

OAI211xp5_ASAP7_75t_L g3087 ( 
.A1(n_3037),
.A2(n_496),
.B(n_494),
.C(n_495),
.Y(n_3087)
);

AOI22xp5_ASAP7_75t_L g3088 ( 
.A1(n_3029),
.A2(n_496),
.B1(n_494),
.B2(n_495),
.Y(n_3088)
);

A2O1A1Ixp33_ASAP7_75t_L g3089 ( 
.A1(n_3038),
.A2(n_3058),
.B(n_3056),
.C(n_3066),
.Y(n_3089)
);

NOR4xp75_ASAP7_75t_L g3090 ( 
.A(n_3041),
.B(n_499),
.C(n_497),
.D(n_498),
.Y(n_3090)
);

OAI211xp5_ASAP7_75t_SL g3091 ( 
.A1(n_3068),
.A2(n_500),
.B(n_498),
.C(n_499),
.Y(n_3091)
);

OAI22xp5_ASAP7_75t_L g3092 ( 
.A1(n_3069),
.A2(n_3049),
.B1(n_3059),
.B2(n_3035),
.Y(n_3092)
);

AOI221xp5_ASAP7_75t_L g3093 ( 
.A1(n_3028),
.A2(n_502),
.B1(n_500),
.B2(n_501),
.C(n_503),
.Y(n_3093)
);

AOI221xp5_ASAP7_75t_L g3094 ( 
.A1(n_3034),
.A2(n_505),
.B1(n_503),
.B2(n_504),
.C(n_506),
.Y(n_3094)
);

OAI22x1_ASAP7_75t_L g3095 ( 
.A1(n_3048),
.A2(n_509),
.B1(n_507),
.B2(n_508),
.Y(n_3095)
);

AOI221x1_ASAP7_75t_L g3096 ( 
.A1(n_3057),
.A2(n_510),
.B1(n_508),
.B2(n_509),
.C(n_511),
.Y(n_3096)
);

OAI22xp5_ASAP7_75t_L g3097 ( 
.A1(n_3062),
.A2(n_516),
.B1(n_514),
.B2(n_515),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_3047),
.B(n_517),
.Y(n_3098)
);

O2A1O1Ixp33_ASAP7_75t_L g3099 ( 
.A1(n_3071),
.A2(n_520),
.B(n_518),
.C(n_519),
.Y(n_3099)
);

AND3x4_ASAP7_75t_L g3100 ( 
.A(n_3044),
.B(n_518),
.C(n_519),
.Y(n_3100)
);

AOI221xp5_ASAP7_75t_SL g3101 ( 
.A1(n_3053),
.A2(n_522),
.B1(n_520),
.B2(n_521),
.C(n_523),
.Y(n_3101)
);

NOR3x2_ASAP7_75t_L g3102 ( 
.A(n_3039),
.B(n_525),
.C(n_526),
.Y(n_3102)
);

AOI211xp5_ASAP7_75t_L g3103 ( 
.A1(n_3054),
.A2(n_528),
.B(n_526),
.C(n_527),
.Y(n_3103)
);

AOI322xp5_ASAP7_75t_L g3104 ( 
.A1(n_3051),
.A2(n_533),
.A3(n_532),
.B1(n_530),
.B2(n_528),
.C1(n_529),
.C2(n_531),
.Y(n_3104)
);

AOI21xp5_ASAP7_75t_L g3105 ( 
.A1(n_3061),
.A2(n_534),
.B(n_535),
.Y(n_3105)
);

AOI22xp5_ASAP7_75t_L g3106 ( 
.A1(n_3052),
.A2(n_538),
.B1(n_536),
.B2(n_537),
.Y(n_3106)
);

AOI211xp5_ASAP7_75t_SL g3107 ( 
.A1(n_3067),
.A2(n_541),
.B(n_539),
.C(n_540),
.Y(n_3107)
);

OAI22xp5_ASAP7_75t_L g3108 ( 
.A1(n_3055),
.A2(n_543),
.B1(n_541),
.B2(n_542),
.Y(n_3108)
);

NAND4xp25_ASAP7_75t_SL g3109 ( 
.A(n_3030),
.B(n_545),
.C(n_542),
.D(n_544),
.Y(n_3109)
);

OAI321xp33_ASAP7_75t_L g3110 ( 
.A1(n_3060),
.A2(n_547),
.A3(n_550),
.B1(n_544),
.B2(n_546),
.C(n_548),
.Y(n_3110)
);

OAI211xp5_ASAP7_75t_SL g3111 ( 
.A1(n_3060),
.A2(n_550),
.B(n_546),
.C(n_548),
.Y(n_3111)
);

OAI211xp5_ASAP7_75t_SL g3112 ( 
.A1(n_3060),
.A2(n_553),
.B(n_551),
.C(n_552),
.Y(n_3112)
);

AOI322xp5_ASAP7_75t_L g3113 ( 
.A1(n_3060),
.A2(n_559),
.A3(n_558),
.B1(n_556),
.B2(n_554),
.C1(n_555),
.C2(n_557),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_3042),
.Y(n_3114)
);

XOR2x2_ASAP7_75t_L g3115 ( 
.A(n_3027),
.B(n_554),
.Y(n_3115)
);

OAI22xp5_ASAP7_75t_L g3116 ( 
.A1(n_3060),
.A2(n_557),
.B1(n_555),
.B2(n_556),
.Y(n_3116)
);

XNOR2xp5_ASAP7_75t_L g3117 ( 
.A(n_3027),
.B(n_559),
.Y(n_3117)
);

OAI322xp33_ASAP7_75t_L g3118 ( 
.A1(n_3063),
.A2(n_566),
.A3(n_564),
.B1(n_562),
.B2(n_560),
.C1(n_561),
.C2(n_563),
.Y(n_3118)
);

HB1xp67_ASAP7_75t_L g3119 ( 
.A(n_3090),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_3086),
.Y(n_3120)
);

NAND4xp75_ASAP7_75t_L g3121 ( 
.A(n_3114),
.B(n_563),
.C(n_560),
.D(n_561),
.Y(n_3121)
);

OA22x2_ASAP7_75t_L g3122 ( 
.A1(n_3106),
.A2(n_567),
.B1(n_564),
.B2(n_566),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_3095),
.Y(n_3123)
);

AO22x2_ASAP7_75t_L g3124 ( 
.A1(n_3092),
.A2(n_3082),
.B1(n_3077),
.B2(n_3078),
.Y(n_3124)
);

AOI21xp5_ASAP7_75t_L g3125 ( 
.A1(n_3089),
.A2(n_567),
.B(n_568),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_3100),
.Y(n_3126)
);

BUFx3_ASAP7_75t_L g3127 ( 
.A(n_3080),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_3102),
.Y(n_3128)
);

NOR2x1p5_ASAP7_75t_L g3129 ( 
.A(n_3098),
.B(n_568),
.Y(n_3129)
);

AND2x4_ASAP7_75t_L g3130 ( 
.A(n_3076),
.B(n_569),
.Y(n_3130)
);

OR2x2_ASAP7_75t_L g3131 ( 
.A(n_3081),
.B(n_569),
.Y(n_3131)
);

OAI21xp33_ASAP7_75t_L g3132 ( 
.A1(n_3117),
.A2(n_570),
.B(n_571),
.Y(n_3132)
);

OAI22xp5_ASAP7_75t_SL g3133 ( 
.A1(n_3075),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_3115),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_3118),
.Y(n_3135)
);

NOR2x1_ASAP7_75t_L g3136 ( 
.A(n_3109),
.B(n_572),
.Y(n_3136)
);

XNOR2x1_ASAP7_75t_L g3137 ( 
.A(n_3088),
.B(n_3108),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_3079),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_3101),
.B(n_573),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_3087),
.Y(n_3140)
);

NOR2xp33_ASAP7_75t_L g3141 ( 
.A(n_3111),
.B(n_573),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_3116),
.Y(n_3142)
);

OAI21xp33_ASAP7_75t_L g3143 ( 
.A1(n_3084),
.A2(n_3091),
.B(n_3085),
.Y(n_3143)
);

INVx4_ASAP7_75t_L g3144 ( 
.A(n_3103),
.Y(n_3144)
);

AOI31xp33_ASAP7_75t_L g3145 ( 
.A1(n_3107),
.A2(n_577),
.A3(n_574),
.B(n_575),
.Y(n_3145)
);

NAND4xp75_ASAP7_75t_L g3146 ( 
.A(n_3096),
.B(n_579),
.C(n_577),
.D(n_578),
.Y(n_3146)
);

NOR3xp33_ASAP7_75t_L g3147 ( 
.A(n_3112),
.B(n_578),
.C(n_579),
.Y(n_3147)
);

AND2x2_ASAP7_75t_L g3148 ( 
.A(n_3074),
.B(n_580),
.Y(n_3148)
);

INVx2_ASAP7_75t_L g3149 ( 
.A(n_3097),
.Y(n_3149)
);

OAI21xp5_ASAP7_75t_L g3150 ( 
.A1(n_3099),
.A2(n_580),
.B(n_581),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_3083),
.Y(n_3151)
);

OAI22x1_ASAP7_75t_L g3152 ( 
.A1(n_3073),
.A2(n_583),
.B1(n_581),
.B2(n_582),
.Y(n_3152)
);

AO211x2_ASAP7_75t_L g3153 ( 
.A1(n_3105),
.A2(n_585),
.B(n_583),
.C(n_584),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_3110),
.Y(n_3154)
);

HB1xp67_ASAP7_75t_L g3155 ( 
.A(n_3094),
.Y(n_3155)
);

HB1xp67_ASAP7_75t_L g3156 ( 
.A(n_3093),
.Y(n_3156)
);

AND2x4_ASAP7_75t_L g3157 ( 
.A(n_3127),
.B(n_3123),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_3133),
.Y(n_3158)
);

HB1xp67_ASAP7_75t_L g3159 ( 
.A(n_3146),
.Y(n_3159)
);

OR3x2_ASAP7_75t_L g3160 ( 
.A(n_3131),
.B(n_3113),
.C(n_3104),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_3122),
.Y(n_3161)
);

INVx2_ASAP7_75t_L g3162 ( 
.A(n_3121),
.Y(n_3162)
);

NAND4xp75_ASAP7_75t_L g3163 ( 
.A(n_3125),
.B(n_586),
.C(n_584),
.D(n_585),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_L g3164 ( 
.A(n_3130),
.B(n_586),
.Y(n_3164)
);

XOR2xp5_ASAP7_75t_L g3165 ( 
.A(n_3119),
.B(n_587),
.Y(n_3165)
);

XNOR2xp5_ASAP7_75t_L g3166 ( 
.A(n_3153),
.B(n_587),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_3129),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_3145),
.B(n_588),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_3139),
.Y(n_3169)
);

INVx4_ASAP7_75t_L g3170 ( 
.A(n_3124),
.Y(n_3170)
);

NAND2xp33_ASAP7_75t_L g3171 ( 
.A(n_3147),
.B(n_589),
.Y(n_3171)
);

OR2x2_ASAP7_75t_L g3172 ( 
.A(n_3126),
.B(n_590),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_3152),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_3124),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_3136),
.Y(n_3175)
);

AND2x2_ASAP7_75t_SL g3176 ( 
.A(n_3128),
.B(n_590),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_3148),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_3135),
.B(n_3141),
.Y(n_3178)
);

XNOR2xp5_ASAP7_75t_L g3179 ( 
.A(n_3137),
.B(n_591),
.Y(n_3179)
);

NOR2x1_ASAP7_75t_L g3180 ( 
.A(n_3140),
.B(n_593),
.Y(n_3180)
);

XNOR2xp5_ASAP7_75t_L g3181 ( 
.A(n_3120),
.B(n_593),
.Y(n_3181)
);

XNOR2xp5_ASAP7_75t_L g3182 ( 
.A(n_3134),
.B(n_3154),
.Y(n_3182)
);

HB1xp67_ASAP7_75t_L g3183 ( 
.A(n_3150),
.Y(n_3183)
);

OAI22xp5_ASAP7_75t_L g3184 ( 
.A1(n_3151),
.A2(n_596),
.B1(n_594),
.B2(n_595),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_3132),
.B(n_3143),
.Y(n_3185)
);

AOI21x1_ASAP7_75t_L g3186 ( 
.A1(n_3180),
.A2(n_3142),
.B(n_3138),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_3165),
.Y(n_3187)
);

HB1xp67_ASAP7_75t_L g3188 ( 
.A(n_3166),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_3179),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_3181),
.Y(n_3190)
);

AOI21xp5_ASAP7_75t_L g3191 ( 
.A1(n_3171),
.A2(n_3155),
.B(n_3156),
.Y(n_3191)
);

INVx2_ASAP7_75t_SL g3192 ( 
.A(n_3176),
.Y(n_3192)
);

OAI22xp5_ASAP7_75t_SL g3193 ( 
.A1(n_3170),
.A2(n_3175),
.B1(n_3168),
.B2(n_3158),
.Y(n_3193)
);

AOI21x1_ASAP7_75t_L g3194 ( 
.A1(n_3159),
.A2(n_3149),
.B(n_3144),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_3172),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_3164),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_3163),
.Y(n_3197)
);

XNOR2xp5_ASAP7_75t_L g3198 ( 
.A(n_3182),
.B(n_594),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_3157),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_3198),
.Y(n_3200)
);

NOR3xp33_ASAP7_75t_L g3201 ( 
.A(n_3193),
.B(n_3174),
.C(n_3185),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_3186),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_3199),
.Y(n_3203)
);

OAI21xp5_ASAP7_75t_L g3204 ( 
.A1(n_3191),
.A2(n_3161),
.B(n_3178),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3188),
.Y(n_3205)
);

OAI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_3197),
.A2(n_3160),
.B1(n_3162),
.B2(n_3173),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_3194),
.Y(n_3207)
);

BUFx2_ASAP7_75t_L g3208 ( 
.A(n_3192),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_3187),
.Y(n_3209)
);

OAI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_3189),
.A2(n_3183),
.B(n_3167),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_3203),
.Y(n_3211)
);

AND2x4_ASAP7_75t_L g3212 ( 
.A(n_3201),
.B(n_3204),
.Y(n_3212)
);

AND2x2_ASAP7_75t_L g3213 ( 
.A(n_3208),
.B(n_3195),
.Y(n_3213)
);

OAI21xp5_ASAP7_75t_L g3214 ( 
.A1(n_3206),
.A2(n_3190),
.B(n_3169),
.Y(n_3214)
);

OAI22xp5_ASAP7_75t_SL g3215 ( 
.A1(n_3207),
.A2(n_3177),
.B1(n_3196),
.B2(n_3184),
.Y(n_3215)
);

OAI22xp5_ASAP7_75t_SL g3216 ( 
.A1(n_3202),
.A2(n_598),
.B1(n_595),
.B2(n_597),
.Y(n_3216)
);

OAI22xp5_ASAP7_75t_L g3217 ( 
.A1(n_3205),
.A2(n_599),
.B1(n_597),
.B2(n_598),
.Y(n_3217)
);

OAI22x1_ASAP7_75t_SL g3218 ( 
.A1(n_3200),
.A2(n_601),
.B1(n_599),
.B2(n_600),
.Y(n_3218)
);

OAI22x1_ASAP7_75t_L g3219 ( 
.A1(n_3209),
.A2(n_605),
.B1(n_602),
.B2(n_604),
.Y(n_3219)
);

AOI22xp5_ASAP7_75t_SL g3220 ( 
.A1(n_3212),
.A2(n_3210),
.B1(n_607),
.B2(n_602),
.Y(n_3220)
);

OAI21xp5_ASAP7_75t_L g3221 ( 
.A1(n_3213),
.A2(n_606),
.B(n_607),
.Y(n_3221)
);

OAI22xp5_ASAP7_75t_L g3222 ( 
.A1(n_3211),
.A2(n_610),
.B1(n_608),
.B2(n_609),
.Y(n_3222)
);

OAI21x1_ASAP7_75t_L g3223 ( 
.A1(n_3214),
.A2(n_608),
.B(n_609),
.Y(n_3223)
);

OAI22xp5_ASAP7_75t_SL g3224 ( 
.A1(n_3215),
.A2(n_612),
.B1(n_610),
.B2(n_611),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_3219),
.Y(n_3225)
);

INVxp67_ASAP7_75t_SL g3226 ( 
.A(n_3218),
.Y(n_3226)
);

AOI22xp5_ASAP7_75t_L g3227 ( 
.A1(n_3216),
.A2(n_615),
.B1(n_613),
.B2(n_614),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3217),
.Y(n_3228)
);

AND2x2_ASAP7_75t_L g3229 ( 
.A(n_3226),
.B(n_616),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_SL g3230 ( 
.A(n_3227),
.B(n_616),
.Y(n_3230)
);

NAND3xp33_ASAP7_75t_L g3231 ( 
.A(n_3220),
.B(n_619),
.C(n_620),
.Y(n_3231)
);

OA21x2_ASAP7_75t_L g3232 ( 
.A1(n_3225),
.A2(n_3228),
.B(n_3223),
.Y(n_3232)
);

OAI22xp5_ASAP7_75t_L g3233 ( 
.A1(n_3224),
.A2(n_623),
.B1(n_621),
.B2(n_622),
.Y(n_3233)
);

INVxp67_ASAP7_75t_L g3234 ( 
.A(n_3229),
.Y(n_3234)
);

XNOR2xp5_ASAP7_75t_L g3235 ( 
.A(n_3231),
.B(n_3221),
.Y(n_3235)
);

AOI222xp33_ASAP7_75t_L g3236 ( 
.A1(n_3230),
.A2(n_3222),
.B1(n_624),
.B2(n_626),
.C1(n_622),
.C2(n_623),
.Y(n_3236)
);

OAI22xp5_ASAP7_75t_SL g3237 ( 
.A1(n_3232),
.A2(n_626),
.B1(n_624),
.B2(n_625),
.Y(n_3237)
);

AO22x2_ASAP7_75t_L g3238 ( 
.A1(n_3233),
.A2(n_629),
.B1(n_625),
.B2(n_627),
.Y(n_3238)
);

OAI221xp5_ASAP7_75t_R g3239 ( 
.A1(n_3235),
.A2(n_3234),
.B1(n_3236),
.B2(n_3238),
.C(n_3237),
.Y(n_3239)
);

AOI22xp5_ASAP7_75t_SL g3240 ( 
.A1(n_3235),
.A2(n_632),
.B1(n_630),
.B2(n_631),
.Y(n_3240)
);

AO21x2_ASAP7_75t_L g3241 ( 
.A1(n_3239),
.A2(n_3240),
.B(n_633),
.Y(n_3241)
);

AOI221xp5_ASAP7_75t_L g3242 ( 
.A1(n_3241),
.A2(n_639),
.B1(n_635),
.B2(n_638),
.C(n_640),
.Y(n_3242)
);

AOI211xp5_ASAP7_75t_L g3243 ( 
.A1(n_3242),
.A2(n_641),
.B(n_638),
.C(n_639),
.Y(n_3243)
);


endmodule