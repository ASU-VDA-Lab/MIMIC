module real_aes_8028_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_717;
wire n_359;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g108 ( .A(n_0), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_1), .A2(n_152), .B(n_157), .C(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g264 ( .A(n_2), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_3), .A2(n_147), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_4), .B(n_224), .Y(n_473) );
AOI21xp33_ASAP7_75t_L g225 ( .A1(n_5), .A2(n_147), .B(n_226), .Y(n_225) );
AND2x6_ASAP7_75t_L g152 ( .A(n_6), .B(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_7), .A2(n_146), .B(n_154), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_8), .B(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_8), .B(n_40), .Y(n_125) );
INVx1_ASAP7_75t_L g562 ( .A(n_9), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_10), .B(n_196), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_11), .B(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g231 ( .A(n_12), .Y(n_231) );
INVx1_ASAP7_75t_L g144 ( .A(n_13), .Y(n_144) );
INVx1_ASAP7_75t_L g164 ( .A(n_14), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_15), .A2(n_165), .B(n_179), .C(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_16), .B(n_224), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_17), .B(n_181), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_18), .B(n_147), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_19), .B(n_486), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_20), .A2(n_212), .B(n_238), .C(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_21), .B(n_224), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_22), .B(n_196), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g160 ( .A1(n_23), .A2(n_161), .B(n_163), .C(n_165), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_24), .B(n_196), .Y(n_459) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_25), .Y(n_490) );
INVx1_ASAP7_75t_L g458 ( .A(n_26), .Y(n_458) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_27), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_28), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_29), .B(n_196), .Y(n_265) );
INVx1_ASAP7_75t_L g483 ( .A(n_30), .Y(n_483) );
INVx1_ASAP7_75t_L g243 ( .A(n_31), .Y(n_243) );
INVx2_ASAP7_75t_L g150 ( .A(n_32), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_33), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_34), .A2(n_212), .B(n_232), .C(n_471), .Y(n_470) );
INVxp67_ASAP7_75t_L g484 ( .A(n_35), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_36), .A2(n_152), .B(n_157), .C(n_176), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_37), .A2(n_157), .B(n_457), .C(n_462), .Y(n_456) );
CKINVDCx14_ASAP7_75t_R g469 ( .A(n_38), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_39), .A2(n_67), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_39), .Y(n_129) );
INVx1_ASAP7_75t_L g114 ( .A(n_40), .Y(n_114) );
INVx1_ASAP7_75t_L g241 ( .A(n_41), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_42), .A2(n_183), .B(n_229), .C(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_43), .B(n_196), .Y(n_195) );
OAI22xp5_ASAP7_75t_SL g721 ( .A1(n_44), .A2(n_83), .B1(n_722), .B2(n_723), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_44), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_45), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_46), .Y(n_480) );
INVx1_ASAP7_75t_L g528 ( .A(n_47), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g244 ( .A(n_48), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_49), .B(n_147), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_50), .A2(n_157), .B1(n_238), .B2(n_240), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_51), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g261 ( .A(n_52), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_53), .A2(n_229), .B(n_230), .C(n_232), .Y(n_228) );
CKINVDCx14_ASAP7_75t_R g559 ( .A(n_54), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_55), .Y(n_200) );
INVx1_ASAP7_75t_L g227 ( .A(n_56), .Y(n_227) );
AOI222xp33_ASAP7_75t_SL g127 ( .A1(n_57), .A2(n_128), .B1(n_131), .B2(n_712), .C1(n_713), .C2(n_714), .Y(n_127) );
INVx1_ASAP7_75t_L g153 ( .A(n_58), .Y(n_153) );
INVx1_ASAP7_75t_L g143 ( .A(n_59), .Y(n_143) );
INVx1_ASAP7_75t_SL g472 ( .A(n_60), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_61), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_62), .B(n_224), .Y(n_532) );
INVx1_ASAP7_75t_L g493 ( .A(n_63), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_SL g251 ( .A1(n_64), .A2(n_181), .B(n_232), .C(n_252), .Y(n_251) );
INVxp67_ASAP7_75t_L g253 ( .A(n_65), .Y(n_253) );
INVx1_ASAP7_75t_L g111 ( .A(n_66), .Y(n_111) );
INVx1_ASAP7_75t_L g130 ( .A(n_67), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_68), .A2(n_147), .B(n_558), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_69), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_70), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_71), .A2(n_147), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g191 ( .A(n_72), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_73), .A2(n_146), .B(n_479), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g455 ( .A(n_74), .Y(n_455) );
INVx1_ASAP7_75t_L g520 ( .A(n_75), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_76), .A2(n_152), .B(n_157), .C(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_77), .A2(n_147), .B(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g523 ( .A(n_78), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_79), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g141 ( .A(n_80), .Y(n_141) );
INVx1_ASAP7_75t_L g512 ( .A(n_81), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_82), .B(n_181), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_83), .Y(n_722) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_84), .A2(n_152), .B(n_157), .C(n_263), .Y(n_262) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_85), .B(n_108), .C(n_109), .Y(n_107) );
OR2x2_ASAP7_75t_L g122 ( .A(n_85), .B(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g444 ( .A(n_85), .Y(n_444) );
OR2x2_ASAP7_75t_L g711 ( .A(n_85), .B(n_124), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_86), .A2(n_157), .B(n_492), .C(n_496), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_87), .B(n_140), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_88), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_89), .A2(n_152), .B(n_157), .C(n_209), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g217 ( .A(n_90), .Y(n_217) );
INVx1_ASAP7_75t_L g250 ( .A(n_91), .Y(n_250) );
CKINVDCx16_ASAP7_75t_R g155 ( .A(n_92), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_93), .B(n_178), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_94), .B(n_169), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_95), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_96), .B(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_97), .A2(n_147), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g531 ( .A(n_98), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_99), .A2(n_102), .B1(n_115), .B2(n_725), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_100), .Y(n_126) );
BUFx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_SL g727 ( .A(n_105), .Y(n_727) );
AND2x2_ASAP7_75t_SL g105 ( .A(n_106), .B(n_112), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g124 ( .A(n_108), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AOI22x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_127), .B1(n_717), .B2(n_719), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_120), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g718 ( .A(n_119), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_120), .A2(n_720), .B(n_724), .Y(n_719) );
NOR2xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_126), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_122), .Y(n_724) );
NOR2x2_ASAP7_75t_L g716 ( .A(n_123), .B(n_444), .Y(n_716) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g443 ( .A(n_124), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g712 ( .A(n_128), .Y(n_712) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_441), .B1(n_445), .B2(n_709), .Y(n_131) );
INVx2_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g713 ( .A1(n_133), .A2(n_443), .B1(n_446), .B2(n_711), .Y(n_713) );
OR4x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_337), .C(n_396), .D(n_423), .Y(n_133) );
NAND3xp33_ASAP7_75t_SL g134 ( .A(n_135), .B(n_279), .C(n_304), .Y(n_134) );
O2A1O1Ixp33_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_202), .B(n_222), .C(n_255), .Y(n_135) );
AOI211xp5_ASAP7_75t_SL g427 ( .A1(n_136), .A2(n_428), .B(n_430), .C(n_433), .Y(n_427) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_171), .Y(n_136) );
INVx1_ASAP7_75t_L g302 ( .A(n_137), .Y(n_302) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g277 ( .A(n_138), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g309 ( .A(n_138), .Y(n_309) );
AND2x2_ASAP7_75t_L g364 ( .A(n_138), .B(n_333), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_138), .B(n_220), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_138), .B(n_221), .Y(n_422) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g283 ( .A(n_139), .Y(n_283) );
AND2x2_ASAP7_75t_L g326 ( .A(n_139), .B(n_189), .Y(n_326) );
AND2x2_ASAP7_75t_L g344 ( .A(n_139), .B(n_221), .Y(n_344) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_145), .B(n_168), .Y(n_139) );
INVx1_ASAP7_75t_L g201 ( .A(n_140), .Y(n_201) );
INVx2_ASAP7_75t_L g206 ( .A(n_140), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g454 ( .A1(n_140), .A2(n_192), .B(n_455), .C(n_456), .Y(n_454) );
OA21x2_ASAP7_75t_L g556 ( .A1(n_140), .A2(n_557), .B(n_563), .Y(n_556) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_L g170 ( .A(n_141), .B(n_142), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
NAND2x1p5_ASAP7_75t_L g192 ( .A(n_148), .B(n_152), .Y(n_192) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx1_ASAP7_75t_L g461 ( .A(n_149), .Y(n_461) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
INVx1_ASAP7_75t_L g239 ( .A(n_150), .Y(n_239) );
INVx1_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_151), .Y(n_162) );
INVx3_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
INVx1_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
INVx4_ASAP7_75t_SL g167 ( .A(n_152), .Y(n_167) );
BUFx3_ASAP7_75t_L g462 ( .A(n_152), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_160), .C(n_167), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_156), .A2(n_167), .B(n_227), .C(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_156), .A2(n_167), .B(n_250), .C(n_251), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_156), .A2(n_167), .B(n_469), .C(n_470), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_SL g479 ( .A1(n_156), .A2(n_167), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g519 ( .A1(n_156), .A2(n_167), .B(n_520), .C(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_SL g527 ( .A1(n_156), .A2(n_167), .B(n_528), .C(n_529), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_SL g558 ( .A1(n_156), .A2(n_167), .B(n_559), .C(n_560), .Y(n_558) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x6_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
BUFx3_ASAP7_75t_L g166 ( .A(n_158), .Y(n_166) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_158), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_161), .B(n_164), .Y(n_163) );
OAI22xp33_ASAP7_75t_L g482 ( .A1(n_161), .A2(n_178), .B1(n_483), .B2(n_484), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_161), .B(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_161), .B(n_531), .Y(n_530) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_SL g240 ( .A1(n_162), .A2(n_241), .B1(n_242), .B2(n_243), .Y(n_240) );
INVx2_ASAP7_75t_L g242 ( .A(n_162), .Y(n_242) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g183 ( .A(n_166), .Y(n_183) );
OAI22xp33_ASAP7_75t_L g236 ( .A1(n_167), .A2(n_192), .B1(n_237), .B2(n_244), .Y(n_236) );
INVx1_ASAP7_75t_L g496 ( .A(n_167), .Y(n_496) );
INVx4_ASAP7_75t_L g188 ( .A(n_169), .Y(n_188) );
OA21x2_ASAP7_75t_L g247 ( .A1(n_169), .A2(n_248), .B(n_254), .Y(n_247) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_169), .Y(n_466) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g185 ( .A(n_170), .Y(n_185) );
INVx4_ASAP7_75t_L g276 ( .A(n_171), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g331 ( .A1(n_171), .A2(n_332), .B(n_334), .Y(n_331) );
AND2x2_ASAP7_75t_L g412 ( .A(n_171), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_189), .Y(n_171) );
INVx1_ASAP7_75t_L g219 ( .A(n_172), .Y(n_219) );
AND2x2_ASAP7_75t_L g281 ( .A(n_172), .B(n_221), .Y(n_281) );
OR2x2_ASAP7_75t_L g310 ( .A(n_172), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g324 ( .A(n_172), .Y(n_324) );
INVx3_ASAP7_75t_L g333 ( .A(n_172), .Y(n_333) );
AND2x2_ASAP7_75t_L g343 ( .A(n_172), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g376 ( .A(n_172), .B(n_282), .Y(n_376) );
AND2x2_ASAP7_75t_L g400 ( .A(n_172), .B(n_356), .Y(n_400) );
OR2x6_ASAP7_75t_L g172 ( .A(n_173), .B(n_186), .Y(n_172) );
AOI21xp5_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_175), .B(n_184), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_180), .B(n_182), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_178), .A2(n_264), .B(n_265), .C(n_266), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_178), .A2(n_458), .B(n_459), .C(n_460), .Y(n_457) );
INVx5_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_179), .B(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_179), .B(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_179), .B(n_562), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_182), .A2(n_195), .B(n_197), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_182), .A2(n_493), .B(n_494), .C(n_495), .Y(n_492) );
O2A1O1Ixp5_ASAP7_75t_L g511 ( .A1(n_182), .A2(n_494), .B(n_512), .C(n_513), .Y(n_511) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g198 ( .A(n_184), .Y(n_198) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_185), .A2(n_236), .B(n_245), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_185), .B(n_246), .Y(n_245) );
AO21x2_ASAP7_75t_L g259 ( .A1(n_185), .A2(n_260), .B(n_267), .Y(n_259) );
NOR2xp33_ASAP7_75t_SL g186 ( .A(n_187), .B(n_188), .Y(n_186) );
INVx3_ASAP7_75t_L g224 ( .A(n_188), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_188), .B(n_464), .Y(n_463) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_188), .A2(n_489), .B(n_497), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_188), .B(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g221 ( .A(n_189), .Y(n_221) );
AND2x2_ASAP7_75t_L g436 ( .A(n_189), .B(n_278), .Y(n_436) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_198), .B(n_199), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_193), .Y(n_190) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_192), .A2(n_261), .B(n_262), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g489 ( .A1(n_192), .A2(n_490), .B(n_491), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_192), .A2(n_509), .B(n_510), .Y(n_508) );
INVx4_ASAP7_75t_L g212 ( .A(n_196), .Y(n_212) );
INVx2_ASAP7_75t_L g229 ( .A(n_196), .Y(n_229) );
INVx1_ASAP7_75t_L g477 ( .A(n_198), .Y(n_477) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_198), .A2(n_502), .B(n_503), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_201), .B(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_201), .B(n_268), .Y(n_267) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_201), .A2(n_508), .B(n_514), .Y(n_507) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_218), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_204), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g356 ( .A(n_204), .B(n_344), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_204), .B(n_333), .Y(n_418) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g278 ( .A(n_205), .Y(n_278) );
AND2x2_ASAP7_75t_L g282 ( .A(n_205), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g323 ( .A(n_205), .B(n_324), .Y(n_323) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_216), .Y(n_205) );
INVx1_ASAP7_75t_L g486 ( .A(n_206), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_206), .B(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_215), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_213), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_212), .B(n_472), .Y(n_471) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx3_ASAP7_75t_L g232 ( .A(n_214), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_218), .B(n_319), .Y(n_341) );
INVx1_ASAP7_75t_L g380 ( .A(n_218), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_218), .B(n_307), .Y(n_424) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
AND2x2_ASAP7_75t_L g287 ( .A(n_219), .B(n_282), .Y(n_287) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_221), .B(n_278), .Y(n_311) );
INVx1_ASAP7_75t_L g390 ( .A(n_221), .Y(n_390) );
AOI322xp5_ASAP7_75t_L g414 ( .A1(n_222), .A2(n_329), .A3(n_389), .B1(n_415), .B2(n_417), .C1(n_419), .C2(n_421), .Y(n_414) );
AND2x2_ASAP7_75t_SL g222 ( .A(n_223), .B(n_234), .Y(n_222) );
AND2x2_ASAP7_75t_L g269 ( .A(n_223), .B(n_247), .Y(n_269) );
INVx1_ASAP7_75t_SL g272 ( .A(n_223), .Y(n_272) );
AND2x2_ASAP7_75t_L g274 ( .A(n_223), .B(n_235), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_223), .B(n_291), .Y(n_297) );
INVx2_ASAP7_75t_L g316 ( .A(n_223), .Y(n_316) );
AND2x2_ASAP7_75t_L g329 ( .A(n_223), .B(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g367 ( .A(n_223), .B(n_291), .Y(n_367) );
BUFx2_ASAP7_75t_L g384 ( .A(n_223), .Y(n_384) );
AND2x2_ASAP7_75t_L g398 ( .A(n_223), .B(n_258), .Y(n_398) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_233), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_234), .B(n_286), .Y(n_313) );
AND2x2_ASAP7_75t_L g440 ( .A(n_234), .B(n_316), .Y(n_440) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_247), .Y(n_234) );
OR2x2_ASAP7_75t_L g285 ( .A(n_235), .B(n_286), .Y(n_285) );
INVx3_ASAP7_75t_L g291 ( .A(n_235), .Y(n_291) );
AND2x2_ASAP7_75t_L g336 ( .A(n_235), .B(n_259), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_235), .B(n_384), .Y(n_383) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_235), .Y(n_420) );
INVx2_ASAP7_75t_L g266 ( .A(n_238), .Y(n_266) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g494 ( .A(n_242), .Y(n_494) );
AND2x2_ASAP7_75t_L g271 ( .A(n_247), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g293 ( .A(n_247), .Y(n_293) );
BUFx2_ASAP7_75t_L g299 ( .A(n_247), .Y(n_299) );
AND2x2_ASAP7_75t_L g318 ( .A(n_247), .B(n_291), .Y(n_318) );
INVx3_ASAP7_75t_L g330 ( .A(n_247), .Y(n_330) );
OR2x2_ASAP7_75t_L g340 ( .A(n_247), .B(n_291), .Y(n_340) );
AOI31xp33_ASAP7_75t_SL g255 ( .A1(n_256), .A2(n_270), .A3(n_273), .B(n_275), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_269), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_257), .B(n_292), .Y(n_303) );
OR2x2_ASAP7_75t_L g327 ( .A(n_257), .B(n_297), .Y(n_327) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_258), .B(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g348 ( .A(n_258), .B(n_340), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_258), .B(n_330), .Y(n_358) );
AND2x2_ASAP7_75t_L g365 ( .A(n_258), .B(n_366), .Y(n_365) );
NAND2x1_ASAP7_75t_L g393 ( .A(n_258), .B(n_329), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_258), .B(n_384), .Y(n_394) );
AND2x2_ASAP7_75t_L g406 ( .A(n_258), .B(n_291), .Y(n_406) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g286 ( .A(n_259), .Y(n_286) );
INVx1_ASAP7_75t_L g352 ( .A(n_269), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_269), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_271), .B(n_347), .Y(n_381) );
AND2x4_ASAP7_75t_L g292 ( .A(n_272), .B(n_293), .Y(n_292) );
CKINVDCx16_ASAP7_75t_R g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx2_ASAP7_75t_L g371 ( .A(n_277), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_277), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g319 ( .A(n_278), .B(n_309), .Y(n_319) );
AND2x2_ASAP7_75t_L g413 ( .A(n_278), .B(n_283), .Y(n_413) );
INVx1_ASAP7_75t_L g438 ( .A(n_278), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_284), .B1(n_287), .B2(n_288), .C(n_294), .Y(n_279) );
CKINVDCx14_ASAP7_75t_R g300 ( .A(n_280), .Y(n_300) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_281), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_284), .B(n_335), .Y(n_354) );
INVx3_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g403 ( .A(n_285), .B(n_299), .Y(n_403) );
AND2x2_ASAP7_75t_L g317 ( .A(n_286), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g347 ( .A(n_286), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_286), .B(n_330), .Y(n_375) );
NOR3xp33_ASAP7_75t_L g417 ( .A(n_286), .B(n_387), .C(n_418), .Y(n_417) );
AOI211xp5_ASAP7_75t_SL g350 ( .A1(n_287), .A2(n_351), .B(n_353), .C(n_361), .Y(n_350) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OAI22xp33_ASAP7_75t_L g339 ( .A1(n_289), .A2(n_340), .B1(n_341), .B2(n_342), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_290), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_290), .B(n_374), .Y(n_373) );
BUFx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g432 ( .A(n_292), .B(n_406), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_300), .B1(n_301), .B2(n_303), .Y(n_294) );
NOR2xp33_ASAP7_75t_SL g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_298), .B(n_347), .Y(n_378) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_301), .A2(n_393), .B1(n_424), .B2(n_431), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_312), .B1(n_314), .B2(n_319), .C(n_320), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_310), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OAI221xp5_ASAP7_75t_L g320 ( .A1(n_310), .A2(n_321), .B1(n_327), .B2(n_328), .C(n_331), .Y(n_320) );
INVx1_ASAP7_75t_L g363 ( .A(n_311), .Y(n_363) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_SL g335 ( .A(n_316), .Y(n_335) );
OR2x2_ASAP7_75t_L g408 ( .A(n_316), .B(n_340), .Y(n_408) );
AND2x2_ASAP7_75t_L g410 ( .A(n_316), .B(n_318), .Y(n_410) );
INVx1_ASAP7_75t_L g349 ( .A(n_319), .Y(n_349) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_325), .Y(n_321) );
AOI21xp33_ASAP7_75t_SL g379 ( .A1(n_322), .A2(n_380), .B(n_381), .Y(n_379) );
OR2x2_ASAP7_75t_L g386 ( .A(n_322), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g360 ( .A(n_323), .B(n_344), .Y(n_360) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp33_ASAP7_75t_SL g377 ( .A(n_328), .B(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_329), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_330), .B(n_366), .Y(n_429) );
O2A1O1Ixp33_ASAP7_75t_L g345 ( .A1(n_333), .A2(n_346), .B(n_348), .C(n_349), .Y(n_345) );
NAND2x1_ASAP7_75t_SL g370 ( .A(n_333), .B(n_371), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_334), .A2(n_383), .B1(n_385), .B2(n_388), .Y(n_382) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_336), .B(n_426), .Y(n_425) );
NAND5xp2_ASAP7_75t_L g337 ( .A(n_338), .B(n_350), .C(n_368), .D(n_382), .E(n_391), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_345), .Y(n_338) );
INVx1_ASAP7_75t_L g395 ( .A(n_341), .Y(n_395) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_343), .A2(n_362), .B1(n_402), .B2(n_404), .C(n_407), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_344), .B(n_438), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_347), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_347), .B(n_413), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_357), .B2(n_359), .Y(n_353) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_365), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
AND2x2_ASAP7_75t_L g435 ( .A(n_364), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_372), .B1(n_376), .B2(n_377), .C(n_379), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g419 ( .A(n_374), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g426 ( .A(n_384), .Y(n_426) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OAI21xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_394), .B(n_395), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI211xp5_ASAP7_75t_SL g396 ( .A1(n_397), .A2(n_399), .B(n_401), .C(n_414), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
A2O1A1Ixp33_ASAP7_75t_L g423 ( .A1(n_399), .A2(n_424), .B(n_425), .C(n_427), .Y(n_423) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_403), .B(n_405), .Y(n_404) );
AOI21xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B(n_411), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI21xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_437), .B(n_439), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
XOR2xp5_ASAP7_75t_L g720 ( .A(n_446), .B(n_721), .Y(n_720) );
OR3x1_ASAP7_75t_L g446 ( .A(n_447), .B(n_620), .C(n_667), .Y(n_446) );
NAND3xp33_ASAP7_75t_SL g447 ( .A(n_448), .B(n_566), .C(n_591), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_506), .B1(n_533), .B2(n_536), .C(n_544), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_474), .B(n_499), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_451), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_451), .B(n_549), .Y(n_664) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_465), .Y(n_451) );
AND2x2_ASAP7_75t_L g535 ( .A(n_452), .B(n_505), .Y(n_535) );
AND2x2_ASAP7_75t_L g584 ( .A(n_452), .B(n_504), .Y(n_584) );
AND2x2_ASAP7_75t_L g605 ( .A(n_452), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g610 ( .A(n_452), .B(n_577), .Y(n_610) );
OR2x2_ASAP7_75t_L g618 ( .A(n_452), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g690 ( .A(n_452), .B(n_487), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_452), .B(n_639), .Y(n_704) );
INVx3_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g550 ( .A(n_453), .B(n_465), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_453), .B(n_487), .Y(n_551) );
AND2x4_ASAP7_75t_L g572 ( .A(n_453), .B(n_505), .Y(n_572) );
AND2x2_ASAP7_75t_L g602 ( .A(n_453), .B(n_476), .Y(n_602) );
AND2x2_ASAP7_75t_L g611 ( .A(n_453), .B(n_601), .Y(n_611) );
AND2x2_ASAP7_75t_L g627 ( .A(n_453), .B(n_488), .Y(n_627) );
OR2x2_ASAP7_75t_L g636 ( .A(n_453), .B(n_619), .Y(n_636) );
AND2x2_ASAP7_75t_L g642 ( .A(n_453), .B(n_577), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_453), .B(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g656 ( .A(n_453), .B(n_501), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_453), .B(n_546), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_453), .B(n_606), .Y(n_695) );
OR2x6_ASAP7_75t_L g453 ( .A(n_454), .B(n_463), .Y(n_453) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_461), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g505 ( .A(n_465), .Y(n_505) );
AND2x2_ASAP7_75t_L g601 ( .A(n_465), .B(n_487), .Y(n_601) );
AND2x2_ASAP7_75t_L g606 ( .A(n_465), .B(n_488), .Y(n_606) );
INVx1_ASAP7_75t_L g662 ( .A(n_465), .Y(n_662) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B(n_473), .Y(n_465) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_466), .A2(n_518), .B(n_524), .Y(n_517) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_466), .A2(n_526), .B(n_532), .Y(n_525) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g571 ( .A(n_475), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_487), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_476), .B(n_535), .Y(n_534) );
BUFx3_ASAP7_75t_L g549 ( .A(n_476), .Y(n_549) );
OR2x2_ASAP7_75t_L g619 ( .A(n_476), .B(n_487), .Y(n_619) );
OR2x2_ASAP7_75t_L g680 ( .A(n_476), .B(n_587), .Y(n_680) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_485), .Y(n_476) );
INVx1_ASAP7_75t_L g502 ( .A(n_478), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_485), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_487), .B(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g639 ( .A(n_487), .B(n_501), .Y(n_639) );
INVx2_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g578 ( .A(n_488), .Y(n_578) );
INVx1_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_500), .A2(n_684), .B1(n_688), .B2(n_691), .C(n_692), .Y(n_683) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_504), .Y(n_500) );
INVx1_ASAP7_75t_SL g547 ( .A(n_501), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_501), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g678 ( .A(n_501), .B(n_535), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_504), .B(n_549), .Y(n_670) );
AND2x2_ASAP7_75t_L g577 ( .A(n_505), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_SL g581 ( .A(n_506), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_506), .B(n_587), .Y(n_617) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_516), .Y(n_506) );
AND2x2_ASAP7_75t_L g543 ( .A(n_507), .B(n_517), .Y(n_543) );
INVx4_ASAP7_75t_L g555 ( .A(n_507), .Y(n_555) );
BUFx3_ASAP7_75t_L g597 ( .A(n_507), .Y(n_597) );
AND3x2_ASAP7_75t_L g612 ( .A(n_507), .B(n_613), .C(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g694 ( .A(n_516), .B(n_608), .Y(n_694) );
AND2x2_ASAP7_75t_L g702 ( .A(n_516), .B(n_587), .Y(n_702) );
INVx1_ASAP7_75t_SL g707 ( .A(n_516), .Y(n_707) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_525), .Y(n_516) );
INVx1_ASAP7_75t_SL g565 ( .A(n_517), .Y(n_565) );
AND2x2_ASAP7_75t_L g588 ( .A(n_517), .B(n_555), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_517), .B(n_539), .Y(n_590) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_517), .Y(n_630) );
OR2x2_ASAP7_75t_L g635 ( .A(n_517), .B(n_555), .Y(n_635) );
INVx2_ASAP7_75t_L g541 ( .A(n_525), .Y(n_541) );
AND2x2_ASAP7_75t_L g575 ( .A(n_525), .B(n_556), .Y(n_575) );
OR2x2_ASAP7_75t_L g595 ( .A(n_525), .B(n_556), .Y(n_595) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_525), .Y(n_615) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
AOI21xp33_ASAP7_75t_L g665 ( .A1(n_534), .A2(n_574), .B(n_666), .Y(n_665) );
AOI322xp5_ASAP7_75t_L g701 ( .A1(n_536), .A2(n_546), .A3(n_572), .B1(n_702), .B2(n_703), .C1(n_705), .C2(n_708), .Y(n_701) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_542), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_538), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_539), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g564 ( .A(n_540), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g632 ( .A(n_541), .B(n_555), .Y(n_632) );
AND2x2_ASAP7_75t_L g699 ( .A(n_541), .B(n_556), .Y(n_699) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g640 ( .A(n_543), .B(n_594), .Y(n_640) );
AOI31xp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_548), .A3(n_551), .B(n_552), .Y(n_544) );
AND2x2_ASAP7_75t_L g599 ( .A(n_546), .B(n_577), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_546), .B(n_569), .Y(n_681) );
AND2x2_ASAP7_75t_L g700 ( .A(n_546), .B(n_605), .Y(n_700) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_549), .B(n_577), .Y(n_589) );
NAND2x1p5_ASAP7_75t_L g623 ( .A(n_549), .B(n_606), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_549), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_549), .B(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_550), .B(n_606), .Y(n_638) );
INVx1_ASAP7_75t_L g682 ( .A(n_550), .Y(n_682) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_564), .Y(n_553) );
INVxp67_ASAP7_75t_L g634 ( .A(n_554), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_555), .B(n_565), .Y(n_570) );
INVx1_ASAP7_75t_L g676 ( .A(n_555), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_555), .B(n_653), .Y(n_687) );
BUFx3_ASAP7_75t_L g587 ( .A(n_556), .Y(n_587) );
AND2x2_ASAP7_75t_L g613 ( .A(n_556), .B(n_565), .Y(n_613) );
INVx2_ASAP7_75t_L g653 ( .A(n_556), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_564), .B(n_686), .Y(n_685) );
AOI211xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_571), .B(n_573), .C(n_582), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_568), .A2(n_617), .B(n_618), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_569), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_569), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g649 ( .A(n_570), .B(n_595), .Y(n_649) );
INVx3_ASAP7_75t_L g580 ( .A(n_572), .Y(n_580) );
OAI22xp5_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_576), .B1(n_579), .B2(n_581), .Y(n_573) );
OAI21xp5_ASAP7_75t_SL g598 ( .A1(n_575), .A2(n_599), .B(n_600), .Y(n_598) );
AND2x2_ASAP7_75t_L g624 ( .A(n_575), .B(n_588), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_575), .B(n_676), .Y(n_675) );
INVxp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g579 ( .A(n_578), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g648 ( .A(n_578), .Y(n_648) );
OAI21xp5_ASAP7_75t_SL g592 ( .A1(n_579), .A2(n_593), .B(n_598), .Y(n_592) );
OAI22xp33_ASAP7_75t_SL g582 ( .A1(n_583), .A2(n_585), .B1(n_589), .B2(n_590), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_584), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g608 ( .A(n_587), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_587), .B(n_630), .Y(n_629) );
NOR3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_603), .C(n_616), .Y(n_591) );
OAI22xp5_ASAP7_75t_SL g658 ( .A1(n_593), .A2(n_659), .B1(n_663), .B2(n_664), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_594), .B(n_596), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g663 ( .A(n_595), .B(n_596), .Y(n_663) );
AND2x2_ASAP7_75t_L g671 ( .A(n_596), .B(n_652), .Y(n_671) );
CKINVDCx16_ASAP7_75t_R g596 ( .A(n_597), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_SL g679 ( .A1(n_597), .A2(n_680), .B(n_681), .C(n_682), .Y(n_679) );
OR2x2_ASAP7_75t_L g706 ( .A(n_597), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_607), .B(n_609), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_L g641 ( .A1(n_605), .A2(n_642), .B(n_643), .C(n_646), .Y(n_641) );
OAI21xp33_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_611), .B(n_612), .Y(n_609) );
AND2x2_ASAP7_75t_L g674 ( .A(n_613), .B(n_632), .Y(n_674) );
INVxp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g652 ( .A(n_615), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g657 ( .A(n_617), .Y(n_657) );
NAND3xp33_ASAP7_75t_SL g620 ( .A(n_621), .B(n_641), .C(n_654), .Y(n_620) );
AOI211xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B(n_625), .C(n_633), .Y(n_621) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g691 ( .A(n_628), .Y(n_691) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g651 ( .A(n_630), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_630), .B(n_699), .Y(n_698) );
INVxp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_635), .B(n_636), .C(n_637), .Y(n_633) );
INVx2_ASAP7_75t_SL g645 ( .A(n_635), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_636), .A2(n_647), .B1(n_649), .B2(n_650), .Y(n_646) );
OAI21xp33_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_639), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
AOI211xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .B(n_658), .C(n_665), .Y(n_654) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVxp33_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g708 ( .A(n_662), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g667 ( .A(n_668), .B(n_683), .C(n_696), .D(n_701), .Y(n_667) );
AOI211xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B(n_672), .C(n_679), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .B(n_677), .Y(n_672) );
AOI21xp33_ASAP7_75t_L g692 ( .A1(n_673), .A2(n_693), .B(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_680), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_700), .Y(n_696) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
endmodule