module fake_jpeg_1735_n_144 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_56),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_69),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_39),
.B1(n_51),
.B2(n_42),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_42),
.B1(n_39),
.B2(n_52),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_42),
.B1(n_51),
.B2(n_50),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_50),
.B1(n_44),
.B2(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_40),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_74),
.Y(n_96)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_44),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_79),
.B1(n_83),
.B2(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_1),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_38),
.B1(n_2),
.B2(n_3),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_38),
.B(n_2),
.C(n_4),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_81),
.B(n_1),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_20),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_21),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_38),
.B1(n_4),
.B2(n_5),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

AO22x1_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_34),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_92),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_95),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_23),
.Y(n_104)
);

AO21x2_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_60),
.B(n_61),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_74),
.B1(n_81),
.B2(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_96),
.B(n_70),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_82),
.B(n_6),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_8),
.B(n_10),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_104),
.Y(n_116)
);

NAND2x1p5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_5),
.Y(n_106)
);

AOI21x1_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_113),
.B(n_7),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_6),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_108),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_26),
.B1(n_33),
.B2(n_31),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_7),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_86),
.C(n_97),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_122),
.C(n_125),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_124),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_30),
.C(n_29),
.Y(n_122)
);

AOI221xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_123),
.B(n_126),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_99),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_106),
.C(n_101),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_27),
.C(n_28),
.Y(n_126)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_11),
.Y(n_136)
);

HB1xp67_ASAP7_75t_SL g133 ( 
.A(n_130),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_133),
.A2(n_136),
.B(n_123),
.C(n_129),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_120),
.B1(n_117),
.B2(n_121),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_135),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_125),
.C(n_117),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_129),
.C(n_132),
.Y(n_139)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_135),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_141),
.A2(n_137),
.B(n_13),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_12),
.B(n_14),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_14),
.Y(n_144)
);


endmodule