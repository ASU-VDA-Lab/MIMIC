module fake_jpeg_18981_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx2_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_1),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_10),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_49),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_36),
.A2(n_27),
.B1(n_22),
.B2(n_23),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_35),
.B1(n_19),
.B2(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_25),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_46),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_22),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_19),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_52),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_23),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_24),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_57),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_55),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_43),
.B1(n_44),
.B2(n_48),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_61),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_13),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_46),
.C(n_21),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_20),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_50),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_73),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_30),
.Y(n_91)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_43),
.B1(n_40),
.B2(n_44),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_79),
.B1(n_48),
.B2(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_41),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_61),
.B(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_21),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_10),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_78),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_81),
.B(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_85),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_64),
.B(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_74),
.C(n_76),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_48),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_76),
.B(n_79),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_66),
.C(n_75),
.Y(n_93)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_88),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_100),
.C(n_103),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_97),
.B(n_98),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_72),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_87),
.C(n_85),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_102),
.B(n_82),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_77),
.C(n_68),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_89),
.B1(n_68),
.B2(n_81),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_109),
.B1(n_26),
.B2(n_15),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_83),
.C(n_86),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_2),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_84),
.B1(n_88),
.B2(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_110),
.B(n_111),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_80),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_7),
.C(n_8),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_112),
.B(n_8),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_99),
.B(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_116),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_0),
.B(n_2),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_117),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_45),
.B1(n_26),
.B2(n_4),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_119),
.B(n_2),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_123),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_124),
.A2(n_113),
.B(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

OAI31xp33_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_118),
.A3(n_119),
.B(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_127),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_106),
.C(n_4),
.Y(n_128)
);

AOI21x1_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_3),
.B(n_4),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_126),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_132),
.A2(n_133),
.B(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_129),
.B(n_5),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_5),
.Y(n_135)
);


endmodule