module fake_jpeg_2554_n_141 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_0),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_13),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_31),
.B(n_25),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_13),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_0),
.Y(n_51)
);

HAxp5_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_42),
.CON(n_60),
.SN(n_60)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_48),
.Y(n_65)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_42),
.Y(n_69)
);

CKINVDCx6p67_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_48),
.B1(n_36),
.B2(n_39),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_36),
.B1(n_35),
.B2(n_43),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_54),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_43),
.B1(n_36),
.B2(n_39),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_34),
.B(n_32),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_79),
.B1(n_64),
.B2(n_62),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_41),
.B1(n_50),
.B2(n_35),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_70),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_61),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_73),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_44),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_41),
.B1(n_44),
.B2(n_47),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_45),
.B1(n_37),
.B2(n_3),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_26),
.Y(n_88)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_88),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_56),
.C(n_4),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_72),
.C(n_7),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_2),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_4),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_5),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_64),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_5),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_6),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_68),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_102),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_67),
.Y(n_99)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_100),
.B(n_18),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_78),
.B(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_83),
.B1(n_93),
.B2(n_92),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_12),
.C(n_14),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_107),
.B(n_110),
.Y(n_115)
);

INVxp33_ASAP7_75t_SL g109 ( 
.A(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_11),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_12),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_117),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_99),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_118),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_14),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_101),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_96),
.C(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_127),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_120),
.A2(n_103),
.B1(n_123),
.B2(n_100),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_109),
.B1(n_105),
.B2(n_15),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_127),
.A2(n_112),
.B(n_117),
.C(n_121),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_134),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_128),
.B1(n_114),
.B2(n_130),
.Y(n_137)
);

AOI322xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_126),
.A3(n_124),
.B1(n_131),
.B2(n_132),
.C1(n_136),
.C2(n_115),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_19),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_24),
.Y(n_141)
);


endmodule