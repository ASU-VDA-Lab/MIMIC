module fake_netlist_5_71_n_81 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_81);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_81;

wire n_24;
wire n_61;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_38;
wire n_80;
wire n_35;
wire n_73;
wire n_30;
wire n_33;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_27;
wire n_64;
wire n_77;
wire n_28;
wire n_70;
wire n_68;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_8),
.A2(n_4),
.B1(n_14),
.B2(n_6),
.Y(n_26)
);

AND2x4_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_2),
.Y(n_27)
);

CKINVDCx8_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

OA21x2_ASAP7_75t_L g30 ( 
.A1(n_9),
.A2(n_2),
.B(n_7),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_1),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_1),
.B(n_3),
.C(n_6),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_7),
.Y(n_37)
);

AND2x4_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_20),
.B(n_21),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_27),
.B(n_30),
.Y(n_42)
);

OAI21x1_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_34),
.B(n_30),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

OAI21x1_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_34),
.B(n_30),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_46),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_25),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_42),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_44),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_44),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_30),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_57),
.A2(n_47),
.B1(n_51),
.B2(n_23),
.Y(n_60)
);

AOI22x1_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_48),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_48),
.B1(n_50),
.B2(n_36),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_63),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_55),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_55),
.B(n_57),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_33),
.B(n_22),
.C(n_25),
.Y(n_71)
);

OAI221xp5_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_56),
.B1(n_28),
.B2(n_29),
.C(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_66),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_61),
.Y(n_75)
);

OAI311xp33_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_58),
.A3(n_43),
.B1(n_28),
.C1(n_19),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_70),
.B(n_67),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_78),
.A2(n_75),
.B1(n_76),
.B2(n_68),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_75),
.B(n_79),
.Y(n_81)
);


endmodule