module fake_jpeg_24268_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_0),
.B(n_8),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_SL g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_8),
.B(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_22),
.Y(n_34)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_14),
.B1(n_15),
.B2(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_16),
.B(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_4),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_27),
.A2(n_14),
.B1(n_10),
.B2(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_25),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_35),
.B1(n_21),
.B2(n_22),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_13),
.C(n_19),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_20),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_21),
.A2(n_20),
.B1(n_13),
.B2(n_14),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_43),
.B1(n_22),
.B2(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_27),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_46),
.B1(n_38),
.B2(n_24),
.Y(n_58)
);

AOI22x1_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_29),
.C(n_44),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_58),
.B1(n_46),
.B2(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_48),
.B(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_37),
.C(n_51),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_57),
.C(n_19),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_19),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_40),
.C(n_39),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_55),
.B1(n_36),
.B2(n_9),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_61),
.Y(n_65)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

OAI21x1_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_60),
.B(n_63),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_67),
.C(n_6),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_65),
.B1(n_7),
.B2(n_9),
.Y(n_71)
);

BUFx24_ASAP7_75t_SL g70 ( 
.A(n_68),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_71),
.B(n_6),
.Y(n_72)
);


endmodule