module fake_jpeg_13907_n_78 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_78);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx13_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_20),
.B(n_13),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_4),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_40),
.Y(n_43)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_1),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_35),
.C(n_28),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_25),
.C(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_23),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_32),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_26),
.B(n_33),
.C(n_25),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B1(n_22),
.B2(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_2),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_39),
.B1(n_22),
.B2(n_5),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_9),
.B1(n_11),
.B2(n_14),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_66),
.A2(n_6),
.B(n_8),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_69),
.C(n_70),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_65),
.C(n_68),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_62),
.C(n_64),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_62),
.Y(n_75)
);

BUFx24_ASAP7_75t_SL g76 ( 
.A(n_75),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_72),
.C(n_18),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_60),
.Y(n_78)
);


endmodule