module fake_netlist_6_531_n_114 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_20, n_7, n_2, n_5, n_19, n_114);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_114;

wire n_52;
wire n_91;
wire n_46;
wire n_21;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_109;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_110;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_20),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_39)
);

AND2x6_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_17),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_2),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_26),
.B(n_3),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_47),
.B(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_23),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_44),
.B(n_25),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_4),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_50),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

OAI21x1_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_46),
.B(n_45),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_39),
.B(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_40),
.Y(n_65)
);

OAI21x1_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_40),
.B(n_12),
.Y(n_66)
);

OAI21x1_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_40),
.B(n_11),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_R g69 ( 
.A(n_60),
.B(n_13),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_R g70 ( 
.A(n_60),
.B(n_15),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_7),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_7),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_R g74 ( 
.A(n_63),
.B(n_9),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_10),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_R g76 ( 
.A(n_63),
.B(n_10),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_R g77 ( 
.A(n_59),
.B(n_65),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_58),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_61),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_75),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_64),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_64),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_88),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_62),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_65),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_61),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_89),
.B(n_76),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_66),
.B1(n_67),
.B2(n_61),
.Y(n_96)
);

AOI221xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_85),
.B1(n_88),
.B2(n_82),
.C(n_86),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_85),
.B(n_86),
.C(n_82),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_79),
.Y(n_99)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_80),
.Y(n_100)
);

OAI221xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_87),
.B1(n_80),
.B2(n_81),
.C(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_99),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_104),
.A2(n_96),
.B(n_92),
.Y(n_108)
);

OAI211xp5_ASAP7_75t_SL g109 ( 
.A1(n_106),
.A2(n_94),
.B(n_66),
.C(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_R g110 ( 
.A(n_107),
.B(n_102),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_110),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_105),
.B1(n_103),
.B2(n_107),
.Y(n_112)
);

AOI222xp33_ASAP7_75t_SL g113 ( 
.A1(n_112),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.C1(n_67),
.C2(n_81),
.Y(n_113)
);

AOI221xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_81),
.B1(n_53),
.B2(n_33),
.C(n_30),
.Y(n_114)
);


endmodule