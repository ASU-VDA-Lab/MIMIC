module fake_aes_4025_n_503 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_503);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_503;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_73;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g70 ( .A(n_31), .Y(n_70) );
INVx2_ASAP7_75t_L g71 ( .A(n_28), .Y(n_71) );
INVxp67_ASAP7_75t_L g72 ( .A(n_13), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_66), .Y(n_73) );
CKINVDCx16_ASAP7_75t_R g74 ( .A(n_41), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_68), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_62), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_32), .Y(n_77) );
INVxp67_ASAP7_75t_L g78 ( .A(n_40), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_50), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_61), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_42), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_33), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_51), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_48), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_0), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_26), .Y(n_86) );
INVx3_ASAP7_75t_L g87 ( .A(n_36), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_45), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_49), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_30), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_67), .Y(n_91) );
HB1xp67_ASAP7_75t_L g92 ( .A(n_69), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_9), .Y(n_93) );
INVxp67_ASAP7_75t_L g94 ( .A(n_43), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_55), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_35), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_47), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_29), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_3), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_37), .Y(n_100) );
INVxp33_ASAP7_75t_L g101 ( .A(n_18), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_7), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_65), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_23), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_74), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_92), .B(n_0), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_74), .Y(n_107) );
AND2x4_ASAP7_75t_L g108 ( .A(n_87), .B(n_1), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_70), .Y(n_109) );
NOR2xp33_ASAP7_75t_R g110 ( .A(n_79), .B(n_24), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_104), .Y(n_111) );
INVx3_ASAP7_75t_L g112 ( .A(n_87), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_87), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_93), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_72), .Y(n_115) );
OAI22xp5_ASAP7_75t_SL g116 ( .A1(n_101), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_93), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_72), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_87), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_93), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_71), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_82), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_99), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_85), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_99), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_78), .B(n_2), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_71), .Y(n_127) );
NOR2xp67_ASAP7_75t_L g128 ( .A(n_94), .B(n_4), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_112), .B(n_80), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_115), .A2(n_99), .B1(n_102), .B2(n_100), .Y(n_130) );
NAND2x1p5_ASAP7_75t_L g131 ( .A(n_108), .B(n_103), .Y(n_131) );
NAND3x1_ASAP7_75t_L g132 ( .A(n_106), .B(n_116), .C(n_126), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_112), .Y(n_133) );
AND3x4_ASAP7_75t_L g134 ( .A(n_128), .B(n_71), .C(n_81), .Y(n_134) );
NOR2x1p5_ASAP7_75t_L g135 ( .A(n_111), .B(n_103), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_112), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_112), .Y(n_137) );
AO22x2_ASAP7_75t_L g138 ( .A1(n_108), .A2(n_100), .B1(n_97), .B2(n_96), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_108), .Y(n_139) );
INVx4_ASAP7_75t_L g140 ( .A(n_108), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_115), .B(n_86), .Y(n_141) );
INVx2_ASAP7_75t_SL g142 ( .A(n_112), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_113), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_113), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_113), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_108), .B(n_86), .Y(n_146) );
INVx2_ASAP7_75t_SL g147 ( .A(n_119), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_119), .Y(n_148) );
INVx4_ASAP7_75t_SL g149 ( .A(n_114), .Y(n_149) );
AND2x4_ASAP7_75t_L g150 ( .A(n_125), .B(n_88), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_124), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_119), .Y(n_152) );
AND2x2_ASAP7_75t_SL g153 ( .A(n_106), .B(n_88), .Y(n_153) );
NAND2xp33_ASAP7_75t_L g154 ( .A(n_110), .B(n_98), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_121), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_137), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_153), .B(n_110), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_150), .B(n_128), .Y(n_158) );
INVx2_ASAP7_75t_SL g159 ( .A(n_131), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_150), .B(n_118), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_137), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_151), .Y(n_162) );
INVx4_ASAP7_75t_L g163 ( .A(n_149), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_150), .B(n_118), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_131), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_143), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_150), .B(n_125), .Y(n_168) );
NOR2xp33_ASAP7_75t_R g169 ( .A(n_151), .B(n_105), .Y(n_169) );
BUFx12f_ASAP7_75t_L g170 ( .A(n_135), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_152), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_146), .B(n_140), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_153), .B(n_126), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
INVx3_ASAP7_75t_SL g175 ( .A(n_149), .Y(n_175) );
AO22x1_ASAP7_75t_L g176 ( .A1(n_134), .A2(n_96), .B1(n_75), .B2(n_76), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_144), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_141), .B(n_105), .Y(n_179) );
INVx1_ASAP7_75t_SL g180 ( .A(n_131), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_139), .Y(n_181) );
NOR2xp33_ASAP7_75t_R g182 ( .A(n_154), .B(n_107), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_153), .B(n_127), .Y(n_183) );
OR2x2_ASAP7_75t_SL g184 ( .A(n_132), .B(n_109), .Y(n_184) );
NOR3xp33_ASAP7_75t_SL g185 ( .A(n_132), .B(n_122), .C(n_116), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_140), .B(n_90), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_135), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_134), .A2(n_127), .B1(n_121), .B2(n_123), .Y(n_188) );
BUFx2_ASAP7_75t_L g189 ( .A(n_138), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_152), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_175), .Y(n_191) );
OR2x2_ASAP7_75t_L g192 ( .A(n_160), .B(n_130), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_189), .A2(n_138), .B1(n_134), .B2(n_146), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_166), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_166), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_167), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_186), .A2(n_140), .B(n_146), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_157), .A2(n_146), .B(n_129), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_180), .B(n_138), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_165), .B(n_139), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_175), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_160), .B(n_138), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_180), .B(n_144), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_164), .B(n_142), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_167), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_178), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_165), .Y(n_207) );
OAI21xp33_ASAP7_75t_L g208 ( .A1(n_183), .A2(n_148), .B(n_145), .Y(n_208) );
INVx5_ASAP7_75t_L g209 ( .A(n_163), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_178), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_165), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_156), .Y(n_212) );
AND2x6_ASAP7_75t_L g213 ( .A(n_172), .B(n_133), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_172), .Y(n_214) );
NAND3xp33_ASAP7_75t_L g215 ( .A(n_188), .B(n_152), .C(n_148), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_172), .A2(n_136), .B(n_147), .Y(n_216) );
BUFx3_ASAP7_75t_L g217 ( .A(n_175), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_169), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_156), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_161), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_161), .Y(n_221) );
BUFx10_ASAP7_75t_L g222 ( .A(n_159), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_188), .A2(n_145), .B1(n_147), .B2(n_155), .Y(n_223) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_193), .A2(n_159), .B1(n_184), .B2(n_168), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_195), .B(n_164), .Y(n_225) );
CKINVDCx11_ASAP7_75t_R g226 ( .A(n_222), .Y(n_226) );
OAI221xp5_ASAP7_75t_L g227 ( .A1(n_193), .A2(n_185), .B1(n_179), .B2(n_173), .C(n_168), .Y(n_227) );
OAI221xp5_ASAP7_75t_L g228 ( .A1(n_192), .A2(n_173), .B1(n_202), .B2(n_204), .C(n_223), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_214), .A2(n_172), .B1(n_162), .B2(n_170), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_198), .A2(n_158), .B(n_177), .Y(n_230) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_215), .A2(n_89), .B(n_81), .Y(n_231) );
OAI222xp33_ASAP7_75t_L g232 ( .A1(n_218), .A2(n_158), .B1(n_184), .B2(n_187), .C1(n_176), .C2(n_77), .Y(n_232) );
AOI221x1_ASAP7_75t_L g233 ( .A1(n_215), .A2(n_158), .B1(n_75), .B2(n_76), .C(n_77), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_207), .B(n_174), .Y(n_234) );
NAND2xp33_ASAP7_75t_SL g235 ( .A(n_191), .B(n_182), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_207), .Y(n_236) );
NAND2xp33_ASAP7_75t_R g237 ( .A(n_199), .B(n_158), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_192), .A2(n_181), .B(n_174), .C(n_155), .Y(n_238) );
CKINVDCx11_ASAP7_75t_R g239 ( .A(n_222), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_194), .A2(n_181), .B(n_174), .C(n_127), .Y(n_240) );
AOI22xp33_ASAP7_75t_SL g241 ( .A1(n_199), .A2(n_170), .B1(n_176), .B2(n_174), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_214), .A2(n_170), .B1(n_152), .B2(n_84), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_223), .A2(n_127), .B1(n_121), .B2(n_120), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_195), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_214), .A2(n_152), .B1(n_83), .B2(n_84), .Y(n_245) );
OAI221xp5_ASAP7_75t_L g246 ( .A1(n_214), .A2(n_114), .B1(n_117), .B2(n_120), .C(n_123), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_195), .B(n_127), .Y(n_247) );
BUFx2_ASAP7_75t_L g248 ( .A(n_213), .Y(n_248) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_194), .A2(n_190), .B(n_177), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_244), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_227), .B(n_232), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_244), .Y(n_252) );
OAI22xp33_ASAP7_75t_L g253 ( .A1(n_224), .A2(n_205), .B1(n_206), .B2(n_207), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_247), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_225), .B(n_196), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_224), .A2(n_200), .B1(n_210), .B2(n_196), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_227), .A2(n_200), .B1(n_210), .B2(n_213), .Y(n_257) );
OAI22xp33_ASAP7_75t_L g258 ( .A1(n_237), .A2(n_206), .B1(n_205), .B2(n_220), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_229), .B(n_211), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_247), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_228), .A2(n_205), .B1(n_206), .B2(n_220), .Y(n_261) );
AOI21x1_ASAP7_75t_L g262 ( .A1(n_231), .A2(n_221), .B(n_220), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_228), .A2(n_203), .B1(n_221), .B2(n_219), .Y(n_263) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_230), .A2(n_208), .B(n_216), .Y(n_264) );
OR2x2_ASAP7_75t_L g265 ( .A(n_225), .B(n_212), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_241), .A2(n_200), .B1(n_213), .B2(n_211), .Y(n_266) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_230), .A2(n_212), .B(n_221), .Y(n_267) );
OAI211xp5_ASAP7_75t_L g268 ( .A1(n_226), .A2(n_212), .B(n_219), .C(n_203), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_246), .A2(n_200), .B1(n_213), .B2(n_211), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_243), .B(n_219), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_246), .A2(n_213), .B1(n_211), .B2(n_208), .Y(n_271) );
AO21x2_ASAP7_75t_L g272 ( .A1(n_261), .A2(n_249), .B(n_243), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_250), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_250), .B(n_231), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_265), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_267), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g277 ( .A1(n_263), .A2(n_233), .B(n_238), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_267), .Y(n_278) );
NAND2xp33_ASAP7_75t_R g279 ( .A(n_251), .B(n_236), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_261), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_252), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_252), .B(n_231), .Y(n_282) );
NAND2xp33_ASAP7_75t_R g283 ( .A(n_265), .B(n_248), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_262), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g285 ( .A1(n_256), .A2(n_117), .B1(n_242), .B2(n_245), .C(n_235), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_262), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_257), .A2(n_239), .B1(n_248), .B2(n_234), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_255), .Y(n_288) );
BUFx10_ASAP7_75t_L g289 ( .A(n_259), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_264), .Y(n_290) );
INVxp67_ASAP7_75t_L g291 ( .A(n_255), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_254), .B(n_231), .Y(n_292) );
INVx5_ASAP7_75t_L g293 ( .A(n_254), .Y(n_293) );
BUFx2_ASAP7_75t_L g294 ( .A(n_284), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_284), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_273), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_275), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_286), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_274), .B(n_263), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_274), .B(n_264), .Y(n_300) );
HB1xp67_ASAP7_75t_SL g301 ( .A(n_280), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_276), .Y(n_302) );
AOI221xp5_ASAP7_75t_L g303 ( .A1(n_291), .A2(n_258), .B1(n_253), .B2(n_268), .C(n_266), .Y(n_303) );
CKINVDCx16_ASAP7_75t_R g304 ( .A(n_283), .Y(n_304) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_277), .A2(n_233), .B(n_268), .Y(n_305) );
NOR4xp25_ASAP7_75t_L g306 ( .A(n_291), .B(n_97), .C(n_83), .D(n_90), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_273), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_286), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_281), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_281), .B(n_270), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_288), .B(n_270), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_274), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_280), .B(n_264), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_282), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_279), .B(n_73), .C(n_91), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_293), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_282), .Y(n_317) );
INVxp67_ASAP7_75t_SL g318 ( .A(n_276), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_272), .B(n_254), .Y(n_319) );
AOI21xp33_ASAP7_75t_L g320 ( .A1(n_277), .A2(n_260), .B(n_271), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_276), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_293), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_288), .A2(n_269), .B1(n_260), .B2(n_240), .Y(n_323) );
INVxp33_ASAP7_75t_L g324 ( .A(n_287), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_278), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_296), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_312), .B(n_272), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_312), .B(n_290), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_299), .B(n_272), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_296), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_295), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_295), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_317), .B(n_272), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_324), .A2(n_289), .B1(n_285), .B2(n_293), .Y(n_334) );
AOI31xp33_ASAP7_75t_L g335 ( .A1(n_315), .A2(n_285), .A3(n_292), .B(n_73), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_307), .Y(n_336) );
OAI31xp33_ASAP7_75t_L g337 ( .A1(n_315), .A2(n_91), .A3(n_95), .B(n_81), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_300), .B(n_290), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_307), .B(n_293), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_295), .Y(n_340) );
NOR2xp67_ASAP7_75t_SL g341 ( .A(n_304), .B(n_293), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_309), .B(n_293), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_299), .B(n_278), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_317), .B(n_278), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_311), .B(n_293), .Y(n_345) );
NAND4xp25_ASAP7_75t_SL g346 ( .A(n_297), .B(n_95), .C(n_292), .D(n_89), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_314), .B(n_290), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_299), .B(n_289), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_314), .B(n_260), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_298), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_316), .Y(n_351) );
NAND2x1p5_ASAP7_75t_L g352 ( .A(n_322), .B(n_217), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_319), .B(n_289), .Y(n_353) );
OR2x6_ASAP7_75t_L g354 ( .A(n_322), .B(n_289), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_298), .Y(n_355) );
NAND3xp33_ASAP7_75t_SL g356 ( .A(n_306), .B(n_89), .C(n_5), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_319), .B(n_4), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_319), .B(n_5), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_300), .B(n_6), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_297), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_303), .A2(n_234), .B1(n_213), .B2(n_249), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_310), .B(n_6), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_300), .B(n_7), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_313), .B(n_8), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_310), .B(n_8), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_311), .B(n_9), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_294), .B(n_10), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_298), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_306), .B(n_10), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_346), .A2(n_303), .B(n_305), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_359), .B(n_313), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_335), .A2(n_301), .B1(n_305), .B2(n_322), .Y(n_372) );
A2O1A1Ixp33_ASAP7_75t_L g373 ( .A1(n_337), .A2(n_294), .B(n_308), .C(n_320), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_326), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_361), .A2(n_320), .B1(n_323), .B2(n_313), .Y(n_375) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_356), .A2(n_308), .B(n_323), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_354), .A2(n_318), .B(n_325), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_334), .A2(n_362), .B1(n_365), .B2(n_301), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_360), .B(n_302), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_351), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_362), .A2(n_318), .B1(n_302), .B2(n_325), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_344), .Y(n_382) );
OAI221xp5_ASAP7_75t_SL g383 ( .A1(n_365), .A2(n_321), .B1(n_302), .B2(n_197), .C(n_14), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_366), .B(n_11), .Y(n_384) );
AOI32xp33_ASAP7_75t_L g385 ( .A1(n_363), .A2(n_302), .A3(n_321), .B1(n_234), .B2(n_14), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_369), .A2(n_321), .B1(n_234), .B2(n_213), .Y(n_386) );
AOI21xp33_ASAP7_75t_L g387 ( .A1(n_367), .A2(n_11), .B(n_12), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_363), .A2(n_213), .B1(n_222), .B2(n_209), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_364), .B(n_12), .Y(n_389) );
AOI21xp33_ASAP7_75t_L g390 ( .A1(n_333), .A2(n_13), .B(n_15), .Y(n_390) );
NOR2x1_ASAP7_75t_L g391 ( .A(n_354), .B(n_217), .Y(n_391) );
INVxp67_ASAP7_75t_L g392 ( .A(n_341), .Y(n_392) );
AOI22x1_ASAP7_75t_L g393 ( .A1(n_357), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_345), .B(n_16), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_364), .B(n_17), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_341), .A2(n_209), .B1(n_217), .B2(n_201), .Y(n_396) );
XOR2x2_ASAP7_75t_L g397 ( .A(n_358), .B(n_348), .Y(n_397) );
NAND2x1_ASAP7_75t_L g398 ( .A(n_354), .B(n_201), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_358), .B(n_201), .Y(n_399) );
AOI311xp33_ASAP7_75t_L g400 ( .A1(n_330), .A2(n_18), .A3(n_19), .B(n_20), .C(n_21), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_343), .B(n_19), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_329), .B(n_20), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_354), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_339), .B(n_201), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_336), .Y(n_405) );
INVx2_ASAP7_75t_SL g406 ( .A(n_352), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_329), .B(n_21), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_348), .B(n_22), .Y(n_408) );
NAND2x1p5_ASAP7_75t_L g409 ( .A(n_349), .B(n_201), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_344), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_342), .B(n_191), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_331), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_353), .B(n_25), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_336), .Y(n_414) );
AOI32xp33_ASAP7_75t_L g415 ( .A1(n_353), .A2(n_27), .A3(n_34), .B1(n_38), .B2(n_39), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_380), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_412), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_398), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_372), .B(n_332), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_374), .Y(n_420) );
NOR3xp33_ASAP7_75t_L g421 ( .A(n_402), .B(n_333), .C(n_327), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_410), .B(n_338), .Y(n_422) );
OAI21xp5_ASAP7_75t_SL g423 ( .A1(n_372), .A2(n_352), .B(n_338), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_371), .B(n_338), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_382), .B(n_338), .Y(n_425) );
AOI32xp33_ASAP7_75t_L g426 ( .A1(n_378), .A2(n_328), .A3(n_355), .B1(n_368), .B2(n_350), .Y(n_426) );
NOR3xp33_ASAP7_75t_SL g427 ( .A(n_370), .B(n_368), .C(n_328), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_407), .B(n_328), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_405), .Y(n_429) );
NOR2xp33_ASAP7_75t_R g430 ( .A(n_403), .B(n_347), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_414), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_403), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_391), .B(n_350), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_409), .Y(n_434) );
NOR3xp33_ASAP7_75t_L g435 ( .A(n_390), .B(n_347), .C(n_340), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_373), .A2(n_332), .B(n_331), .Y(n_436) );
NAND2xp33_ASAP7_75t_SL g437 ( .A(n_406), .B(n_340), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_401), .Y(n_438) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_377), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_381), .Y(n_440) );
NOR2x1_ASAP7_75t_L g441 ( .A(n_376), .B(n_191), .Y(n_441) );
NAND2xp33_ASAP7_75t_SL g442 ( .A(n_397), .B(n_191), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_394), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_392), .B(n_191), .Y(n_444) );
AOI211x1_ASAP7_75t_L g445 ( .A1(n_387), .A2(n_395), .B(n_389), .C(n_376), .Y(n_445) );
OAI21xp33_ASAP7_75t_SL g446 ( .A1(n_385), .A2(n_163), .B(n_46), .Y(n_446) );
INVxp67_ASAP7_75t_L g447 ( .A(n_379), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_409), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_399), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_375), .B(n_44), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_404), .Y(n_451) );
AOI21xp33_ASAP7_75t_L g452 ( .A1(n_446), .A2(n_384), .B(n_393), .Y(n_452) );
INVx1_ASAP7_75t_SL g453 ( .A(n_430), .Y(n_453) );
OAI22xp33_ASAP7_75t_L g454 ( .A1(n_423), .A2(n_388), .B1(n_386), .B2(n_413), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_426), .B(n_400), .C(n_415), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g456 ( .A1(n_441), .A2(n_383), .B(n_408), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_440), .B(n_411), .Y(n_457) );
XNOR2xp5_ASAP7_75t_L g458 ( .A(n_443), .B(n_396), .Y(n_458) );
CKINVDCx6p67_ASAP7_75t_R g459 ( .A(n_418), .Y(n_459) );
NOR2x1_ASAP7_75t_L g460 ( .A(n_418), .B(n_163), .Y(n_460) );
O2A1O1Ixp5_ASAP7_75t_SL g461 ( .A1(n_419), .A2(n_52), .B(n_53), .C(n_54), .Y(n_461) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_427), .A2(n_209), .B(n_190), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_439), .B(n_56), .Y(n_463) );
XNOR2xp5_ASAP7_75t_L g464 ( .A(n_438), .B(n_57), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_425), .B(n_58), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_420), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_429), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_430), .B(n_59), .Y(n_468) );
XNOR2x2_ASAP7_75t_L g469 ( .A(n_419), .B(n_60), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_442), .A2(n_209), .B(n_171), .Y(n_470) );
AOI322xp5_ASAP7_75t_L g471 ( .A1(n_453), .A2(n_416), .A3(n_421), .B1(n_437), .B2(n_424), .C1(n_428), .C2(n_422), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_455), .A2(n_445), .B1(n_428), .B2(n_447), .C(n_435), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_452), .B(n_431), .Y(n_473) );
OAI21xp33_ASAP7_75t_L g474 ( .A1(n_458), .A2(n_432), .B(n_449), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_457), .B(n_467), .Y(n_475) );
NAND2xp33_ASAP7_75t_L g476 ( .A(n_464), .B(n_433), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_457), .B(n_436), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_452), .A2(n_433), .B(n_448), .C(n_444), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_SL g479 ( .A1(n_454), .A2(n_444), .B(n_450), .C(n_432), .Y(n_479) );
NOR2x1_ASAP7_75t_L g480 ( .A(n_454), .B(n_434), .Y(n_480) );
NAND3xp33_ASAP7_75t_L g481 ( .A(n_463), .B(n_451), .C(n_434), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_459), .Y(n_482) );
OAI21xp5_ASAP7_75t_SL g483 ( .A1(n_456), .A2(n_417), .B(n_63), .Y(n_483) );
OAI21x1_ASAP7_75t_SL g484 ( .A1(n_469), .A2(n_417), .B(n_64), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_466), .Y(n_485) );
INVxp33_ASAP7_75t_SL g486 ( .A(n_468), .Y(n_486) );
OAI221xp5_ASAP7_75t_L g487 ( .A1(n_470), .A2(n_149), .B1(n_462), .B2(n_460), .C(n_465), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_470), .A2(n_454), .B1(n_455), .B2(n_453), .Y(n_488) );
NOR4xp25_ASAP7_75t_L g489 ( .A(n_461), .B(n_360), .C(n_455), .D(n_453), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_459), .Y(n_490) );
NAND4xp75_ASAP7_75t_L g491 ( .A(n_480), .B(n_488), .C(n_472), .D(n_473), .Y(n_491) );
NAND3xp33_ASAP7_75t_SL g492 ( .A(n_489), .B(n_478), .C(n_490), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_475), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_477), .B(n_473), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_485), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_494), .B(n_471), .Y(n_496) );
AO22x2_ASAP7_75t_L g497 ( .A1(n_491), .A2(n_484), .B1(n_481), .B2(n_483), .Y(n_497) );
AOI22xp33_ASAP7_75t_SL g498 ( .A1(n_493), .A2(n_482), .B1(n_486), .B2(n_476), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_496), .B(n_492), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_498), .B(n_495), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_500), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_501), .A2(n_492), .B1(n_499), .B2(n_497), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_L g503 ( .A1(n_502), .A2(n_479), .B(n_474), .C(n_487), .Y(n_503) );
endmodule