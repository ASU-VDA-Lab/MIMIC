module real_jpeg_23334_n_3 (n_1, n_0, n_2, n_3);

input n_1;
input n_0;
input n_2;

output n_3;

wire n_5;
wire n_4;
wire n_6;
wire n_7;

AO21x1_ASAP7_75t_L g3 ( 
.A1(n_0),
.A2(n_4),
.B(n_7),
.Y(n_3)
);

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_1),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g5 ( 
.A(n_2),
.Y(n_5)
);

NAND2xp5_ASAP7_75t_L g4 ( 
.A(n_5),
.B(n_6),
.Y(n_4)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_5),
.B(n_6),
.Y(n_7)
);


endmodule