module real_jpeg_13201_n_3 (n_1, n_0, n_2, n_3);

input n_1;
input n_0;
input n_2;

output n_3;

wire n_5;
wire n_4;
wire n_8;
wire n_6;
wire n_7;

NAND2xp5_ASAP7_75t_L g5 ( 
.A(n_0),
.B(n_2),
.Y(n_5)
);

OAI21xp5_ASAP7_75t_L g3 ( 
.A1(n_1),
.A2(n_4),
.B(n_6),
.Y(n_3)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVxp67_ASAP7_75t_L g4 ( 
.A(n_5),
.Y(n_4)
);

NOR2xp33_ASAP7_75t_SL g7 ( 
.A(n_5),
.B(n_8),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_7),
.Y(n_6)
);


endmodule