module fake_jpeg_7185_n_77 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_77);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_13),
.B(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_SL g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_53),
.Y(n_60)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_57),
.B1(n_48),
.B2(n_46),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_0),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_61)
);

NOR4xp25_ASAP7_75t_SL g55 ( 
.A(n_34),
.B(n_14),
.C(n_2),
.D(n_3),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_0),
.B1(n_5),
.B2(n_7),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_33),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_58)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_65),
.Y(n_68)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_62),
.B1(n_60),
.B2(n_40),
.Y(n_69)
);

NOR2xp67_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_70),
.B(n_61),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_68),
.C(n_36),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_72),
.A2(n_35),
.B1(n_19),
.B2(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_74),
.B(n_32),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_12),
.B1(n_26),
.B2(n_28),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_30),
.Y(n_77)
);


endmodule