module real_jpeg_24030_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_1),
.A2(n_19),
.B1(n_20),
.B2(n_25),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_1),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_2),
.A2(n_19),
.B1(n_20),
.B2(n_45),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_45),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_2),
.A2(n_23),
.B1(n_26),
.B2(n_45),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_4),
.A2(n_23),
.B1(n_26),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_4),
.A2(n_32),
.B1(n_39),
.B2(n_40),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_4),
.A2(n_18),
.B(n_26),
.C(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_4),
.B(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_4),
.A2(n_19),
.B1(n_20),
.B2(n_32),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_4),
.B(n_38),
.C(n_39),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_4),
.B(n_16),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_4),
.B(n_9),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_4),
.B(n_36),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_9),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_87),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_85),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_58),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_13),
.B(n_58),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_33),
.C(n_46),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_14),
.B(n_33),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_27),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_22),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_17),
.B(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_17)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_21),
.B1(n_23),
.B2(n_26),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_19),
.A2(n_20),
.B1(n_37),
.B2(n_38),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_19),
.A2(n_21),
.B(n_32),
.Y(n_56)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_20),
.B(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_SL g75 ( 
.A(n_22),
.Y(n_75)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_23),
.A2(n_26),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_29),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_41),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_34),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_35),
.B(n_42),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_36),
.B(n_44),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_39),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_39),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_42),
.B(n_81),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_46),
.B(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_55),
.B2(n_57),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_55),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B(n_54),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_49),
.B(n_110),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_49),
.B(n_69),
.Y(n_116)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_53),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_55),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_76),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_71),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_66),
.B(n_109),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_84),
.B(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_134),
.B(n_138),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_113),
.B(n_133),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_96),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_90),
.B(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_93),
.B1(n_94),
.B2(n_121),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_91),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_104),
.B2(n_112),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_99),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_103),
.C(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_111),
.B(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_122),
.B(n_132),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_120),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_128),
.B(n_131),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_129),
.B(n_130),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_135),
.B(n_136),
.Y(n_138)
);


endmodule