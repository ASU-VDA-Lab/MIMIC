module fake_jpeg_23753_n_38 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_38);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_10),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_15),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_5),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_7),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_16),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_19),
.B(n_22),
.C(n_0),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_32),
.B(n_30),
.C(n_12),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_1),
.B(n_4),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_29),
.C(n_31),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_34),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_37),
.Y(n_38)
);


endmodule