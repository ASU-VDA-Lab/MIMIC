module fake_aes_10084_n_631 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_631);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_631;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_L g86 ( .A(n_44), .Y(n_86) );
BUFx3_ASAP7_75t_L g87 ( .A(n_72), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_83), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_23), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_63), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_35), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_24), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_69), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_62), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_43), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_28), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_32), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_2), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_21), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_7), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_67), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_17), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_74), .Y(n_103) );
BUFx2_ASAP7_75t_L g104 ( .A(n_77), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_10), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_45), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_55), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_47), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_70), .Y(n_109) );
INVxp67_ASAP7_75t_L g110 ( .A(n_50), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_59), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_18), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_26), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_76), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_41), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_51), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_17), .Y(n_118) );
XNOR2x1_ASAP7_75t_L g119 ( .A(n_15), .B(n_16), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_18), .Y(n_120) );
CKINVDCx14_ASAP7_75t_R g121 ( .A(n_33), .Y(n_121) );
INVx2_ASAP7_75t_SL g122 ( .A(n_64), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_48), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_20), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_27), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_40), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_21), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_58), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_92), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_92), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_126), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_93), .Y(n_132) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_89), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_104), .B(n_0), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_112), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_126), .Y(n_136) );
BUFx8_ASAP7_75t_L g137 ( .A(n_104), .Y(n_137) );
NOR2xp33_ASAP7_75t_R g138 ( .A(n_121), .B(n_37), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_120), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_87), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_94), .Y(n_142) );
INVx6_ASAP7_75t_L g143 ( .A(n_87), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_122), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_122), .B(n_1), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_112), .B(n_3), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_94), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_91), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_89), .B(n_3), .Y(n_149) );
NOR2xp33_ASAP7_75t_SL g150 ( .A(n_106), .B(n_39), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_107), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_115), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_98), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_119), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_140), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g156 ( .A1(n_134), .A2(n_119), .B1(n_127), .B2(n_102), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_140), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_141), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_144), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_140), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_134), .Y(n_161) );
BUFx4f_ASAP7_75t_L g162 ( .A(n_134), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_148), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_147), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_129), .B(n_86), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_134), .B(n_99), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_147), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_147), .Y(n_168) );
INVx4_ASAP7_75t_L g169 ( .A(n_146), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_131), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_141), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_131), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_131), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_129), .B(n_99), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_130), .B(n_110), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_146), .Y(n_177) );
INVxp67_ASAP7_75t_L g178 ( .A(n_133), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_146), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_146), .Y(n_180) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_137), .Y(n_181) );
INVx4_ASAP7_75t_SL g182 ( .A(n_143), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_141), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
NAND2xp33_ASAP7_75t_L g185 ( .A(n_138), .B(n_97), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_162), .A2(n_145), .B(n_132), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_169), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_162), .B(n_137), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_155), .Y(n_189) );
NAND2xp33_ASAP7_75t_L g190 ( .A(n_181), .B(n_144), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
NOR3xp33_ASAP7_75t_SL g192 ( .A(n_163), .B(n_152), .C(n_151), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_161), .B(n_137), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_181), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_159), .Y(n_195) );
AOI22xp33_ASAP7_75t_SL g196 ( .A1(n_166), .A2(n_137), .B1(n_124), .B2(n_150), .Y(n_196) );
NOR3xp33_ASAP7_75t_L g197 ( .A(n_178), .B(n_149), .C(n_154), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_162), .A2(n_132), .B1(n_142), .B2(n_130), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_174), .B(n_142), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_178), .B(n_111), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_157), .Y(n_201) );
NOR2x1p5_ASAP7_75t_L g202 ( .A(n_161), .B(n_154), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_157), .Y(n_203) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_162), .Y(n_204) );
BUFx2_ASAP7_75t_L g205 ( .A(n_161), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_176), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_161), .B(n_136), .Y(n_207) );
BUFx4f_ASAP7_75t_L g208 ( .A(n_180), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_176), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_169), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_161), .B(n_136), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_160), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_160), .Y(n_213) );
BUFx4f_ASAP7_75t_L g214 ( .A(n_180), .Y(n_214) );
INVx2_ASAP7_75t_SL g215 ( .A(n_174), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_164), .Y(n_216) );
BUFx4f_ASAP7_75t_L g217 ( .A(n_180), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_169), .A2(n_144), .B1(n_143), .B2(n_100), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_164), .Y(n_219) );
INVx2_ASAP7_75t_SL g220 ( .A(n_174), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_167), .Y(n_221) );
AOI22xp33_ASAP7_75t_SL g222 ( .A1(n_166), .A2(n_100), .B1(n_135), .B2(n_118), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_169), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_169), .B(n_97), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_177), .B(n_103), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_176), .Y(n_226) );
OAI222xp33_ASAP7_75t_L g227 ( .A1(n_196), .A2(n_139), .B1(n_156), .B2(n_153), .C1(n_166), .C2(n_179), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_202), .A2(n_180), .B1(n_177), .B2(n_179), .Y(n_228) );
BUFx3_ASAP7_75t_L g229 ( .A(n_195), .Y(n_229) );
NAND2x1p5_ASAP7_75t_L g230 ( .A(n_215), .B(n_167), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_215), .B(n_156), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_186), .A2(n_165), .B(n_175), .Y(n_232) );
BUFx4f_ASAP7_75t_L g233 ( .A(n_220), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_186), .A2(n_165), .B(n_175), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_199), .B(n_168), .Y(n_235) );
AOI222xp33_ASAP7_75t_L g236 ( .A1(n_202), .A2(n_105), .B1(n_114), .B2(n_135), .C1(n_168), .C2(n_185), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_208), .B(n_184), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_195), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_197), .B(n_139), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_220), .A2(n_172), .B1(n_170), .B2(n_173), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_198), .A2(n_196), .B1(n_193), .B2(n_199), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_207), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_188), .B(n_182), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_194), .A2(n_128), .B1(n_113), .B2(n_103), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_207), .A2(n_184), .B(n_159), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_204), .B(n_113), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_200), .B(n_170), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_187), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_193), .B(n_182), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_187), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_205), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_211), .A2(n_184), .B(n_159), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_205), .Y(n_253) );
AND3x1_ASAP7_75t_SL g254 ( .A(n_192), .B(n_116), .C(n_95), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_222), .A2(n_128), .B1(n_172), .B2(n_173), .Y(n_255) );
INVxp67_ASAP7_75t_L g256 ( .A(n_224), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_195), .Y(n_257) );
AOI221xp5_ASAP7_75t_L g258 ( .A1(n_222), .A2(n_135), .B1(n_144), .B2(n_96), .C(n_101), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_187), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_208), .B(n_184), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_224), .B(n_135), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_189), .A2(n_143), .B1(n_141), .B2(n_101), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_189), .B(n_143), .Y(n_263) );
BUFx12f_ASAP7_75t_L g264 ( .A(n_209), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_191), .B(n_182), .Y(n_265) );
BUFx12f_ASAP7_75t_L g266 ( .A(n_209), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_211), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_233), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_242), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_248), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_232), .A2(n_226), .B(n_206), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_234), .A2(n_213), .B(n_201), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_233), .Y(n_273) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_261), .A2(n_116), .B(n_95), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_230), .B(n_191), .Y(n_275) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_241), .A2(n_226), .B(n_206), .Y(n_276) );
OAI21x1_ASAP7_75t_L g277 ( .A1(n_263), .A2(n_226), .B(n_206), .Y(n_277) );
AOI21x1_ASAP7_75t_L g278 ( .A1(n_265), .A2(n_183), .B(n_171), .Y(n_278) );
NOR4xp25_ASAP7_75t_L g279 ( .A(n_227), .B(n_125), .C(n_96), .D(n_88), .Y(n_279) );
OAI21x1_ASAP7_75t_L g280 ( .A1(n_240), .A2(n_171), .B(n_183), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_230), .A2(n_171), .B(n_183), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_248), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_250), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_267), .B(n_201), .Y(n_284) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_262), .A2(n_158), .B(n_213), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_250), .Y(n_286) );
BUFx3_ASAP7_75t_L g287 ( .A(n_266), .Y(n_287) );
OAI221xp5_ASAP7_75t_L g288 ( .A1(n_228), .A2(n_225), .B1(n_203), .B2(n_221), .C(n_219), .Y(n_288) );
CKINVDCx8_ASAP7_75t_R g289 ( .A(n_251), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_238), .B(n_203), .Y(n_290) );
A2O1A1Ixp33_ASAP7_75t_L g291 ( .A1(n_256), .A2(n_216), .B(n_212), .C(n_219), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_259), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_259), .Y(n_293) );
AO21x2_ASAP7_75t_L g294 ( .A1(n_245), .A2(n_158), .B(n_125), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_231), .A2(n_216), .B1(n_221), .B2(n_212), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_262), .A2(n_158), .B(n_108), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_235), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_239), .A2(n_208), .B1(n_214), .B2(n_217), .Y(n_298) );
OA21x2_ASAP7_75t_L g299 ( .A1(n_258), .A2(n_109), .B(n_117), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_253), .B(n_223), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_287), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_297), .A2(n_231), .B1(n_236), .B2(n_228), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_297), .B(n_269), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_297), .B(n_247), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_287), .Y(n_305) );
OR2x6_ASAP7_75t_L g306 ( .A(n_287), .B(n_253), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_288), .A2(n_246), .B1(n_217), .B2(n_208), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_295), .B(n_255), .Y(n_308) );
AOI222xp33_ASAP7_75t_L g309 ( .A1(n_269), .A2(n_246), .B1(n_217), .B2(n_214), .C1(n_190), .C2(n_90), .Y(n_309) );
AOI21xp33_ASAP7_75t_L g310 ( .A1(n_288), .A2(n_249), .B(n_243), .Y(n_310) );
OAI221xp5_ASAP7_75t_L g311 ( .A1(n_279), .A2(n_244), .B1(n_217), .B2(n_214), .C(n_218), .Y(n_311) );
OAI22xp33_ASAP7_75t_L g312 ( .A1(n_289), .A2(n_214), .B1(n_254), .B2(n_266), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_287), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_272), .A2(n_260), .B(n_237), .Y(n_314) );
OAI222xp33_ASAP7_75t_L g315 ( .A1(n_289), .A2(n_254), .B1(n_123), .B2(n_260), .C1(n_237), .C2(n_243), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_295), .A2(n_229), .B1(n_257), .B2(n_238), .Y(n_316) );
OAI211xp5_ASAP7_75t_SL g317 ( .A1(n_289), .A2(n_252), .B(n_210), .C(n_223), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_284), .B(n_187), .Y(n_318) );
INVxp67_ASAP7_75t_L g319 ( .A(n_284), .Y(n_319) );
AO31x2_ASAP7_75t_L g320 ( .A1(n_291), .A2(n_141), .A3(n_176), .B(n_264), .Y(n_320) );
AOI22xp33_ASAP7_75t_SL g321 ( .A1(n_299), .A2(n_229), .B1(n_238), .B2(n_257), .Y(n_321) );
OAI221xp5_ASAP7_75t_L g322 ( .A1(n_279), .A2(n_210), .B1(n_223), .B2(n_141), .C(n_238), .Y(n_322) );
OA21x2_ASAP7_75t_L g323 ( .A1(n_276), .A2(n_249), .B(n_176), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_284), .B(n_223), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_291), .B(n_210), .Y(n_325) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_275), .B(n_257), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_300), .A2(n_210), .B1(n_257), .B2(n_176), .Y(n_327) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_298), .A2(n_176), .B1(n_209), .B2(n_6), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_303), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_323), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_320), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_319), .B(n_274), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_323), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_304), .B(n_272), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_320), .Y(n_335) );
AND2x2_ASAP7_75t_SL g336 ( .A(n_308), .B(n_274), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_302), .A2(n_299), .B1(n_274), .B2(n_294), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_323), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_320), .Y(n_339) );
BUFx6f_ASAP7_75t_SL g340 ( .A(n_313), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_320), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_318), .B(n_274), .Y(n_342) );
INVxp67_ASAP7_75t_SL g343 ( .A(n_316), .Y(n_343) );
INVx5_ASAP7_75t_L g344 ( .A(n_313), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_314), .B(n_276), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_326), .Y(n_346) );
INVxp67_ASAP7_75t_SL g347 ( .A(n_304), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_318), .B(n_274), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_308), .B(n_274), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_306), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_324), .B(n_270), .Y(n_351) );
INVxp67_ASAP7_75t_L g352 ( .A(n_301), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_306), .B(n_276), .Y(n_353) );
AO31x2_ASAP7_75t_L g354 ( .A1(n_325), .A2(n_270), .A3(n_282), .B(n_283), .Y(n_354) );
INVx4_ASAP7_75t_L g355 ( .A(n_313), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_342), .B(n_348), .Y(n_356) );
AND2x4_ASAP7_75t_SL g357 ( .A(n_355), .B(n_313), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_354), .Y(n_358) );
NAND4xp25_ASAP7_75t_L g359 ( .A(n_337), .B(n_307), .C(n_322), .D(n_309), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_347), .Y(n_360) );
AND2x4_ASAP7_75t_SL g361 ( .A(n_355), .B(n_306), .Y(n_361) );
OAI21xp5_ASAP7_75t_L g362 ( .A1(n_337), .A2(n_315), .B(n_312), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_330), .A2(n_275), .B(n_321), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_344), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_354), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_342), .B(n_294), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_347), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_350), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_354), .Y(n_369) );
NAND2xp33_ASAP7_75t_R g370 ( .A(n_342), .B(n_305), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_352), .Y(n_371) );
OR2x2_ASAP7_75t_SL g372 ( .A(n_350), .B(n_299), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_354), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_353), .B(n_294), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_348), .B(n_294), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_354), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_354), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_354), .Y(n_378) );
INVx4_ASAP7_75t_L g379 ( .A(n_344), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_336), .A2(n_311), .B1(n_310), .B2(n_317), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_329), .B(n_305), .Y(n_381) );
INVx2_ASAP7_75t_SL g382 ( .A(n_344), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_349), .B(n_306), .Y(n_383) );
AOI222xp33_ASAP7_75t_SL g384 ( .A1(n_329), .A2(n_4), .B1(n_5), .B2(n_7), .C1(n_8), .C2(n_9), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_352), .B(n_268), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_349), .B(n_294), .Y(n_386) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_330), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_351), .B(n_324), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_356), .B(n_331), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_358), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_356), .B(n_331), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_366), .B(n_375), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_366), .B(n_335), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_375), .B(n_335), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_374), .B(n_365), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_360), .B(n_349), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_367), .B(n_334), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_374), .B(n_358), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_381), .B(n_268), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_374), .B(n_339), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_374), .B(n_341), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_358), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_365), .B(n_334), .Y(n_403) );
NOR2xp67_ASAP7_75t_L g404 ( .A(n_379), .B(n_333), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_369), .B(n_341), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_379), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_369), .B(n_332), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_373), .B(n_333), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_373), .B(n_332), .Y(n_409) );
NAND3xp33_ASAP7_75t_SL g410 ( .A(n_384), .B(n_332), .C(n_273), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_386), .B(n_338), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_378), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_386), .B(n_338), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_383), .B(n_353), .Y(n_414) );
INVxp67_ASAP7_75t_L g415 ( .A(n_387), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_371), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_376), .B(n_339), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_376), .B(n_339), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_377), .B(n_336), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_378), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_379), .B(n_336), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_377), .B(n_348), .Y(n_422) );
AOI21xp33_ASAP7_75t_L g423 ( .A1(n_362), .A2(n_353), .B(n_343), .Y(n_423) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_370), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_378), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_372), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_372), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_383), .B(n_345), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_368), .B(n_345), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_388), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_379), .B(n_345), .Y(n_431) );
INVx1_ASAP7_75t_SL g432 ( .A(n_364), .Y(n_432) );
INVxp67_ASAP7_75t_SL g433 ( .A(n_363), .Y(n_433) );
NOR3xp33_ASAP7_75t_L g434 ( .A(n_385), .B(n_328), .C(n_355), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_382), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_382), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_430), .B(n_380), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_392), .B(n_345), .Y(n_438) );
AOI211xp5_ASAP7_75t_L g439 ( .A1(n_423), .A2(n_359), .B(n_343), .C(n_351), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_416), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_416), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_411), .B(n_361), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_430), .B(n_361), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_406), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_411), .B(n_361), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_392), .B(n_345), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_396), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_389), .B(n_351), .Y(n_448) );
INVxp67_ASAP7_75t_L g449 ( .A(n_413), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_395), .B(n_346), .Y(n_450) );
NAND4xp25_ASAP7_75t_L g451 ( .A(n_423), .B(n_359), .C(n_298), .D(n_327), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_395), .B(n_346), .Y(n_452) );
NOR3xp33_ASAP7_75t_L g453 ( .A(n_410), .B(n_355), .C(n_346), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_406), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_396), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_389), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_413), .B(n_391), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_391), .B(n_357), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_397), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_404), .B(n_357), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_422), .B(n_355), .Y(n_461) );
HB1xp67_ASAP7_75t_SL g462 ( .A(n_424), .Y(n_462) );
NOR3xp33_ASAP7_75t_L g463 ( .A(n_410), .B(n_290), .C(n_273), .Y(n_463) );
NAND4xp25_ASAP7_75t_SL g464 ( .A(n_424), .B(n_340), .C(n_357), .D(n_344), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_401), .B(n_344), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_393), .B(n_344), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_397), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_422), .B(n_344), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_402), .Y(n_469) );
NAND2x1_ASAP7_75t_SL g470 ( .A(n_404), .B(n_340), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_415), .Y(n_471) );
NAND2x1p5_ASAP7_75t_L g472 ( .A(n_406), .B(n_344), .Y(n_472) );
NAND3xp33_ASAP7_75t_L g473 ( .A(n_426), .B(n_299), .C(n_290), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_402), .Y(n_474) );
NOR2xp67_ASAP7_75t_SL g475 ( .A(n_406), .B(n_340), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_415), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_426), .B(n_8), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_393), .B(n_9), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_394), .B(n_10), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_414), .B(n_11), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_401), .B(n_271), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_408), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_408), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_394), .B(n_271), .Y(n_484) );
NOR2x1_ASAP7_75t_L g485 ( .A(n_421), .B(n_340), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_398), .B(n_271), .Y(n_486) );
AOI21xp5_ASAP7_75t_SL g487 ( .A1(n_433), .A2(n_299), .B(n_326), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_414), .Y(n_488) );
INVxp67_ASAP7_75t_L g489 ( .A(n_435), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_398), .B(n_280), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_402), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_405), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_398), .B(n_280), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_398), .B(n_280), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_459), .B(n_405), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_462), .A2(n_427), .B1(n_433), .B2(n_419), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_485), .A2(n_427), .B1(n_409), .B2(n_407), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_457), .B(n_407), .Y(n_498) );
OAI322xp33_ASAP7_75t_L g499 ( .A1(n_449), .A2(n_427), .A3(n_409), .B1(n_419), .B2(n_403), .C1(n_425), .C2(n_390), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_456), .B(n_429), .Y(n_500) );
OAI22xp33_ASAP7_75t_L g501 ( .A1(n_472), .A2(n_436), .B1(n_435), .B2(n_432), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_464), .A2(n_487), .B(n_439), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_437), .A2(n_429), .B1(n_434), .B2(n_428), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_476), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_476), .Y(n_505) );
INVx2_ASAP7_75t_SL g506 ( .A(n_458), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_440), .Y(n_507) );
NOR2xp33_ASAP7_75t_R g508 ( .A(n_468), .B(n_399), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_467), .B(n_403), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_438), .B(n_428), .Y(n_510) );
OAI321xp33_ASAP7_75t_L g511 ( .A1(n_451), .A2(n_436), .A3(n_431), .B1(n_390), .B2(n_425), .C(n_417), .Y(n_511) );
OAI21xp5_ASAP7_75t_SL g512 ( .A1(n_460), .A2(n_434), .B(n_431), .Y(n_512) );
INVxp67_ASAP7_75t_SL g513 ( .A(n_454), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_447), .B(n_418), .Y(n_514) );
INVxp67_ASAP7_75t_L g515 ( .A(n_441), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_460), .B(n_432), .Y(n_516) );
AOI32xp33_ASAP7_75t_L g517 ( .A1(n_477), .A2(n_400), .A3(n_418), .B1(n_417), .B2(n_412), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_471), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_455), .B(n_420), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_492), .B(n_420), .Y(n_520) );
NOR2xp67_ASAP7_75t_L g521 ( .A(n_454), .B(n_412), .Y(n_521) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_454), .A2(n_400), .B1(n_412), .B2(n_299), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_488), .Y(n_523) );
OAI21xp5_ASAP7_75t_SL g524 ( .A1(n_460), .A2(n_400), .B(n_300), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_438), .B(n_400), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_482), .Y(n_526) );
NAND3xp33_ASAP7_75t_SL g527 ( .A(n_453), .B(n_11), .C(n_12), .Y(n_527) );
OAI21xp5_ASAP7_75t_SL g528 ( .A1(n_472), .A2(n_300), .B(n_293), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_478), .B(n_12), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_483), .B(n_13), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_444), .B(n_296), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_463), .A2(n_293), .B1(n_300), .B2(n_283), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_477), .A2(n_293), .B1(n_300), .B2(n_270), .Y(n_533) );
XOR2x1_ASAP7_75t_L g534 ( .A(n_480), .B(n_13), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_448), .B(n_14), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_470), .Y(n_536) );
NAND2xp33_ASAP7_75t_L g537 ( .A(n_444), .B(n_270), .Y(n_537) );
AOI32xp33_ASAP7_75t_L g538 ( .A1(n_446), .A2(n_296), .A3(n_300), .B1(n_281), .B2(n_286), .Y(n_538) );
OAI32xp33_ASAP7_75t_L g539 ( .A1(n_442), .A2(n_282), .A3(n_283), .B1(n_286), .B2(n_292), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_446), .B(n_15), .Y(n_540) );
NAND4xp25_ASAP7_75t_L g541 ( .A(n_479), .B(n_16), .C(n_19), .D(n_20), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_465), .B(n_450), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_465), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_445), .A2(n_286), .B1(n_282), .B2(n_283), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_489), .Y(n_545) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_527), .A2(n_487), .B(n_473), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_511), .B(n_484), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_504), .Y(n_548) );
INVxp33_ASAP7_75t_L g549 ( .A(n_508), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_505), .B(n_484), .Y(n_550) );
INVx2_ASAP7_75t_SL g551 ( .A(n_506), .Y(n_551) );
OAI21xp33_ASAP7_75t_L g552 ( .A1(n_512), .A2(n_466), .B(n_443), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_525), .B(n_450), .Y(n_553) );
OAI211xp5_ASAP7_75t_L g554 ( .A1(n_528), .A2(n_461), .B(n_493), .C(n_490), .Y(n_554) );
INVx2_ASAP7_75t_SL g555 ( .A(n_542), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_518), .Y(n_556) );
AOI221xp5_ASAP7_75t_L g557 ( .A1(n_499), .A2(n_452), .B1(n_481), .B2(n_486), .C(n_490), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_500), .Y(n_558) );
NOR3xp33_ASAP7_75t_L g559 ( .A(n_541), .B(n_486), .C(n_469), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g560 ( .A(n_511), .B(n_481), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g561 ( .A1(n_496), .A2(n_452), .B1(n_475), .B2(n_493), .C(n_494), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_498), .B(n_491), .Y(n_562) );
AO22x1_ASAP7_75t_L g563 ( .A1(n_536), .A2(n_494), .B1(n_491), .B2(n_474), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_514), .B(n_474), .Y(n_564) );
NOR2xp67_ASAP7_75t_SL g565 ( .A(n_524), .B(n_469), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_545), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_519), .Y(n_567) );
AOI222xp33_ASAP7_75t_SL g568 ( .A1(n_496), .A2(n_19), .B1(n_22), .B2(n_23), .C1(n_292), .C2(n_286), .Y(n_568) );
AND2x4_ASAP7_75t_L g569 ( .A(n_516), .B(n_22), .Y(n_569) );
XNOR2x1_ASAP7_75t_L g570 ( .A(n_534), .B(n_296), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_509), .B(n_277), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_507), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_520), .Y(n_573) );
XOR2xp5_ASAP7_75t_L g574 ( .A(n_503), .B(n_25), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_497), .A2(n_292), .B1(n_282), .B2(n_285), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_523), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_540), .Y(n_577) );
AO22x2_ASAP7_75t_L g578 ( .A1(n_513), .A2(n_292), .B1(n_30), .B2(n_31), .Y(n_578) );
NOR2xp67_ASAP7_75t_L g579 ( .A(n_502), .B(n_29), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_526), .Y(n_580) );
AO21x1_ASAP7_75t_L g581 ( .A1(n_549), .A2(n_501), .B(n_537), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_564), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_559), .A2(n_529), .B1(n_543), .B2(n_532), .Y(n_583) );
NOR2x1_ASAP7_75t_SL g584 ( .A(n_554), .B(n_544), .Y(n_584) );
AOI322xp5_ASAP7_75t_L g585 ( .A1(n_557), .A2(n_510), .A3(n_536), .B1(n_530), .B2(n_495), .C1(n_515), .C2(n_533), .Y(n_585) );
NAND3xp33_ASAP7_75t_SL g586 ( .A(n_568), .B(n_517), .C(n_522), .Y(n_586) );
OAI221xp5_ASAP7_75t_L g587 ( .A1(n_561), .A2(n_535), .B1(n_538), .B2(n_521), .C(n_544), .Y(n_587) );
NOR3x1_ASAP7_75t_L g588 ( .A(n_560), .B(n_531), .C(n_539), .Y(n_588) );
NAND2xp33_ASAP7_75t_SL g589 ( .A(n_565), .B(n_34), .Y(n_589) );
A2O1A1Ixp33_ASAP7_75t_L g590 ( .A1(n_561), .A2(n_281), .B(n_277), .C(n_285), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_550), .B(n_277), .Y(n_591) );
AOI31xp33_ASAP7_75t_L g592 ( .A1(n_570), .A2(n_36), .A3(n_38), .B(n_42), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_547), .A2(n_285), .B1(n_281), .B2(n_182), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_548), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_567), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_546), .A2(n_209), .B1(n_49), .B2(n_52), .C(n_53), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_552), .A2(n_209), .B1(n_54), .B2(n_56), .C(n_57), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_550), .Y(n_598) );
OAI21xp33_ASAP7_75t_L g599 ( .A1(n_546), .A2(n_278), .B(n_60), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g600 ( .A1(n_569), .A2(n_46), .B(n_61), .C(n_65), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_573), .A2(n_278), .B(n_68), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_585), .B(n_566), .Y(n_602) );
AOI211x1_ASAP7_75t_SL g603 ( .A1(n_586), .A2(n_579), .B(n_568), .C(n_571), .Y(n_603) );
INVx2_ASAP7_75t_SL g604 ( .A(n_582), .Y(n_604) );
AOI31xp33_ASAP7_75t_L g605 ( .A1(n_581), .A2(n_569), .A3(n_574), .B(n_551), .Y(n_605) );
BUFx2_ASAP7_75t_L g606 ( .A(n_589), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_592), .B(n_575), .Y(n_607) );
NAND3xp33_ASAP7_75t_L g608 ( .A(n_587), .B(n_563), .C(n_556), .Y(n_608) );
XNOR2x1_ASAP7_75t_L g609 ( .A(n_584), .B(n_578), .Y(n_609) );
OAI21xp33_ASAP7_75t_L g610 ( .A1(n_587), .A2(n_571), .B(n_576), .Y(n_610) );
OAI211xp5_ASAP7_75t_L g611 ( .A1(n_583), .A2(n_577), .B(n_572), .C(n_558), .Y(n_611) );
AOI222xp33_ASAP7_75t_L g612 ( .A1(n_595), .A2(n_580), .B1(n_555), .B2(n_578), .C1(n_553), .C2(n_562), .Y(n_612) );
AOI211xp5_ASAP7_75t_L g613 ( .A1(n_590), .A2(n_66), .B(n_71), .C(n_73), .Y(n_613) );
NAND3xp33_ASAP7_75t_SL g614 ( .A(n_603), .B(n_596), .C(n_600), .Y(n_614) );
NAND4xp75_ASAP7_75t_L g615 ( .A(n_602), .B(n_588), .C(n_596), .D(n_597), .Y(n_615) );
AO22x2_ASAP7_75t_L g616 ( .A1(n_609), .A2(n_594), .B1(n_598), .B2(n_591), .Y(n_616) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_605), .B(n_599), .C(n_601), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_604), .B(n_608), .Y(n_618) );
OAI322xp33_ASAP7_75t_SL g619 ( .A1(n_605), .A2(n_593), .A3(n_75), .B1(n_78), .B2(n_79), .C1(n_80), .C2(n_81), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_618), .B(n_606), .Y(n_620) );
OA22x2_ASAP7_75t_L g621 ( .A1(n_616), .A2(n_610), .B1(n_611), .B2(n_607), .Y(n_621) );
A2O1A1Ixp33_ASAP7_75t_L g622 ( .A1(n_614), .A2(n_617), .B(n_615), .C(n_619), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_618), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_623), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_620), .Y(n_625) );
OAI221xp5_ASAP7_75t_L g626 ( .A1(n_625), .A2(n_622), .B1(n_621), .B2(n_612), .C(n_613), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_625), .Y(n_627) );
NAND4xp25_ASAP7_75t_L g628 ( .A(n_626), .B(n_624), .C(n_620), .D(n_84), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_628), .A2(n_627), .B1(n_182), .B2(n_209), .Y(n_629) );
OR2x6_ASAP7_75t_L g630 ( .A(n_629), .B(n_278), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_630), .A2(n_182), .B1(n_82), .B2(n_85), .Y(n_631) );
endmodule