module fake_ariane_498_n_667 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_667);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_667;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_226;
wire n_220;
wire n_261;
wire n_663;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_665;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_566;
wire n_578;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_661;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_616;
wire n_658;
wire n_617;
wire n_630;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_147;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;

INVx1_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_81),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_134),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_86),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_13),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_9),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_72),
.Y(n_153)
);

BUFx2_ASAP7_75t_SL g154 ( 
.A(n_136),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_89),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_15),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_41),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_117),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_12),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_56),
.Y(n_161)
);

BUFx2_ASAP7_75t_SL g162 ( 
.A(n_39),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_130),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_48),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_49),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_58),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_113),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_63),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_43),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_84),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_52),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_124),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_51),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_87),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_80),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_7),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_17),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_91),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_92),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_78),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_17),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_36),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_7),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_69),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_98),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_82),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_114),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_108),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_33),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_60),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_115),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_76),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_101),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_25),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_75),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_70),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_27),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_55),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_61),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_137),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_32),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_35),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_102),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_133),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_140),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_13),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_111),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_109),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_31),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_28),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_119),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_151),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_145),
.B(n_0),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_199),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_152),
.Y(n_222)
);

INVxp67_ASAP7_75t_SL g223 ( 
.A(n_193),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_169),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_160),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_169),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_159),
.B(n_0),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_180),
.B(n_1),
.Y(n_228)
);

NOR2xp67_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_1),
.Y(n_229)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_161),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g231 ( 
.A(n_161),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_181),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_183),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_191),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_196),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_146),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_147),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g242 ( 
.A(n_207),
.Y(n_242)
);

INVxp33_ASAP7_75t_SL g243 ( 
.A(n_213),
.Y(n_243)
);

NOR2xp67_ASAP7_75t_L g244 ( 
.A(n_165),
.B(n_2),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_198),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_202),
.B(n_2),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_149),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_153),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_209),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_165),
.B(n_3),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_155),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_213),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_157),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_158),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_163),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_257),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_215),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_221),
.B(n_166),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_148),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_166),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_171),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_222),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_217),
.B(n_225),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_233),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_244),
.B(n_164),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_223),
.B(n_167),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_257),
.B(n_154),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_222),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_240),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_259),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_233),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_241),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_235),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_253),
.B(n_210),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_235),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_219),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_250),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_251),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_219),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_243),
.B(n_168),
.Y(n_291)
);

BUFx8_ASAP7_75t_L g292 ( 
.A(n_232),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_255),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_234),
.B(n_162),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_254),
.Y(n_295)
);

AND2x6_ASAP7_75t_L g296 ( 
.A(n_238),
.B(n_150),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_260),
.B(n_170),
.Y(n_297)
);

AOI22x1_ASAP7_75t_SL g298 ( 
.A1(n_214),
.A2(n_206),
.B1(n_205),
.B2(n_204),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_239),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_248),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_245),
.B(n_172),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_214),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_230),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_220),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_231),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_259),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_255),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_220),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_236),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_228),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_237),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_237),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_271),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_264),
.B(n_216),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_242),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_271),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_247),
.Y(n_320)
);

INVx6_ASAP7_75t_L g321 ( 
.A(n_292),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_276),
.A2(n_227),
.B1(n_218),
.B2(n_229),
.Y(n_322)
);

INVx4_ASAP7_75t_SL g323 ( 
.A(n_296),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_262),
.Y(n_324)
);

INVx6_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

AND2x6_ASAP7_75t_L g326 ( 
.A(n_270),
.B(n_150),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_279),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_283),
.B(n_173),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_300),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_300),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_150),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_313),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_271),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_284),
.A2(n_286),
.B1(n_265),
.B2(n_268),
.Y(n_335)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_300),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_272),
.Y(n_337)
);

BUFx8_ASAP7_75t_SL g338 ( 
.A(n_313),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_300),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_272),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_311),
.B(n_174),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_150),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_L g344 ( 
.A1(n_267),
.A2(n_203),
.B1(n_200),
.B2(n_197),
.Y(n_344)
);

BUFx4f_ASAP7_75t_L g345 ( 
.A(n_294),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_284),
.A2(n_195),
.B1(n_194),
.B2(n_192),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_272),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_288),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_265),
.B(n_286),
.Y(n_349)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_289),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_295),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_301),
.Y(n_352)
);

NAND2x1p5_ASAP7_75t_L g353 ( 
.A(n_290),
.B(n_175),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_303),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_178),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_290),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_272),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_308),
.B(n_3),
.Y(n_359)
);

NAND3x1_ASAP7_75t_L g360 ( 
.A(n_291),
.B(n_263),
.C(n_266),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_274),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_282),
.B(n_179),
.Y(n_362)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_296),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_278),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_281),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_292),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_282),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_282),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_302),
.B(n_182),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_312),
.B(n_269),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_275),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_296),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_296),
.Y(n_373)
);

INVxp33_ASAP7_75t_L g374 ( 
.A(n_277),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_307),
.B(n_4),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_261),
.A2(n_280),
.B1(n_285),
.B2(n_273),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_285),
.B(n_184),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_297),
.B(n_185),
.Y(n_378)
);

INVx6_ASAP7_75t_L g379 ( 
.A(n_296),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_261),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_273),
.B(n_188),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_315),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_189),
.Y(n_383)
);

A2O1A1Ixp33_ASAP7_75t_L g384 ( 
.A1(n_322),
.A2(n_280),
.B(n_190),
.C(n_309),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_345),
.B(n_350),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_361),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_327),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_378),
.B(n_296),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_4),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_342),
.B(n_5),
.Y(n_391)
);

NAND3xp33_ASAP7_75t_L g392 ( 
.A(n_342),
.B(n_298),
.C(n_305),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_320),
.B(n_5),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_349),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_320),
.B(n_6),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_355),
.Y(n_396)
);

NAND3xp33_ASAP7_75t_L g397 ( 
.A(n_344),
.B(n_305),
.C(n_303),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_361),
.Y(n_398)
);

AND2x2_ASAP7_75t_SL g399 ( 
.A(n_322),
.B(n_6),
.Y(n_399)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_379),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_368),
.B(n_8),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_345),
.B(n_8),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_364),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_343),
.B(n_9),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_344),
.B(n_377),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_343),
.B(n_10),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_L g407 ( 
.A1(n_324),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_341),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_360),
.B(n_11),
.Y(n_409)
);

OR2x2_ASAP7_75t_SL g410 ( 
.A(n_333),
.B(n_14),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_352),
.B(n_14),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_364),
.B(n_365),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_364),
.B(n_15),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_354),
.B(n_16),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_L g415 ( 
.A(n_348),
.B(n_21),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_365),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_365),
.B(n_16),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_367),
.B(n_18),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_316),
.B(n_18),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_329),
.B(n_356),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_328),
.B(n_19),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_314),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_377),
.B(n_19),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_326),
.B(n_20),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_326),
.B(n_20),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_326),
.B(n_144),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_314),
.B(n_22),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_376),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_326),
.B(n_29),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_353),
.B(n_143),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_366),
.B(n_30),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_L g433 ( 
.A1(n_376),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_314),
.B(n_40),
.Y(n_434)
);

NAND3xp33_ASAP7_75t_L g435 ( 
.A(n_351),
.B(n_42),
.C(n_44),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_349),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_317),
.Y(n_437)
);

OAI22xp33_ASAP7_75t_L g438 ( 
.A1(n_359),
.A2(n_353),
.B1(n_381),
.B2(n_332),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_330),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_381),
.B(n_142),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_336),
.B(n_318),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_321),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_336),
.B(n_45),
.Y(n_443)
);

OR2x6_ASAP7_75t_L g444 ( 
.A(n_321),
.B(n_46),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_318),
.B(n_47),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_363),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_446)
);

A2O1A1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_332),
.A2(n_57),
.B(n_59),
.C(n_62),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_319),
.B(n_139),
.Y(n_448)
);

NAND2x1p5_ASAP7_75t_L g449 ( 
.A(n_400),
.B(n_363),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_388),
.B(n_380),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_405),
.B(n_369),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_405),
.B(n_394),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_399),
.B(n_325),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_408),
.Y(n_454)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_444),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_319),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_394),
.B(n_362),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_382),
.B(n_374),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_388),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_382),
.B(n_325),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_R g461 ( 
.A(n_442),
.B(n_370),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_396),
.B(n_362),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_421),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_400),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_399),
.A2(n_339),
.B1(n_331),
.B2(n_346),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_439),
.Y(n_466)
);

INVx5_ASAP7_75t_L g467 ( 
.A(n_444),
.Y(n_467)
);

AO22x1_ASAP7_75t_L g468 ( 
.A1(n_432),
.A2(n_338),
.B1(n_375),
.B2(n_373),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_432),
.B(n_373),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_422),
.Y(n_470)
);

AOI211xp5_ASAP7_75t_L g471 ( 
.A1(n_397),
.A2(n_334),
.B(n_337),
.C(n_347),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_423),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_411),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_419),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_390),
.A2(n_346),
.B1(n_340),
.B2(n_357),
.Y(n_475)
);

INVx5_ASAP7_75t_L g476 ( 
.A(n_444),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_418),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_437),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_384),
.B(n_335),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_420),
.B(n_340),
.Y(n_480)
);

NAND2x1p5_ASAP7_75t_L g481 ( 
.A(n_386),
.B(n_373),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_393),
.B(n_335),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_395),
.B(n_357),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_385),
.A2(n_403),
.B1(n_398),
.B2(n_416),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_386),
.B(n_357),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_438),
.B(n_372),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_438),
.B(n_372),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_410),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_409),
.Y(n_489)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_423),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_414),
.B(n_379),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_387),
.B(n_323),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_452),
.A2(n_389),
.B(n_440),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_457),
.A2(n_391),
.B(n_424),
.Y(n_494)
);

OAI21x1_ASAP7_75t_SL g495 ( 
.A1(n_451),
.A2(n_429),
.B(n_433),
.Y(n_495)
);

OA21x2_ASAP7_75t_L g496 ( 
.A1(n_486),
.A2(n_448),
.B(n_445),
.Y(n_496)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_483),
.A2(n_443),
.B(n_412),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_458),
.B(n_383),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_462),
.A2(n_401),
.B(n_441),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_453),
.B(n_402),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_456),
.A2(n_431),
.B(n_402),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_492),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_453),
.B(n_415),
.Y(n_503)
);

A2O1A1Ixp33_ASAP7_75t_L g504 ( 
.A1(n_482),
.A2(n_433),
.B(n_429),
.C(n_407),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_454),
.B(n_455),
.Y(n_505)
);

AO31x2_ASAP7_75t_L g506 ( 
.A1(n_477),
.A2(n_413),
.A3(n_417),
.B(n_406),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_465),
.B(n_425),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_456),
.A2(n_404),
.B(n_426),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_455),
.B(n_407),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_455),
.B(n_392),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_450),
.Y(n_511)
);

OA21x2_ASAP7_75t_L g512 ( 
.A1(n_487),
.A2(n_428),
.B(n_434),
.Y(n_512)
);

A2O1A1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_473),
.A2(n_446),
.B(n_435),
.C(n_447),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_450),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_463),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_492),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_474),
.B(n_434),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_467),
.B(n_428),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_481),
.A2(n_430),
.B(n_427),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_464),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_461),
.Y(n_521)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_481),
.A2(n_485),
.B(n_484),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_466),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_516),
.B(n_479),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_504),
.A2(n_498),
.B1(n_500),
.B2(n_517),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_497),
.A2(n_475),
.B(n_446),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_495),
.A2(n_467),
.B1(n_476),
.B2(n_470),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_523),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_515),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_504),
.A2(n_475),
.B(n_480),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_519),
.A2(n_472),
.B(n_449),
.Y(n_531)
);

A2O1A1Ixp33_ASAP7_75t_L g532 ( 
.A1(n_517),
.A2(n_465),
.B(n_471),
.C(n_489),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_506),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_512),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_506),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_519),
.A2(n_472),
.B(n_449),
.Y(n_536)
);

O2A1O1Ixp33_ASAP7_75t_SL g537 ( 
.A1(n_513),
.A2(n_471),
.B(n_464),
.C(n_490),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_SL g538 ( 
.A1(n_509),
.A2(n_476),
.B1(n_467),
.B2(n_469),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_516),
.B(n_476),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_502),
.Y(n_540)
);

AO21x2_ASAP7_75t_L g541 ( 
.A1(n_507),
.A2(n_460),
.B(n_469),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_513),
.A2(n_490),
.B(n_469),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_493),
.A2(n_490),
.B(n_469),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_502),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_507),
.A2(n_488),
.B1(n_478),
.B2(n_459),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_521),
.A2(n_478),
.B1(n_491),
.B2(n_468),
.Y(n_546)
);

A2O1A1Ixp33_ASAP7_75t_L g547 ( 
.A1(n_518),
.A2(n_323),
.B(n_65),
.C(n_66),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_514),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_514),
.B(n_323),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_L g550 ( 
.A1(n_505),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_548),
.B(n_511),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_524),
.A2(n_510),
.B1(n_503),
.B2(n_518),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_540),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_548),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_540),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_528),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_528),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_529),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_543),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_540),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_524),
.B(n_502),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_SL g562 ( 
.A(n_532),
.B(n_494),
.C(n_499),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_529),
.B(n_506),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_525),
.B(n_527),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_534),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_545),
.A2(n_520),
.B1(n_502),
.B2(n_501),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_540),
.Y(n_567)
);

OAI221xp5_ASAP7_75t_L g568 ( 
.A1(n_530),
.A2(n_508),
.B1(n_512),
.B2(n_520),
.C(n_496),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_544),
.B(n_522),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_546),
.B(n_71),
.Y(n_570)
);

AOI21xp33_ASAP7_75t_L g571 ( 
.A1(n_530),
.A2(n_512),
.B(n_496),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_539),
.B(n_506),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_526),
.A2(n_496),
.B(n_74),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_541),
.A2(n_138),
.B1(n_77),
.B2(n_83),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_533),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_542),
.A2(n_73),
.B(n_85),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_538),
.A2(n_88),
.B1(n_90),
.B2(n_94),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_542),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_578)
);

AND2x2_ASAP7_75t_SL g579 ( 
.A(n_540),
.B(n_99),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_540),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_541),
.Y(n_581)
);

NAND2x1p5_ASAP7_75t_L g582 ( 
.A(n_579),
.B(n_544),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_569),
.B(n_541),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_554),
.B(n_539),
.Y(n_584)
);

OAI221xp5_ASAP7_75t_L g585 ( 
.A1(n_570),
.A2(n_552),
.B1(n_564),
.B2(n_574),
.C(n_562),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_554),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_556),
.B(n_533),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_579),
.A2(n_535),
.B1(n_550),
.B2(n_534),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_563),
.B(n_535),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_569),
.B(n_544),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_579),
.A2(n_561),
.B1(n_566),
.B2(n_578),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_558),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_576),
.A2(n_537),
.B(n_543),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_557),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_551),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_561),
.B(n_544),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_563),
.A2(n_534),
.B1(n_526),
.B2(n_549),
.Y(n_597)
);

AOI33xp33_ASAP7_75t_L g598 ( 
.A1(n_574),
.A2(n_547),
.A3(n_103),
.B1(n_104),
.B2(n_105),
.B3(n_106),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_568),
.A2(n_536),
.B(n_531),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_SL g600 ( 
.A1(n_581),
.A2(n_536),
.B1(n_531),
.B2(n_116),
.Y(n_600)
);

AOI221xp5_ASAP7_75t_L g601 ( 
.A1(n_571),
.A2(n_100),
.B1(n_107),
.B2(n_118),
.C(n_120),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_561),
.B(n_121),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_555),
.Y(n_603)
);

INVx6_ASAP7_75t_L g604 ( 
.A(n_553),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_586),
.B(n_572),
.Y(n_605)
);

OR2x2_ASAP7_75t_SL g606 ( 
.A(n_595),
.B(n_580),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_586),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_584),
.B(n_555),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_594),
.B(n_575),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_592),
.B(n_575),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_590),
.B(n_567),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_587),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_590),
.B(n_567),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_589),
.B(n_581),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_590),
.B(n_560),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_596),
.B(n_560),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_583),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_583),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_583),
.Y(n_619)
);

BUFx10_ASAP7_75t_L g620 ( 
.A(n_607),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_609),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_609),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_614),
.B(n_589),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_605),
.B(n_603),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_611),
.B(n_603),
.Y(n_625)
);

AOI322xp5_ASAP7_75t_L g626 ( 
.A1(n_614),
.A2(n_588),
.A3(n_591),
.B1(n_585),
.B2(n_601),
.C1(n_600),
.C2(n_598),
.Y(n_626)
);

OAI211xp5_ASAP7_75t_L g627 ( 
.A1(n_610),
.A2(n_588),
.B(n_593),
.C(n_599),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_623),
.B(n_612),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_621),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_625),
.B(n_613),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_622),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_624),
.B(n_605),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_620),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_620),
.B(n_615),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_629),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_633),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_634),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_629),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_630),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_636),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_636),
.B(n_620),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_635),
.Y(n_642)
);

OAI32xp33_ASAP7_75t_L g643 ( 
.A1(n_638),
.A2(n_632),
.A3(n_631),
.B1(n_628),
.B2(n_582),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_639),
.Y(n_644)
);

AOI222xp33_ASAP7_75t_L g645 ( 
.A1(n_640),
.A2(n_627),
.B1(n_626),
.B2(n_610),
.C1(n_637),
.C2(n_608),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_640),
.A2(n_627),
.B1(n_606),
.B2(n_582),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_642),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_645),
.A2(n_641),
.B1(n_644),
.B2(n_602),
.Y(n_648)
);

OAI211xp5_ASAP7_75t_L g649 ( 
.A1(n_647),
.A2(n_641),
.B(n_643),
.C(n_577),
.Y(n_649)
);

AOI21xp33_ASAP7_75t_L g650 ( 
.A1(n_649),
.A2(n_646),
.B(n_569),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_650),
.B(n_648),
.Y(n_651)
);

NOR3xp33_ASAP7_75t_L g652 ( 
.A(n_651),
.B(n_598),
.C(n_553),
.Y(n_652)
);

NAND3xp33_ASAP7_75t_L g653 ( 
.A(n_652),
.B(n_580),
.C(n_553),
.Y(n_653)
);

XNOR2x1_ASAP7_75t_L g654 ( 
.A(n_653),
.B(n_122),
.Y(n_654)
);

NOR4xp25_ASAP7_75t_L g655 ( 
.A(n_654),
.B(n_616),
.C(n_559),
.D(n_597),
.Y(n_655)
);

BUFx4f_ASAP7_75t_SL g656 ( 
.A(n_655),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_656),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_657),
.A2(n_573),
.B(n_559),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_658),
.Y(n_659)
);

XOR2xp5_ASAP7_75t_L g660 ( 
.A(n_659),
.B(n_123),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_659),
.A2(n_573),
.B(n_127),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_660),
.A2(n_580),
.B1(n_604),
.B2(n_559),
.Y(n_662)
);

OR2x6_ASAP7_75t_L g663 ( 
.A(n_661),
.B(n_580),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_SL g664 ( 
.A1(n_663),
.A2(n_580),
.B1(n_128),
.B2(n_129),
.Y(n_664)
);

AOI222xp33_ASAP7_75t_L g665 ( 
.A1(n_662),
.A2(n_619),
.B1(n_618),
.B2(n_617),
.C1(n_135),
.C2(n_125),
.Y(n_665)
);

OAI221xp5_ASAP7_75t_R g666 ( 
.A1(n_664),
.A2(n_131),
.B1(n_132),
.B2(n_604),
.C(n_597),
.Y(n_666)
);

AOI211xp5_ASAP7_75t_L g667 ( 
.A1(n_666),
.A2(n_665),
.B(n_604),
.C(n_565),
.Y(n_667)
);


endmodule