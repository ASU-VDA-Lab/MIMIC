module fake_jpeg_32135_n_81 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_81);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_81;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_27),
.B(n_32),
.C(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_3),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_27),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_28),
.C(n_30),
.Y(n_41)
);

A2O1A1O1Ixp25_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_50),
.B(n_27),
.C(n_29),
.D(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_6),
.B1(n_10),
.B2(n_12),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_26),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_59),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_SL g60 ( 
.A(n_54),
.B(n_13),
.C(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_25),
.B1(n_7),
.B2(n_9),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_44),
.B1(n_49),
.B2(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_61),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g61 ( 
.A(n_58),
.B(n_48),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_67),
.Y(n_71)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_16),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_23),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_65),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_72),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_75),
.B(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_77),
.B(n_70),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_61),
.B1(n_69),
.B2(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);


endmodule