module real_jpeg_6013_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g129 ( 
.A(n_0),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_1),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_1),
.A2(n_81),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_1),
.A2(n_81),
.B1(n_309),
.B2(n_311),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_1),
.A2(n_81),
.B1(n_291),
.B2(n_296),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_2),
.A2(n_55),
.B1(n_59),
.B2(n_62),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_2),
.A2(n_62),
.B1(n_166),
.B2(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_4),
.A2(n_68),
.B1(n_72),
.B2(n_73),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_4),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_4),
.A2(n_72),
.B1(n_231),
.B2(n_233),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_5),
.A2(n_38),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_5),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_5),
.A2(n_133),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_5),
.A2(n_133),
.B1(n_291),
.B2(n_296),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_5),
.A2(n_133),
.B1(n_349),
.B2(n_351),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_6),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_6),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_7),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_7),
.Y(n_237)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_8),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_9),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_9),
.Y(n_265)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_9),
.Y(n_322)
);

INVx8_ASAP7_75t_L g337 ( 
.A(n_9),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_10),
.A2(n_42),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_10),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_10),
.A2(n_94),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_10),
.A2(n_94),
.B1(n_166),
.B2(n_190),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_10),
.A2(n_94),
.B1(n_300),
.B2(n_304),
.Y(n_299)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_13),
.A2(n_41),
.B1(n_192),
.B2(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_13),
.B(n_286),
.C(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_13),
.B(n_122),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_13),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_13),
.B(n_174),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_13),
.B(n_364),
.Y(n_363)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_14),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_14),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_14),
.Y(n_97)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_15),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_15),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_16),
.A2(n_166),
.B1(n_169),
.B2(n_172),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_16),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_16),
.A2(n_172),
.B1(n_214),
.B2(n_218),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_16),
.A2(n_172),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_245),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_244),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_204),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_21),
.B(n_204),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_141),
.C(n_186),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_22),
.B(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_75),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_23),
.B(n_76),
.C(n_105),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_44),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_24),
.A2(n_44),
.B1(n_45),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_24),
.Y(n_254)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.A3(n_33),
.B1(n_35),
.B2(n_40),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_29),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_30),
.Y(n_135)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_39),
.Y(n_201)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_39),
.Y(n_361)
);

OAI21xp33_ASAP7_75t_SL g195 ( 
.A1(n_40),
.A2(n_41),
.B(n_42),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_41),
.B(n_85),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_41),
.A2(n_46),
.B(n_298),
.Y(n_323)
);

OAI21xp33_ASAP7_75t_SL g358 ( 
.A1(n_41),
.A2(n_359),
.B(n_362),
.Y(n_358)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_53),
.B1(n_63),
.B2(n_66),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_46),
.A2(n_63),
.B1(n_180),
.B2(n_236),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_46),
.A2(n_290),
.B(n_298),
.Y(n_289)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_47),
.A2(n_67),
.B1(n_179),
.B2(n_184),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_47),
.A2(n_54),
.B1(n_259),
.B2(n_263),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_47),
.B(n_299),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_47),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_52),
.Y(n_162)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_52),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_52),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_52),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_52),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_57),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_58),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_58),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_60),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.Y(n_158)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_61),
.Y(n_261)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_64),
.B(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_104),
.B2(n_105),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_83),
.B(n_92),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_78),
.A2(n_85),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_82),
.Y(n_223)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_84),
.B(n_93),
.Y(n_197)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_89),
.Y(n_219)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.Y(n_92)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_97),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_98),
.A2(n_195),
.B(n_196),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_98),
.Y(n_221)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_131),
.B(n_136),
.Y(n_105)
);

AOI22x1_ASAP7_75t_L g210 ( 
.A1(n_106),
.A2(n_122),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_106),
.B(n_211),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_106),
.A2(n_136),
.B(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_107),
.A2(n_132),
.B1(n_140),
.B2(n_199),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_122),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_112),
.B1(n_116),
.B2(n_121),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_110),
.Y(n_376)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_111),
.Y(n_381)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_115),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_115),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

AO22x2_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_130),
.Y(n_122)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_126),
.Y(n_234)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_128),
.Y(n_350)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_129),
.Y(n_232)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_129),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_130),
.Y(n_279)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx6_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_137),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_140),
.A2(n_199),
.B(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_141),
.A2(n_142),
.B1(n_186),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_178),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_143),
.B(n_178),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_165),
.B1(n_173),
.B2(n_175),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_144),
.A2(n_277),
.B(n_280),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_144),
.A2(n_173),
.B1(n_308),
.B2(n_348),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_144),
.A2(n_280),
.B(n_348),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_145),
.A2(n_174),
.B1(n_176),
.B2(n_230),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_158),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_150),
.B1(n_153),
.B2(n_156),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_149),
.Y(n_284)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_149),
.Y(n_310)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_157),
.Y(n_312)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_158),
.A2(n_188),
.B(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_160),
.Y(n_286)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_165),
.A2(n_173),
.B(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_171),
.Y(n_373)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_174),
.B(n_189),
.Y(n_280)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_186),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.C(n_198),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_187),
.B(n_198),
.Y(n_250)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_193),
.A2(n_194),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_228),
.B1(n_242),
.B2(n_243),
.Y(n_206)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_220),
.B1(n_226),
.B2(n_227),
.Y(n_209)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_215),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI32xp33_ASAP7_75t_L g371 ( 
.A1(n_218),
.A2(n_363),
.A3(n_372),
.B1(n_374),
.B2(n_377),
.Y(n_371)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_220),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_235),
.Y(n_228)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_241),
.Y(n_297)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_241),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_270),
.B(n_400),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_267),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_248),
.B(n_267),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.C(n_255),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_249),
.B(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_255),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.C(n_266),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_256),
.B(n_391),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_258),
.B(n_266),
.Y(n_391)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_259),
.Y(n_368)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_265),
.Y(n_370)
);

AOI21x1_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_394),
.B(n_399),
.Y(n_270)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_383),
.B(n_393),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_342),
.B(n_382),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_315),
.B(n_341),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_288),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_275),
.B(n_288),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_276),
.A2(n_281),
.B1(n_282),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_276),
.Y(n_339)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_305),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_289),
.B(n_306),
.C(n_314),
.Y(n_343)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_290),
.Y(n_334)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_295),
.Y(n_303)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_296),
.Y(n_319)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_313),
.B2(n_314),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_309),
.Y(n_378)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_331),
.B(n_340),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_324),
.B(n_330),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_323),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_322),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_329),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_327),
.B(n_328),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_326),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_328),
.A2(n_368),
.B(n_369),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_338),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_338),
.Y(n_340)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_343),
.B(n_344),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_366),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_356),
.B2(n_357),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_347),
.B(n_356),
.C(n_366),
.Y(n_384)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx5_ASAP7_75t_SL g352 ( 
.A(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVxp33_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx6_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_371),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_371),
.Y(n_389)
);

INVx3_ASAP7_75t_SL g369 ( 
.A(n_370),
.Y(n_369)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NAND2xp33_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_384),
.B(n_385),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_387),
.B1(n_390),
.B2(n_392),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_389),
.C(n_392),
.Y(n_395)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_390),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_395),
.B(n_396),
.Y(n_399)
);


endmodule