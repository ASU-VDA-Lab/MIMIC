module fake_jpeg_20230_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

AOI21xp33_ASAP7_75t_L g7 ( 
.A1(n_0),
.A2(n_2),
.B(n_4),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_4),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_0),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

AND2x4_ASAP7_75t_SL g15 ( 
.A(n_7),
.B(n_12),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_15),
.A2(n_9),
.B(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_16),
.B(n_10),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_6),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_17),
.A2(n_7),
.B1(n_9),
.B2(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

AO21x2_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_12),
.B(n_10),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_21),
.B1(n_15),
.B2(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_16),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_15),
.C(n_19),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_25),
.B(n_21),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_27),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_15),
.C(n_18),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_27),
.A2(n_21),
.B1(n_14),
.B2(n_11),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_11),
.B1(n_3),
.B2(n_5),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_21),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_32),
.B(n_28),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_33),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_3),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_30),
.B(n_5),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_33),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_36),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_37),
.Y(n_39)
);


endmodule