module fake_jpeg_26550_n_154 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_154);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_1),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_29),
.C(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_34),
.Y(n_47)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_1),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_1),
.C(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_30),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_3),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_41),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_19),
.Y(n_62)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_65),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_20),
.B1(n_17),
.B2(n_25),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_17),
.B(n_20),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_24),
.C(n_15),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_16),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_25),
.B1(n_27),
.B2(n_15),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_27),
.B1(n_24),
.B2(n_14),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_19),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_23),
.Y(n_65)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_23),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_69),
.Y(n_80)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_70),
.B(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

OR2x2_ASAP7_75t_SL g92 ( 
.A(n_73),
.B(n_81),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g102 ( 
.A(n_75),
.B(n_84),
.C(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_14),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_56),
.C(n_59),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_63),
.C(n_18),
.Y(n_105)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_19),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_41),
.B1(n_33),
.B2(n_38),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_89),
.Y(n_94)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_45),
.B1(n_42),
.B2(n_35),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_13),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_3),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_45),
.B1(n_18),
.B2(n_35),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_67),
.B(n_66),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_104),
.Y(n_110)
);

AO22x1_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_55),
.B1(n_69),
.B2(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_101),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_57),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_99),
.B(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_4),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_107),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_106),
.A2(n_104),
.B1(n_97),
.B2(n_94),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_63),
.C(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_5),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_84),
.B(n_98),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_79),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_78),
.C(n_72),
.Y(n_128)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_95),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_117),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_83),
.B(n_73),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_116),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_84),
.B1(n_74),
.B2(n_55),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_74),
.B1(n_81),
.B2(n_89),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_122),
.B(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_111),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_133),
.Y(n_141)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_101),
.B(n_108),
.C(n_92),
.D(n_105),
.Y(n_126)
);

XNOR2x1_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_130),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_129),
.C(n_131),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_72),
.C(n_86),
.Y(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_5),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_10),
.C(n_7),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_9),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_138),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_116),
.B1(n_119),
.B2(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_112),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_139),
.B(n_141),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_126),
.C(n_10),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_137),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_145),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_147),
.A2(n_135),
.B(n_144),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_150),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_10),
.B(n_139),
.C(n_143),
.D(n_145),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_148),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_153),
.Y(n_154)
);


endmodule