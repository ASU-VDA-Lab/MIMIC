module fake_jpeg_52_n_226 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_226);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx11_ASAP7_75t_SL g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_1),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_14),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_82),
.Y(n_87)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_84),
.B(n_76),
.C(n_58),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_84),
.B(n_86),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_86),
.A2(n_77),
.B1(n_60),
.B2(n_75),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_88),
.A2(n_95),
.B1(n_97),
.B2(n_83),
.Y(n_113)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_55),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_74),
.Y(n_115)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_55),
.B1(n_66),
.B2(n_59),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_83),
.B1(n_56),
.B2(n_63),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_77),
.B1(n_60),
.B2(n_75),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_60),
.B1(n_76),
.B2(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_102),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_67),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_54),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_105),
.B(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_69),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_61),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_116),
.B1(n_58),
.B2(n_51),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_83),
.B1(n_74),
.B2(n_72),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_114),
.A2(n_71),
.B1(n_57),
.B2(n_96),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_117),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_63),
.B1(n_71),
.B2(n_56),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_73),
.C(n_65),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_68),
.Y(n_125)
);

AOI22x1_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_96),
.B1(n_68),
.B2(n_53),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_140),
.Y(n_148)
);

CKINVDCx12_ASAP7_75t_R g121 ( 
.A(n_117),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_121),
.B(n_127),
.Y(n_153)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_126),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_0),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_0),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_58),
.B1(n_2),
.B2(n_3),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_130),
.A2(n_119),
.B1(n_7),
.B2(n_9),
.Y(n_144)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_101),
.B(n_1),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_133),
.Y(n_145)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_135),
.B(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_102),
.B(n_5),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_109),
.B(n_112),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_24),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_164),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_25),
.B1(n_48),
.B2(n_45),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_162),
.B1(n_160),
.B2(n_157),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_122),
.A2(n_6),
.B(n_9),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_157),
.B(n_14),
.Y(n_168)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_152),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_23),
.C(n_44),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_161),
.C(n_165),
.Y(n_178)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_155),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_123),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_50),
.B(n_43),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_6),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_158),
.B(n_13),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_10),
.B(n_11),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_40),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_137),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_39),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_168),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_15),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_171),
.A2(n_176),
.B(n_182),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_15),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_175),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_16),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_28),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_183),
.C(n_185),
.Y(n_187)
);

OAI321xp33_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_31),
.A3(n_35),
.B1(n_34),
.B2(n_32),
.C(n_38),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_16),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_184),
.A2(n_186),
.B1(n_144),
.B2(n_162),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_18),
.C(n_19),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_147),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_196),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_172),
.A2(n_164),
.B(n_146),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_172),
.B(n_180),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_147),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_180),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_200),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_183),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_207),
.C(n_205),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_167),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_202),
.B(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_206),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_169),
.B1(n_165),
.B2(n_178),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_178),
.C(n_177),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_212),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_194),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_187),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_200),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_215),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_209),
.A2(n_198),
.B1(n_199),
.B2(n_189),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_210),
.B1(n_211),
.B2(n_193),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_SL g220 ( 
.A1(n_219),
.A2(n_216),
.B(n_214),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_218),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_185),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_222),
.Y(n_223)
);

OAI31xp33_ASAP7_75t_SL g224 ( 
.A1(n_223),
.A2(n_18),
.A3(n_19),
.B(n_20),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_21),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_21),
.Y(n_226)
);


endmodule