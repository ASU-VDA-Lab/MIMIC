module real_aes_8719_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_722, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_722;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g465 ( .A1(n_0), .A2(n_203), .B(n_466), .C(n_469), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_1), .B(n_460), .Y(n_470) );
INVx1_ASAP7_75t_L g116 ( .A(n_2), .Y(n_116) );
INVx1_ASAP7_75t_L g238 ( .A(n_3), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_4), .B(n_155), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_5), .A2(n_455), .B(n_543), .Y(n_542) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_6), .A2(n_178), .B(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_7), .A2(n_38), .B1(n_148), .B2(n_172), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_8), .B(n_178), .Y(n_250) );
AND2x6_ASAP7_75t_L g163 ( .A(n_9), .B(n_164), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_10), .A2(n_163), .B(n_446), .C(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_11), .B(n_39), .Y(n_117) );
INVx1_ASAP7_75t_L g144 ( .A(n_12), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_13), .B(n_153), .Y(n_186) );
INVx1_ASAP7_75t_L g230 ( .A(n_14), .Y(n_230) );
OAI22xp5_ASAP7_75t_SL g711 ( .A1(n_15), .A2(n_76), .B1(n_712), .B2(n_713), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_15), .Y(n_713) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_16), .B(n_155), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_17), .B(n_179), .Y(n_217) );
AO32x2_ASAP7_75t_L g200 ( .A1(n_18), .A2(n_177), .A3(n_178), .B1(n_201), .B2(n_205), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_19), .B(n_148), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_20), .B(n_179), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_21), .A2(n_55), .B1(n_148), .B2(n_172), .Y(n_204) );
AOI22xp33_ASAP7_75t_SL g175 ( .A1(n_22), .A2(n_83), .B1(n_148), .B2(n_153), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_23), .B(n_148), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_24), .A2(n_177), .B(n_446), .C(n_493), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_25), .A2(n_177), .B(n_446), .C(n_508), .Y(n_507) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_26), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_27), .B(n_140), .Y(n_259) );
OAI22xp5_ASAP7_75t_SL g700 ( .A1(n_28), .A2(n_94), .B1(n_701), .B2(n_702), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_28), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_29), .A2(n_699), .B1(n_700), .B2(n_703), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_29), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_30), .A2(n_455), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_31), .B(n_140), .Y(n_165) );
INVx2_ASAP7_75t_L g150 ( .A(n_32), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_33), .A2(n_452), .B(n_478), .C(n_479), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_34), .B(n_148), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_35), .B(n_140), .Y(n_193) );
OAI22xp5_ASAP7_75t_SL g716 ( .A1(n_36), .A2(n_43), .B1(n_436), .B2(n_717), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_36), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_37), .B(n_188), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_40), .B(n_491), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_41), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_42), .B(n_155), .Y(n_531) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_43), .A2(n_131), .B1(n_436), .B2(n_437), .Y(n_130) );
INVx1_ASAP7_75t_L g436 ( .A(n_43), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_44), .B(n_455), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_45), .A2(n_452), .B(n_478), .C(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_46), .B(n_148), .Y(n_245) );
INVx1_ASAP7_75t_L g467 ( .A(n_47), .Y(n_467) );
AOI22xp5_ASAP7_75t_SL g127 ( .A1(n_48), .A2(n_114), .B1(n_128), .B2(n_706), .Y(n_127) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_49), .A2(n_92), .B1(n_172), .B2(n_173), .Y(n_171) );
INVx1_ASAP7_75t_L g530 ( .A(n_50), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_51), .B(n_148), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_52), .B(n_148), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_53), .B(n_455), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_54), .B(n_236), .Y(n_249) );
AOI22xp33_ASAP7_75t_SL g221 ( .A1(n_56), .A2(n_60), .B1(n_148), .B2(n_153), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_57), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_58), .B(n_148), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_59), .B(n_148), .Y(n_258) );
INVx1_ASAP7_75t_L g164 ( .A(n_61), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_62), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_63), .B(n_460), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_64), .A2(n_233), .B(n_236), .C(n_546), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_65), .A2(n_105), .B1(n_118), .B2(n_719), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_66), .B(n_148), .Y(n_239) );
INVx1_ASAP7_75t_L g143 ( .A(n_67), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_68), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_69), .B(n_155), .Y(n_483) );
AO32x2_ASAP7_75t_L g169 ( .A1(n_70), .A2(n_170), .A3(n_176), .B1(n_177), .B2(n_178), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_71), .B(n_156), .Y(n_520) );
INVx1_ASAP7_75t_L g257 ( .A(n_72), .Y(n_257) );
INVx1_ASAP7_75t_L g151 ( .A(n_73), .Y(n_151) );
CKINVDCx16_ASAP7_75t_R g463 ( .A(n_74), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_75), .B(n_482), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_76), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_L g445 ( .A1(n_77), .A2(n_446), .B(n_448), .C(n_452), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_78), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_79), .B(n_153), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g544 ( .A(n_80), .Y(n_544) );
INVx1_ASAP7_75t_L g110 ( .A(n_81), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_82), .B(n_481), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_84), .B(n_172), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_85), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_86), .B(n_153), .Y(n_160) );
INVx2_ASAP7_75t_L g141 ( .A(n_87), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_88), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_89), .B(n_174), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_90), .B(n_153), .Y(n_246) );
INVx2_ASAP7_75t_L g113 ( .A(n_91), .Y(n_113) );
OR2x2_ASAP7_75t_L g125 ( .A(n_91), .B(n_114), .Y(n_125) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_93), .A2(n_103), .B1(n_153), .B2(n_154), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_94), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_95), .B(n_455), .Y(n_476) );
INVx1_ASAP7_75t_L g480 ( .A(n_96), .Y(n_480) );
INVxp67_ASAP7_75t_L g547 ( .A(n_97), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_98), .B(n_153), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_99), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g449 ( .A(n_100), .Y(n_449) );
INVx1_ASAP7_75t_L g516 ( .A(n_101), .Y(n_516) );
AND2x2_ASAP7_75t_L g532 ( .A(n_102), .B(n_140), .Y(n_532) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx12_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g720 ( .A(n_108), .Y(n_720) );
OR2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
INVx1_ASAP7_75t_SL g706 ( .A(n_111), .Y(n_706) );
INVx3_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
NOR2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AO22x2_ASAP7_75t_SL g129 ( .A1(n_113), .A2(n_130), .B1(n_438), .B2(n_697), .Y(n_129) );
INVx1_ASAP7_75t_L g697 ( .A(n_113), .Y(n_697) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
AOI22x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_127), .B1(n_707), .B2(n_708), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_123), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_SL g707 ( .A(n_121), .Y(n_707) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_123), .A2(n_709), .B(n_718), .Y(n_708) );
NOR2xp33_ASAP7_75t_SL g123 ( .A(n_124), .B(n_126), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx2_ASAP7_75t_L g718 ( .A(n_125), .Y(n_718) );
OAI22xp33_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_698), .B1(n_704), .B2(n_705), .Y(n_128) );
INVx1_ASAP7_75t_L g704 ( .A(n_129), .Y(n_704) );
INVx1_ASAP7_75t_L g437 ( .A(n_131), .Y(n_437) );
OAI22xp5_ASAP7_75t_SL g714 ( .A1(n_131), .A2(n_437), .B1(n_715), .B2(n_716), .Y(n_714) );
OR2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_357), .Y(n_131) );
NAND3xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_306), .C(n_348), .Y(n_132) );
AOI211xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_211), .B(n_260), .C(n_282), .Y(n_133) );
OAI211xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_166), .B(n_194), .C(n_206), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_136), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g369 ( .A(n_136), .B(n_286), .Y(n_369) );
BUFx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g271 ( .A(n_137), .B(n_197), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_137), .B(n_182), .Y(n_388) );
INVx1_ASAP7_75t_L g406 ( .A(n_137), .Y(n_406) );
AND2x2_ASAP7_75t_L g415 ( .A(n_137), .B(n_303), .Y(n_415) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g298 ( .A(n_138), .B(n_182), .Y(n_298) );
AND2x2_ASAP7_75t_L g356 ( .A(n_138), .B(n_303), .Y(n_356) );
INVx1_ASAP7_75t_L g400 ( .A(n_138), .Y(n_400) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g277 ( .A(n_139), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g285 ( .A(n_139), .Y(n_285) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_139), .Y(n_325) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_145), .B(n_165), .Y(n_139) );
INVx2_ASAP7_75t_L g176 ( .A(n_140), .Y(n_176) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_140), .A2(n_183), .B(n_193), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_140), .A2(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g499 ( .A(n_140), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_140), .A2(n_527), .B(n_528), .Y(n_526) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_L g179 ( .A(n_141), .B(n_142), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
OAI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_158), .B(n_163), .Y(n_145) );
O2A1O1Ixp5_ASAP7_75t_SL g146 ( .A1(n_147), .A2(n_151), .B(n_152), .C(n_155), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_148), .Y(n_451) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g172 ( .A(n_149), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
AND2x6_ASAP7_75t_L g446 ( .A(n_149), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g154 ( .A(n_150), .Y(n_154) );
INVx1_ASAP7_75t_L g237 ( .A(n_150), .Y(n_237) );
INVx2_ASAP7_75t_L g231 ( .A(n_153), .Y(n_231) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g203 ( .A(n_155), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_155), .A2(n_245), .B(n_246), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_155), .A2(n_254), .B(n_255), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_155), .B(n_547), .Y(n_546) );
INVx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OAI22xp5_ASAP7_75t_SL g170 ( .A1(n_156), .A2(n_171), .B1(n_174), .B2(n_175), .Y(n_170) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_157), .Y(n_162) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_157), .Y(n_174) );
INVx1_ASAP7_75t_L g188 ( .A(n_157), .Y(n_188) );
INVx1_ASAP7_75t_L g447 ( .A(n_157), .Y(n_447) );
AND2x2_ASAP7_75t_L g456 ( .A(n_157), .B(n_237), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_161), .Y(n_158) );
INVx1_ASAP7_75t_L g233 ( .A(n_161), .Y(n_233) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g482 ( .A(n_162), .Y(n_482) );
BUFx3_ASAP7_75t_L g177 ( .A(n_163), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_163), .A2(n_184), .B(n_189), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_163), .A2(n_229), .B(n_234), .Y(n_228) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_163), .A2(n_244), .B(n_247), .Y(n_243) );
INVx4_ASAP7_75t_SL g453 ( .A(n_163), .Y(n_453) );
AND2x4_ASAP7_75t_L g455 ( .A(n_163), .B(n_456), .Y(n_455) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_163), .B(n_456), .Y(n_517) );
INVxp67_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_180), .Y(n_167) );
AND2x2_ASAP7_75t_L g264 ( .A(n_168), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g297 ( .A(n_168), .Y(n_297) );
OR2x2_ASAP7_75t_L g423 ( .A(n_168), .B(n_424), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_168), .B(n_182), .Y(n_427) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g197 ( .A(n_169), .Y(n_197) );
INVx1_ASAP7_75t_L g209 ( .A(n_169), .Y(n_209) );
AND2x2_ASAP7_75t_L g286 ( .A(n_169), .B(n_199), .Y(n_286) );
AND2x2_ASAP7_75t_L g326 ( .A(n_169), .B(n_200), .Y(n_326) );
INVx2_ASAP7_75t_L g469 ( .A(n_173), .Y(n_469) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_173), .Y(n_484) );
INVx2_ASAP7_75t_L g192 ( .A(n_174), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_174), .A2(n_202), .B1(n_203), .B2(n_204), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_174), .A2(n_203), .B1(n_220), .B2(n_221), .Y(n_219) );
INVx4_ASAP7_75t_L g468 ( .A(n_174), .Y(n_468) );
INVx1_ASAP7_75t_L g496 ( .A(n_176), .Y(n_496) );
NAND3xp33_ASAP7_75t_L g218 ( .A(n_177), .B(n_219), .C(n_222), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_177), .A2(n_253), .B(n_256), .Y(n_252) );
INVx4_ASAP7_75t_L g222 ( .A(n_178), .Y(n_222) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_178), .A2(n_243), .B(n_250), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_178), .A2(n_506), .B(n_507), .Y(n_505) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_178), .Y(n_541) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g205 ( .A(n_179), .Y(n_205) );
INVxp67_ASAP7_75t_L g368 ( .A(n_180), .Y(n_368) );
AND2x4_ASAP7_75t_L g393 ( .A(n_180), .B(n_286), .Y(n_393) );
BUFx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_SL g284 ( .A(n_181), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g198 ( .A(n_182), .B(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g272 ( .A(n_182), .B(n_200), .Y(n_272) );
INVx1_ASAP7_75t_L g278 ( .A(n_182), .Y(n_278) );
INVx2_ASAP7_75t_L g304 ( .A(n_182), .Y(n_304) );
AND2x2_ASAP7_75t_L g320 ( .A(n_182), .B(n_321), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .Y(n_184) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_192), .Y(n_189) );
O2A1O1Ixp5_ASAP7_75t_L g256 ( .A1(n_192), .A2(n_235), .B(n_257), .C(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_195), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_198), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
BUFx2_ASAP7_75t_L g275 ( .A(n_197), .Y(n_275) );
AND2x2_ASAP7_75t_L g383 ( .A(n_197), .B(n_199), .Y(n_383) );
AND2x2_ASAP7_75t_L g300 ( .A(n_198), .B(n_285), .Y(n_300) );
AND2x2_ASAP7_75t_L g399 ( .A(n_198), .B(n_400), .Y(n_399) );
NOR2xp67_ASAP7_75t_L g321 ( .A(n_199), .B(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g424 ( .A(n_199), .B(n_285), .Y(n_424) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
BUFx2_ASAP7_75t_L g210 ( .A(n_200), .Y(n_210) );
AND2x2_ASAP7_75t_L g303 ( .A(n_200), .B(n_304), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_203), .A2(n_235), .B(n_238), .C(n_239), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_203), .A2(n_248), .B(n_249), .Y(n_247) );
INVx2_ASAP7_75t_L g227 ( .A(n_205), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_205), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_210), .Y(n_207) );
AND2x2_ASAP7_75t_L g349 ( .A(n_208), .B(n_284), .Y(n_349) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_209), .B(n_285), .Y(n_334) );
INVx2_ASAP7_75t_L g333 ( .A(n_210), .Y(n_333) );
OAI222xp33_ASAP7_75t_L g337 ( .A1(n_210), .A2(n_277), .B1(n_338), .B2(n_340), .C1(n_341), .C2(n_344), .Y(n_337) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_223), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g262 ( .A(n_215), .Y(n_262) );
OR2x2_ASAP7_75t_L g373 ( .A(n_215), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx3_ASAP7_75t_L g295 ( .A(n_216), .Y(n_295) );
NOR2x1_ASAP7_75t_L g346 ( .A(n_216), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g352 ( .A(n_216), .B(n_266), .Y(n_352) );
AND2x4_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
INVx1_ASAP7_75t_L g313 ( .A(n_217), .Y(n_313) );
AO21x1_ASAP7_75t_L g312 ( .A1(n_219), .A2(n_222), .B(n_313), .Y(n_312) );
AO21x2_ASAP7_75t_L g443 ( .A1(n_222), .A2(n_444), .B(n_457), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_222), .B(n_458), .Y(n_457) );
INVx3_ASAP7_75t_L g460 ( .A(n_222), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_222), .B(n_486), .Y(n_485) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_222), .A2(n_515), .B(n_522), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_223), .A2(n_316), .B1(n_355), .B2(n_356), .Y(n_354) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_241), .Y(n_223) );
INVx3_ASAP7_75t_L g288 ( .A(n_224), .Y(n_288) );
OR2x2_ASAP7_75t_L g421 ( .A(n_224), .B(n_297), .Y(n_421) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g294 ( .A(n_225), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g310 ( .A(n_225), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g318 ( .A(n_225), .B(n_266), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_225), .B(n_242), .Y(n_374) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g265 ( .A(n_226), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g269 ( .A(n_226), .B(n_242), .Y(n_269) );
AND2x2_ASAP7_75t_L g345 ( .A(n_226), .B(n_292), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_226), .B(n_251), .Y(n_385) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_240), .Y(n_226) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_227), .A2(n_252), .B(n_259), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_232), .C(n_233), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_231), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_231), .A2(n_520), .B(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_L g448 ( .A1(n_233), .A2(n_449), .B(n_450), .C(n_451), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_235), .A2(n_494), .B(n_495), .Y(n_493) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_241), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g301 ( .A(n_241), .B(n_262), .Y(n_301) );
AND2x2_ASAP7_75t_L g305 ( .A(n_241), .B(n_295), .Y(n_305) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_251), .Y(n_241) );
INVx3_ASAP7_75t_L g266 ( .A(n_242), .Y(n_266) );
AND2x2_ASAP7_75t_L g291 ( .A(n_242), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g426 ( .A(n_242), .B(n_409), .Y(n_426) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_251), .Y(n_280) );
INVx2_ASAP7_75t_L g292 ( .A(n_251), .Y(n_292) );
AND2x2_ASAP7_75t_L g336 ( .A(n_251), .B(n_312), .Y(n_336) );
INVx1_ASAP7_75t_L g379 ( .A(n_251), .Y(n_379) );
OR2x2_ASAP7_75t_L g410 ( .A(n_251), .B(n_312), .Y(n_410) );
AND2x2_ASAP7_75t_L g430 ( .A(n_251), .B(n_266), .Y(n_430) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_263), .B(n_267), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g268 ( .A(n_262), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_262), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g387 ( .A(n_264), .Y(n_387) );
INVx2_ASAP7_75t_SL g281 ( .A(n_265), .Y(n_281) );
AND2x2_ASAP7_75t_L g401 ( .A(n_265), .B(n_295), .Y(n_401) );
INVx2_ASAP7_75t_L g347 ( .A(n_266), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_266), .B(n_379), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_270), .B1(n_273), .B2(n_279), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_269), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g435 ( .A(n_269), .Y(n_435) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g360 ( .A(n_271), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_271), .B(n_303), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_272), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g376 ( .A(n_272), .B(n_325), .Y(n_376) );
INVx2_ASAP7_75t_L g432 ( .A(n_272), .Y(n_432) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x2_ASAP7_75t_L g302 ( .A(n_275), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_275), .B(n_320), .Y(n_353) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_277), .B(n_297), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g414 ( .A(n_280), .Y(n_414) );
O2A1O1Ixp33_ASAP7_75t_SL g364 ( .A1(n_281), .A2(n_365), .B(n_367), .C(n_370), .Y(n_364) );
OR2x2_ASAP7_75t_L g391 ( .A(n_281), .B(n_295), .Y(n_391) );
OAI221xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_287), .B1(n_289), .B2(n_296), .C(n_299), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_284), .B(n_286), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_284), .B(n_333), .Y(n_340) );
AND2x2_ASAP7_75t_L g382 ( .A(n_284), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g418 ( .A(n_284), .Y(n_418) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_285), .Y(n_309) );
INVx1_ASAP7_75t_L g322 ( .A(n_285), .Y(n_322) );
NOR2xp67_ASAP7_75t_L g342 ( .A(n_288), .B(n_343), .Y(n_342) );
INVxp67_ASAP7_75t_L g396 ( .A(n_288), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_288), .B(n_336), .Y(n_412) );
INVx2_ASAP7_75t_L g398 ( .A(n_289), .Y(n_398) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g339 ( .A(n_291), .B(n_310), .Y(n_339) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_291), .A2(n_307), .B(n_349), .C(n_350), .Y(n_348) );
AND2x2_ASAP7_75t_L g317 ( .A(n_292), .B(n_312), .Y(n_317) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_296), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
OR2x2_ASAP7_75t_L g365 ( .A(n_297), .B(n_366), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B1(n_302), .B2(n_305), .Y(n_299) );
INVx1_ASAP7_75t_L g419 ( .A(n_301), .Y(n_419) );
INVx1_ASAP7_75t_L g366 ( .A(n_303), .Y(n_366) );
INVx1_ASAP7_75t_L g417 ( .A(n_305), .Y(n_417) );
AOI211xp5_ASAP7_75t_SL g306 ( .A1(n_307), .A2(n_310), .B(n_314), .C(n_337), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g329 ( .A(n_309), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g380 ( .A(n_310), .Y(n_380) );
AND2x2_ASAP7_75t_L g429 ( .A(n_310), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OAI21xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_319), .B(n_327), .Y(n_314) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx2_ASAP7_75t_L g343 ( .A(n_317), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_317), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g335 ( .A(n_318), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g411 ( .A(n_318), .Y(n_411) );
OAI32xp33_ASAP7_75t_L g422 ( .A1(n_318), .A2(n_370), .A3(n_377), .B1(n_418), .B2(n_423), .Y(n_422) );
NOR2xp33_ASAP7_75t_SL g319 ( .A(n_320), .B(n_323), .Y(n_319) );
INVx1_ASAP7_75t_SL g390 ( .A(n_320), .Y(n_390) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g330 ( .A(n_326), .Y(n_330) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_331), .B(n_335), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI22xp33_ASAP7_75t_L g402 ( .A1(n_329), .A2(n_377), .B1(n_403), .B2(n_405), .Y(n_402) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_333), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g370 ( .A(n_336), .Y(n_370) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g363 ( .A(n_347), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_353), .B(n_354), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_356), .A2(n_398), .B1(n_399), .B2(n_401), .C(n_402), .Y(n_397) );
NAND5xp2_ASAP7_75t_L g357 ( .A(n_358), .B(n_381), .C(n_397), .D(n_407), .E(n_425), .Y(n_357) );
AOI211xp5_ASAP7_75t_SL g358 ( .A1(n_359), .A2(n_361), .B(n_364), .C(n_371), .Y(n_358) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g428 ( .A(n_365), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
OAI22xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B1(n_375), .B2(n_377), .Y(n_371) );
INVx1_ASAP7_75t_SL g404 ( .A(n_374), .Y(n_404) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI322xp33_ASAP7_75t_L g386 ( .A1(n_377), .A2(n_387), .A3(n_388), .B1(n_389), .B2(n_390), .C1(n_391), .C2(n_392), .Y(n_386) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx1_ASAP7_75t_L g389 ( .A(n_379), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_379), .B(n_404), .Y(n_403) );
AOI211xp5_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_384), .B(n_386), .C(n_394), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_390), .A2(n_417), .B1(n_418), .B2(n_419), .Y(n_416) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g433 ( .A(n_400), .Y(n_433) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_415), .B1(n_416), .B2(n_420), .C(n_422), .Y(n_407) );
OAI211xp5_ASAP7_75t_SL g408 ( .A1(n_409), .A2(n_411), .B(n_412), .C(n_413), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g434 ( .A(n_410), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B1(n_428), .B2(n_429), .C(n_431), .Y(n_425) );
AOI21xp33_ASAP7_75t_SL g431 ( .A1(n_432), .A2(n_433), .B(n_434), .Y(n_431) );
NAND2x1p5_ASAP7_75t_L g438 ( .A(n_439), .B(n_640), .Y(n_438) );
AND4x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_580), .C(n_595), .D(n_620), .Y(n_439) );
NOR2xp33_ASAP7_75t_SL g440 ( .A(n_441), .B(n_553), .Y(n_440) );
OAI21xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_471), .B(n_533), .Y(n_441) );
AND2x2_ASAP7_75t_L g583 ( .A(n_442), .B(n_488), .Y(n_583) );
AND2x2_ASAP7_75t_L g596 ( .A(n_442), .B(n_487), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_442), .B(n_472), .Y(n_646) );
INVx1_ASAP7_75t_L g650 ( .A(n_442), .Y(n_650) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_459), .Y(n_442) );
INVx2_ASAP7_75t_L g567 ( .A(n_443), .Y(n_567) );
BUFx2_ASAP7_75t_L g594 ( .A(n_443), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_454), .Y(n_444) );
INVx5_ASAP7_75t_L g464 ( .A(n_446), .Y(n_464) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_SL g462 ( .A1(n_453), .A2(n_463), .B(n_464), .C(n_465), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_453), .A2(n_464), .B(n_544), .C(n_545), .Y(n_543) );
BUFx2_ASAP7_75t_L g491 ( .A(n_455), .Y(n_491) );
AND2x2_ASAP7_75t_L g534 ( .A(n_459), .B(n_488), .Y(n_534) );
INVx2_ASAP7_75t_L g550 ( .A(n_459), .Y(n_550) );
AND2x2_ASAP7_75t_L g559 ( .A(n_459), .B(n_487), .Y(n_559) );
AND2x2_ASAP7_75t_L g638 ( .A(n_459), .B(n_567), .Y(n_638) );
OA21x2_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B(n_470), .Y(n_459) );
INVx2_ASAP7_75t_L g478 ( .A(n_464), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_500), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_472), .B(n_565), .Y(n_603) );
INVx1_ASAP7_75t_L g691 ( .A(n_472), .Y(n_691) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_487), .Y(n_472) );
AND2x2_ASAP7_75t_L g549 ( .A(n_473), .B(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g563 ( .A(n_473), .B(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_473), .Y(n_592) );
OR2x2_ASAP7_75t_L g624 ( .A(n_473), .B(n_566), .Y(n_624) );
AND2x2_ASAP7_75t_L g632 ( .A(n_473), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g665 ( .A(n_473), .B(n_634), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_473), .B(n_534), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_473), .B(n_594), .Y(n_690) );
AND2x2_ASAP7_75t_L g696 ( .A(n_473), .B(n_583), .Y(n_696) );
INVx5_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g556 ( .A(n_474), .Y(n_556) );
AND2x2_ASAP7_75t_L g586 ( .A(n_474), .B(n_566), .Y(n_586) );
AND2x2_ASAP7_75t_L g619 ( .A(n_474), .B(n_579), .Y(n_619) );
AND2x2_ASAP7_75t_L g639 ( .A(n_474), .B(n_488), .Y(n_639) );
AND2x2_ASAP7_75t_L g673 ( .A(n_474), .B(n_539), .Y(n_673) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_485), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B(n_483), .C(n_484), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_481), .A2(n_484), .B(n_530), .C(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x4_ASAP7_75t_L g579 ( .A(n_487), .B(n_550), .Y(n_579) );
AND2x2_ASAP7_75t_L g590 ( .A(n_487), .B(n_586), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_487), .B(n_566), .Y(n_629) );
INVx2_ASAP7_75t_L g644 ( .A(n_487), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_487), .B(n_578), .Y(n_667) );
AND2x2_ASAP7_75t_L g686 ( .A(n_487), .B(n_638), .Y(n_686) );
INVx5_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_488), .Y(n_585) );
AND2x2_ASAP7_75t_L g593 ( .A(n_488), .B(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g634 ( .A(n_488), .B(n_550), .Y(n_634) );
OR2x6_ASAP7_75t_L g488 ( .A(n_489), .B(n_497), .Y(n_488) );
AOI21xp5_ASAP7_75t_SL g489 ( .A1(n_490), .A2(n_492), .B(n_496), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_511), .Y(n_501) );
AND2x2_ASAP7_75t_L g557 ( .A(n_502), .B(n_540), .Y(n_557) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_503), .B(n_514), .Y(n_537) );
OR2x2_ASAP7_75t_L g570 ( .A(n_503), .B(n_540), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_503), .B(n_540), .Y(n_575) );
AND2x2_ASAP7_75t_L g602 ( .A(n_503), .B(n_539), .Y(n_602) );
AND2x2_ASAP7_75t_L g654 ( .A(n_503), .B(n_513), .Y(n_654) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_504), .B(n_524), .Y(n_562) );
AND2x2_ASAP7_75t_L g598 ( .A(n_504), .B(n_514), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_511), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OR2x2_ASAP7_75t_L g588 ( .A(n_512), .B(n_570), .Y(n_588) );
OR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_524), .Y(n_512) );
OAI322xp33_ASAP7_75t_L g553 ( .A1(n_513), .A2(n_554), .A3(n_558), .B1(n_560), .B2(n_563), .C1(n_568), .C2(n_576), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_513), .B(n_539), .Y(n_561) );
OR2x2_ASAP7_75t_L g571 ( .A(n_513), .B(n_525), .Y(n_571) );
AND2x2_ASAP7_75t_L g573 ( .A(n_513), .B(n_525), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_513), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_513), .B(n_540), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_513), .B(n_669), .Y(n_668) );
INVx5_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_514), .B(n_557), .Y(n_683) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_518), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_524), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g551 ( .A(n_524), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_524), .B(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g613 ( .A(n_524), .B(n_540), .Y(n_613) );
AOI211xp5_ASAP7_75t_SL g641 ( .A1(n_524), .A2(n_642), .B(n_645), .C(n_657), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_524), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g679 ( .A(n_524), .B(n_654), .Y(n_679) );
INVx5_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g607 ( .A(n_525), .B(n_540), .Y(n_607) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_525), .Y(n_616) );
AND2x2_ASAP7_75t_L g656 ( .A(n_525), .B(n_654), .Y(n_656) );
AND2x2_ASAP7_75t_SL g687 ( .A(n_525), .B(n_557), .Y(n_687) );
AND2x2_ASAP7_75t_L g694 ( .A(n_525), .B(n_653), .Y(n_694) );
OR2x6_ASAP7_75t_L g525 ( .A(n_526), .B(n_532), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B1(n_549), .B2(n_551), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_534), .B(n_556), .Y(n_604) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g552 ( .A(n_537), .Y(n_552) );
OR2x2_ASAP7_75t_L g612 ( .A(n_537), .B(n_613), .Y(n_612) );
OAI221xp5_ASAP7_75t_SL g660 ( .A1(n_537), .A2(n_661), .B1(n_663), .B2(n_664), .C(n_666), .Y(n_660) );
INVx2_ASAP7_75t_L g599 ( .A(n_538), .Y(n_599) );
AND2x2_ASAP7_75t_L g572 ( .A(n_539), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g662 ( .A(n_539), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_539), .B(n_654), .Y(n_675) );
INVx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVxp67_ASAP7_75t_L g617 ( .A(n_540), .Y(n_617) );
AND2x2_ASAP7_75t_L g653 ( .A(n_540), .B(n_654), .Y(n_653) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B(n_548), .Y(n_540) );
AND2x2_ASAP7_75t_L g655 ( .A(n_549), .B(n_594), .Y(n_655) );
AND2x2_ASAP7_75t_L g565 ( .A(n_550), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_550), .B(n_623), .Y(n_622) );
NOR2xp33_ASAP7_75t_SL g636 ( .A(n_552), .B(n_599), .Y(n_636) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g642 ( .A(n_555), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
OR2x2_ASAP7_75t_L g628 ( .A(n_556), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g693 ( .A(n_556), .B(n_638), .Y(n_693) );
INVx2_ASAP7_75t_L g626 ( .A(n_557), .Y(n_626) );
NAND4xp25_ASAP7_75t_SL g689 ( .A(n_558), .B(n_690), .C(n_691), .D(n_692), .Y(n_689) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_559), .B(n_623), .Y(n_658) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_SL g695 ( .A(n_562), .Y(n_695) );
O2A1O1Ixp33_ASAP7_75t_SL g657 ( .A1(n_563), .A2(n_626), .B(n_630), .C(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g652 ( .A(n_565), .B(n_644), .Y(n_652) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_566), .Y(n_578) );
INVx1_ASAP7_75t_L g633 ( .A(n_566), .Y(n_633) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_567), .Y(n_610) );
AOI211xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_571), .B(n_572), .C(n_574), .Y(n_568) );
AND2x2_ASAP7_75t_L g589 ( .A(n_569), .B(n_573), .Y(n_589) );
OAI322xp33_ASAP7_75t_SL g627 ( .A1(n_569), .A2(n_628), .A3(n_630), .B1(n_631), .B2(n_635), .C1(n_636), .C2(n_637), .Y(n_627) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g649 ( .A(n_571), .B(n_575), .Y(n_649) );
INVx1_ASAP7_75t_L g630 ( .A(n_573), .Y(n_630) );
INVx1_ASAP7_75t_SL g648 ( .A(n_575), .Y(n_648) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AOI222xp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_587), .B1(n_589), .B2(n_590), .C1(n_591), .C2(n_722), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_582), .B(n_584), .Y(n_581) );
OAI322xp33_ASAP7_75t_L g670 ( .A1(n_582), .A2(n_644), .A3(n_649), .B1(n_671), .B2(n_672), .C1(n_674), .C2(n_675), .Y(n_670) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_583), .A2(n_597), .B1(n_621), .B2(n_625), .C(n_627), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
OAI222xp33_ASAP7_75t_L g600 ( .A1(n_588), .A2(n_601), .B1(n_603), .B2(n_604), .C1(n_605), .C2(n_608), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_590), .A2(n_597), .B1(n_667), .B2(n_668), .Y(n_666) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AOI211xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B(n_600), .C(n_611), .Y(n_595) );
O2A1O1Ixp33_ASAP7_75t_L g676 ( .A1(n_597), .A2(n_634), .B(n_677), .C(n_680), .Y(n_676) );
AND2x4_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g606 ( .A(n_598), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g669 ( .A(n_602), .Y(n_669) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_609), .B(n_634), .Y(n_663) );
BUFx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AOI21xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_614), .B(n_618), .Y(n_611) );
OAI221xp5_ASAP7_75t_SL g680 ( .A1(n_612), .A2(n_681), .B1(n_682), .B2(n_683), .C(n_684), .Y(n_680) );
INVxp33_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_616), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_623), .B(n_634), .Y(n_674) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
AND2x2_ASAP7_75t_L g685 ( .A(n_638), .B(n_644), .Y(n_685) );
AND4x1_ASAP7_75t_L g640 ( .A(n_641), .B(n_659), .C(n_676), .D(n_688), .Y(n_640) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI221xp5_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_647), .B1(n_649), .B2(n_650), .C(n_651), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_655), .B2(n_656), .Y(n_651) );
INVx1_ASAP7_75t_L g681 ( .A(n_652), .Y(n_681) );
INVx1_ASAP7_75t_SL g671 ( .A(n_656), .Y(n_671) );
NOR2xp33_ASAP7_75t_SL g659 ( .A(n_660), .B(n_670), .Y(n_659) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_672), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_679), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_694), .B1(n_695), .B2(n_696), .Y(n_688) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g705 ( .A(n_698), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
XNOR2xp5_ASAP7_75t_SL g710 ( .A(n_711), .B(n_714), .Y(n_710) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
endmodule