module real_aes_5541_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_976, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_974, n_9, n_23, n_72, n_132, n_119, n_160, n_973, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_975, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_976;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_974;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_973;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_975;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_260;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_938;
wire n_744;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_281;
wire n_962;
wire n_468;
wire n_746;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_298;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_296;
wire n_954;
wire n_702;
wire n_969;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_265;
wire n_354;
wire n_968;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_0), .A2(n_681), .B(n_683), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_1), .A2(n_128), .B1(n_376), .B2(n_377), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_2), .A2(n_129), .B1(n_490), .B2(n_492), .Y(n_489) );
INVx1_ASAP7_75t_L g621 ( .A(n_3), .Y(n_621) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_4), .Y(n_700) );
AND2x4_ASAP7_75t_L g713 ( .A(n_4), .B(n_714), .Y(n_713) );
AND2x4_ASAP7_75t_L g721 ( .A(n_4), .B(n_242), .Y(n_721) );
AOI22xp33_ASAP7_75t_SL g751 ( .A1(n_5), .A2(n_43), .B1(n_737), .B2(n_738), .Y(n_751) );
INVx1_ASAP7_75t_SL g923 ( .A(n_5), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_5), .A2(n_952), .B1(n_967), .B2(n_969), .Y(n_951) );
AOI221x1_ASAP7_75t_L g522 ( .A1(n_6), .A2(n_59), .B1(n_523), .B2(n_524), .C(n_525), .Y(n_522) );
INVx1_ASAP7_75t_L g447 ( .A(n_7), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_8), .A2(n_208), .B1(n_363), .B2(n_372), .Y(n_964) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_9), .A2(n_48), .B1(n_353), .B2(n_355), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_10), .A2(n_220), .B1(n_370), .B2(n_376), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_11), .A2(n_45), .B1(n_463), .B2(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_12), .A2(n_102), .B1(n_727), .B2(n_728), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_13), .A2(n_24), .B1(n_372), .B2(n_373), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_14), .A2(n_198), .B1(n_414), .B2(n_415), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_15), .A2(n_236), .B1(n_660), .B2(n_661), .Y(n_659) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_16), .Y(n_536) );
INVx1_ASAP7_75t_L g940 ( .A(n_17), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_18), .A2(n_89), .B1(n_338), .B2(n_344), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_19), .A2(n_78), .B1(n_363), .B2(n_384), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_20), .A2(n_71), .B1(n_369), .B2(n_372), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_21), .Y(n_539) );
INVx1_ASAP7_75t_L g601 ( .A(n_22), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_23), .A2(n_139), .B1(n_296), .B2(n_688), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_25), .A2(n_213), .B1(n_363), .B2(n_364), .Y(n_362) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_26), .A2(n_50), .B1(n_428), .B2(n_432), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_27), .A2(n_58), .B1(n_263), .B2(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_28), .B(n_461), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_29), .A2(n_152), .B1(n_412), .B2(n_461), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_30), .A2(n_94), .B1(n_733), .B2(n_735), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_31), .A2(n_75), .B1(n_520), .B2(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_32), .A2(n_247), .B1(n_404), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_33), .A2(n_63), .B1(n_423), .B2(n_512), .Y(n_630) );
INVx1_ASAP7_75t_L g274 ( .A(n_34), .Y(n_274) );
INVxp67_ASAP7_75t_L g293 ( .A(n_34), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_34), .B(n_190), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_35), .A2(n_36), .B1(n_443), .B2(n_444), .C(n_446), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_37), .A2(n_140), .B1(n_364), .B2(n_373), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_38), .A2(n_224), .B1(n_656), .B2(n_657), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_39), .A2(n_175), .B1(n_737), .B2(n_738), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_40), .A2(n_228), .B1(n_720), .B2(n_722), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_41), .A2(n_203), .B1(n_463), .B2(n_629), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_42), .A2(n_68), .B1(n_435), .B2(n_437), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_44), .B(n_269), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_46), .A2(n_226), .B1(n_381), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_47), .A2(n_114), .B1(n_727), .B2(n_728), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_49), .A2(n_144), .B1(n_463), .B2(n_464), .Y(n_462) );
INVx2_ASAP7_75t_L g698 ( .A(n_51), .Y(n_698) );
INVx1_ASAP7_75t_L g712 ( .A(n_52), .Y(n_712) );
AND2x4_ASAP7_75t_L g717 ( .A(n_52), .B(n_698), .Y(n_717) );
INVx1_ASAP7_75t_SL g734 ( .A(n_52), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_53), .A2(n_179), .B1(n_306), .B2(n_414), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_54), .A2(n_117), .B1(n_366), .B2(n_367), .Y(n_566) );
INVx1_ASAP7_75t_L g943 ( .A(n_55), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_56), .A2(n_187), .B1(n_451), .B2(n_452), .Y(n_450) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_57), .A2(n_167), .B1(n_642), .B2(n_644), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_60), .A2(n_116), .B1(n_437), .B2(n_466), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_61), .A2(n_195), .B1(n_329), .B2(n_454), .Y(n_674) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_62), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_64), .A2(n_93), .B1(n_347), .B2(n_349), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_65), .A2(n_204), .B1(n_664), .B2(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g689 ( .A(n_66), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_67), .B(n_379), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_69), .A2(n_149), .B1(n_737), .B2(n_738), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_70), .A2(n_98), .B1(n_369), .B2(n_370), .Y(n_963) );
INVx1_ASAP7_75t_L g769 ( .A(n_72), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_73), .B(n_377), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_74), .A2(n_134), .B1(n_263), .B2(n_285), .Y(n_262) );
INVx1_ASAP7_75t_SL g521 ( .A(n_76), .Y(n_521) );
NOR3xp33_ASAP7_75t_L g547 ( .A(n_76), .B(n_548), .C(n_549), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_77), .A2(n_109), .B1(n_458), .B2(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_79), .B(n_651), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_80), .A2(n_245), .B1(n_733), .B2(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g934 ( .A(n_81), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_82), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g280 ( .A(n_83), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_83), .B(n_189), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_84), .A2(n_202), .B1(n_366), .B2(n_367), .Y(n_965) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_85), .A2(n_91), .B1(n_733), .B2(n_735), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_86), .A2(n_177), .B1(n_366), .B2(n_367), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_87), .A2(n_135), .B1(n_485), .B2(n_487), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_88), .A2(n_180), .B1(n_353), .B2(n_355), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_90), .A2(n_243), .B1(n_418), .B2(n_419), .Y(n_417) );
INVx1_ASAP7_75t_L g440 ( .A(n_91), .Y(n_440) );
OAI222xp33_ASAP7_75t_L g455 ( .A1(n_91), .A2(n_456), .B1(n_462), .B2(n_465), .C1(n_973), .C2(n_974), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_91), .B(n_465), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_92), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_95), .A2(n_196), .B1(n_338), .B2(n_344), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_96), .A2(n_99), .B1(n_376), .B2(n_382), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_97), .A2(n_237), .B1(n_466), .B2(n_627), .Y(n_673) );
INVx1_ASAP7_75t_L g481 ( .A(n_100), .Y(n_481) );
AOI21xp33_ASAP7_75t_L g599 ( .A1(n_101), .A2(n_381), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g386 ( .A(n_103), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_104), .A2(n_173), .B1(n_369), .B2(n_370), .Y(n_930) );
AOI21xp33_ASAP7_75t_L g383 ( .A1(n_105), .A2(n_384), .B(n_385), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_106), .A2(n_244), .B1(n_423), .B2(n_425), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_107), .A2(n_238), .B1(n_369), .B2(n_370), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_108), .A2(n_130), .B1(n_370), .B2(n_373), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_110), .A2(n_192), .B1(n_722), .B2(n_737), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_111), .A2(n_145), .B1(n_304), .B2(n_306), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_112), .A2(n_142), .B1(n_384), .B2(n_561), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_113), .A2(n_235), .B1(n_463), .B2(n_464), .Y(n_508) );
INVxp33_ASAP7_75t_SL g774 ( .A(n_115), .Y(n_774) );
AO22x1_ASAP7_75t_L g453 ( .A1(n_118), .A2(n_121), .B1(n_423), .B2(n_454), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_119), .A2(n_178), .B1(n_372), .B2(n_373), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_120), .A2(n_206), .B1(n_427), .B2(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g619 ( .A(n_122), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_123), .A2(n_218), .B1(n_466), .B2(n_627), .Y(n_626) );
XNOR2x1_ASAP7_75t_L g634 ( .A(n_124), .B(n_635), .Y(n_634) );
XNOR2x2_ASAP7_75t_SL g690 ( .A(n_124), .B(n_635), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_125), .A2(n_138), .B1(n_366), .B2(n_367), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_126), .A2(n_158), .B1(n_638), .B2(n_639), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_127), .A2(n_156), .B1(n_710), .B2(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_131), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g684 ( .A(n_132), .Y(n_684) );
INVx1_ASAP7_75t_L g941 ( .A(n_133), .Y(n_941) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_136), .A2(n_150), .B1(n_347), .B2(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_137), .A2(n_230), .B1(n_364), .B2(n_369), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_141), .A2(n_160), .B1(n_419), .B2(n_654), .Y(n_653) );
XOR2xp5_ASAP7_75t_L g554 ( .A(n_143), .B(n_555), .Y(n_554) );
XOR2xp5_ASAP7_75t_L g574 ( .A(n_143), .B(n_555), .Y(n_574) );
INVx1_ASAP7_75t_L g772 ( .A(n_146), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_147), .A2(n_186), .B1(n_315), .B2(n_317), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_148), .A2(n_165), .B1(n_500), .B2(n_501), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_151), .A2(n_181), .B1(n_410), .B2(n_411), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_153), .A2(n_166), .B1(n_505), .B2(n_506), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_154), .A2(n_159), .B1(n_382), .B2(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_155), .A2(n_157), .B1(n_329), .B2(n_454), .Y(n_625) );
AOI21xp33_ASAP7_75t_L g645 ( .A1(n_161), .A2(n_646), .B(n_648), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_162), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g938 ( .A(n_163), .Y(n_938) );
INVx1_ASAP7_75t_L g357 ( .A(n_164), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_168), .A2(n_248), .B1(n_423), .B2(n_676), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_169), .A2(n_397), .B(n_401), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_170), .A2(n_222), .B1(n_363), .B2(n_372), .Y(n_931) );
OA22x2_ASAP7_75t_L g284 ( .A1(n_171), .A2(n_190), .B1(n_269), .B2(n_283), .Y(n_284) );
INVx1_ASAP7_75t_L g312 ( .A(n_171), .Y(n_312) );
AOI21xp5_ASAP7_75t_SL g936 ( .A1(n_172), .A2(n_379), .B(n_937), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_174), .A2(n_234), .B1(n_379), .B2(n_686), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_176), .A2(n_240), .B1(n_710), .B2(n_730), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_182), .A2(n_210), .B1(n_451), .B2(n_466), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_183), .Y(n_534) );
AND2x2_ASAP7_75t_L g525 ( .A(n_184), .B(n_501), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_185), .A2(n_212), .B1(n_329), .B2(n_334), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_188), .A2(n_209), .B1(n_381), .B2(n_382), .Y(n_380) );
INVx1_ASAP7_75t_L g276 ( .A(n_189), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_189), .B(n_310), .Y(n_326) );
OAI21xp33_ASAP7_75t_L g313 ( .A1(n_190), .A2(n_205), .B(n_294), .Y(n_313) );
INVx1_ASAP7_75t_L g718 ( .A(n_191), .Y(n_718) );
XNOR2x2_ASAP7_75t_SL g359 ( .A(n_193), .B(n_360), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_194), .A2(n_219), .B1(n_363), .B2(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_197), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g585 ( .A(n_199), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_199), .A2(n_211), .B1(n_733), .B2(n_735), .Y(n_747) );
INVx1_ASAP7_75t_L g715 ( .A(n_200), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g928 ( .A1(n_201), .A2(n_223), .B1(n_364), .B2(n_373), .Y(n_928) );
INVx1_ASAP7_75t_L g282 ( .A(n_205), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_205), .B(n_233), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_207), .B(n_381), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_214), .A2(n_215), .B1(n_510), .B2(n_512), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_216), .A2(n_953), .B1(n_954), .B2(n_966), .Y(n_952) );
CKINVDCx5p33_ASAP7_75t_R g953 ( .A(n_216), .Y(n_953) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_217), .Y(n_604) );
INVx1_ASAP7_75t_L g402 ( .A(n_221), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_225), .B(n_406), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_227), .A2(n_239), .B1(n_443), .B2(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g649 ( .A(n_229), .Y(n_649) );
INVx1_ASAP7_75t_L g608 ( .A(n_231), .Y(n_608) );
INVx1_ASAP7_75t_L g613 ( .A(n_232), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_233), .B(n_268), .Y(n_267) );
XOR2x2_ASAP7_75t_L g393 ( .A(n_240), .B(n_394), .Y(n_393) );
INVxp33_ASAP7_75t_L g768 ( .A(n_241), .Y(n_768) );
INVx1_ASAP7_75t_L g714 ( .A(n_242), .Y(n_714) );
INVx1_ASAP7_75t_L g616 ( .A(n_246), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_701), .B(n_704), .Y(n_249) );
AOI21xp33_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_577), .B(n_693), .Y(n_250) );
INVxp67_ASAP7_75t_SL g703 ( .A(n_251), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_477), .B1(n_478), .B2(n_576), .Y(n_251) );
INVx1_ASAP7_75t_L g576 ( .A(n_252), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_391), .B1(n_475), .B2(n_476), .Y(n_252) );
INVx1_ASAP7_75t_L g476 ( .A(n_253), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_358), .B1(n_387), .B2(n_390), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
BUFx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g389 ( .A(n_257), .Y(n_389) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
XOR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_357), .Y(n_259) );
NOR2x1_ASAP7_75t_L g260 ( .A(n_261), .B(n_327), .Y(n_260) );
NAND4xp25_ASAP7_75t_L g261 ( .A(n_262), .B(n_295), .C(n_303), .D(n_314), .Y(n_261) );
BUFx2_ASAP7_75t_L g415 ( .A(n_263), .Y(n_415) );
INVx2_ASAP7_75t_L g640 ( .A(n_263), .Y(n_640) );
BUFx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g494 ( .A(n_264), .Y(n_494) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_264), .Y(n_596) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_277), .Y(n_264) );
AND2x4_ASAP7_75t_L g305 ( .A(n_265), .B(n_299), .Y(n_305) );
AND2x4_ASAP7_75t_L g354 ( .A(n_265), .B(n_340), .Y(n_354) );
AND2x4_ASAP7_75t_L g366 ( .A(n_265), .B(n_340), .Y(n_366) );
AND2x4_ASAP7_75t_L g376 ( .A(n_265), .B(n_277), .Y(n_376) );
AND2x4_ASAP7_75t_L g384 ( .A(n_265), .B(n_299), .Y(n_384) );
AND2x4_ASAP7_75t_L g265 ( .A(n_266), .B(n_271), .Y(n_265) );
AND2x2_ASAP7_75t_L g287 ( .A(n_266), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g302 ( .A(n_266), .Y(n_302) );
OR2x2_ASAP7_75t_L g332 ( .A(n_266), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g342 ( .A(n_266), .B(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g266 ( .A(n_267), .B(n_270), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_268), .B(n_274), .Y(n_273) );
INVxp67_ASAP7_75t_L g310 ( .A(n_268), .Y(n_310) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp33_ASAP7_75t_L g275 ( .A(n_269), .B(n_276), .Y(n_275) );
NAND2xp33_ASAP7_75t_L g279 ( .A(n_269), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g283 ( .A(n_269), .Y(n_283) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_269), .Y(n_289) );
INVx1_ASAP7_75t_L g294 ( .A(n_269), .Y(n_294) );
NAND3xp33_ASAP7_75t_L g325 ( .A(n_270), .B(n_309), .C(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g301 ( .A(n_271), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g333 ( .A(n_272), .Y(n_333) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
AND2x2_ASAP7_75t_L g316 ( .A(n_277), .B(n_301), .Y(n_316) );
AND2x4_ASAP7_75t_L g335 ( .A(n_277), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g348 ( .A(n_277), .B(n_342), .Y(n_348) );
AND2x4_ASAP7_75t_L g363 ( .A(n_277), .B(n_342), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_277), .B(n_331), .Y(n_364) );
AND2x2_ASAP7_75t_L g381 ( .A(n_277), .B(n_301), .Y(n_381) );
AND2x2_ASAP7_75t_L g424 ( .A(n_277), .B(n_342), .Y(n_424) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_284), .Y(n_277) );
INVx1_ASAP7_75t_L g300 ( .A(n_278), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_280), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g292 ( .A1(n_282), .A2(n_293), .B(n_294), .Y(n_292) );
AND2x2_ASAP7_75t_L g291 ( .A(n_284), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g299 ( .A(n_284), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g341 ( .A(n_284), .Y(n_341) );
BUFx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx4f_ASAP7_75t_L g404 ( .A(n_286), .Y(n_404) );
INVx5_ASAP7_75t_L g459 ( .A(n_286), .Y(n_459) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_291), .Y(n_286) );
AND2x4_ASAP7_75t_L g377 ( .A(n_287), .B(n_291), .Y(n_377) );
AND2x2_ASAP7_75t_L g561 ( .A(n_287), .B(n_291), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g321 ( .A(n_289), .Y(n_321) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g410 ( .A(n_297), .Y(n_410) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx3_ASAP7_75t_L g461 ( .A(n_298), .Y(n_461) );
INVx2_ASAP7_75t_L g486 ( .A(n_298), .Y(n_486) );
BUFx8_ASAP7_75t_SL g523 ( .A(n_298), .Y(n_523) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_298), .Y(n_558) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_298), .Y(n_643) );
AND2x4_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
AND2x2_ASAP7_75t_L g379 ( .A(n_299), .B(n_301), .Y(n_379) );
AND2x4_ASAP7_75t_L g340 ( .A(n_300), .B(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g307 ( .A(n_301), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g356 ( .A(n_301), .B(n_340), .Y(n_356) );
AND2x4_ASAP7_75t_L g367 ( .A(n_301), .B(n_340), .Y(n_367) );
AND2x4_ASAP7_75t_L g382 ( .A(n_301), .B(n_308), .Y(n_382) );
BUFx2_ASAP7_75t_L g638 ( .A(n_304), .Y(n_638) );
BUFx3_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx3_ASAP7_75t_L g414 ( .A(n_305), .Y(n_414) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_305), .Y(n_443) );
INVx1_ASAP7_75t_L g491 ( .A(n_305), .Y(n_491) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_307), .Y(n_412) );
INVx3_ASAP7_75t_L g488 ( .A(n_307), .Y(n_488) );
AND2x4_ASAP7_75t_L g330 ( .A(n_308), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g351 ( .A(n_308), .B(n_342), .Y(n_351) );
AND2x4_ASAP7_75t_L g372 ( .A(n_308), .B(n_342), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_308), .B(n_331), .Y(n_373) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_313), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx2_ASAP7_75t_L g445 ( .A(n_315), .Y(n_445) );
BUFx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx3_ASAP7_75t_L g400 ( .A(n_316), .Y(n_400) );
INVx2_ASAP7_75t_L g498 ( .A(n_316), .Y(n_498) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_318), .B(n_601), .Y(n_600) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_319), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_SL g563 ( .A(n_319), .Y(n_563) );
INVx2_ASAP7_75t_L g686 ( .A(n_319), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g937 ( .A(n_319), .B(n_938), .Y(n_937) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx3_ASAP7_75t_L g408 ( .A(n_320), .Y(n_408) );
AO21x2_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B(n_325), .Y(n_320) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_322), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
NAND4xp25_ASAP7_75t_L g327 ( .A(n_328), .B(n_337), .C(n_346), .D(n_352), .Y(n_327) );
BUFx12f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx6_ASAP7_75t_L g421 ( .A(n_330), .Y(n_421) );
AND2x4_ASAP7_75t_L g345 ( .A(n_331), .B(n_340), .Y(n_345) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g336 ( .A(n_332), .Y(n_336) );
INVx1_ASAP7_75t_L g343 ( .A(n_333), .Y(n_343) );
BUFx3_ASAP7_75t_L g425 ( .A(n_334), .Y(n_425) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_335), .Y(n_454) );
BUFx3_ASAP7_75t_L g505 ( .A(n_335), .Y(n_505) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_335), .Y(n_520) );
BUFx12f_ASAP7_75t_L g658 ( .A(n_335), .Y(n_658) );
AND2x4_ASAP7_75t_L g370 ( .A(n_336), .B(n_340), .Y(n_370) );
INVx1_ASAP7_75t_L g436 ( .A(n_338), .Y(n_436) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_338), .Y(n_664) );
BUFx12f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_339), .Y(n_466) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
AND2x4_ASAP7_75t_L g369 ( .A(n_340), .B(n_342), .Y(n_369) );
BUFx3_ASAP7_75t_L g418 ( .A(n_344), .Y(n_418) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_345), .Y(n_451) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_345), .Y(n_627) );
BUFx4f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx4_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx4_ASAP7_75t_L g437 ( .A(n_350), .Y(n_437) );
INVx1_ASAP7_75t_L g512 ( .A(n_350), .Y(n_512) );
INVx2_ASAP7_75t_SL g591 ( .A(n_350), .Y(n_591) );
INVx1_ASAP7_75t_L g666 ( .A(n_350), .Y(n_666) );
INVx4_ASAP7_75t_L g676 ( .A(n_350), .Y(n_676) );
INVx8_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_353), .Y(n_660) );
BUFx12f_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx3_ASAP7_75t_L g429 ( .A(n_354), .Y(n_429) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_354), .Y(n_463) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g433 ( .A(n_356), .Y(n_433) );
BUFx5_ASAP7_75t_L g464 ( .A(n_356), .Y(n_464) );
BUFx3_ASAP7_75t_L g662 ( .A(n_356), .Y(n_662) );
INVx2_ASAP7_75t_L g390 ( .A(n_358), .Y(n_390) );
BUFx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_374), .Y(n_360) );
NAND4xp25_ASAP7_75t_L g361 ( .A(n_362), .B(n_365), .C(n_368), .D(n_371), .Y(n_361) );
NAND4xp25_ASAP7_75t_L g374 ( .A(n_375), .B(n_378), .C(n_380), .D(n_383), .Y(n_374) );
INVx2_ASAP7_75t_L g542 ( .A(n_376), .Y(n_542) );
INVx1_ASAP7_75t_L g944 ( .A(n_376), .Y(n_944) );
INVx4_ASAP7_75t_L g535 ( .A(n_377), .Y(n_535) );
INVx2_ASAP7_75t_L g935 ( .A(n_381), .Y(n_935) );
INVx2_ASAP7_75t_L g537 ( .A(n_382), .Y(n_537) );
INVx2_ASAP7_75t_L g540 ( .A(n_384), .Y(n_540) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g475 ( .A(n_391), .Y(n_475) );
AO22x2_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_393), .B1(n_438), .B2(n_474), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NOR2x1_ASAP7_75t_L g394 ( .A(n_395), .B(n_416), .Y(n_394) );
NAND3xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_409), .C(n_413), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g524 ( .A(n_400), .Y(n_524) );
INVx2_ASAP7_75t_L g647 ( .A(n_400), .Y(n_647) );
OAI21xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_405), .Y(n_401) );
INVx2_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_407), .B(n_447), .Y(n_446) );
INVx4_ASAP7_75t_L g611 ( .A(n_407), .Y(n_611) );
INVx1_ASAP7_75t_L g651 ( .A(n_407), .Y(n_651) );
INVx4_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx3_ASAP7_75t_L g502 ( .A(n_408), .Y(n_502) );
BUFx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx4_ASAP7_75t_L g617 ( .A(n_412), .Y(n_617) );
NAND4xp25_ASAP7_75t_L g416 ( .A(n_417), .B(n_422), .C(n_426), .D(n_434), .Y(n_416) );
BUFx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g452 ( .A(n_421), .Y(n_452) );
INVx1_ASAP7_75t_L g506 ( .A(n_421), .Y(n_506) );
INVx2_ASAP7_75t_L g589 ( .A(n_421), .Y(n_589) );
BUFx8_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_424), .Y(n_511) );
BUFx4f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_432), .Y(n_629) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g474 ( .A(n_438), .Y(n_474) );
AND2x4_ASAP7_75t_L g438 ( .A(n_439), .B(n_467), .Y(n_438) );
AOI21x1_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B(n_455), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_448), .Y(n_441) );
BUFx2_ASAP7_75t_L g468 ( .A(n_442), .Y(n_468) );
INVx4_ASAP7_75t_L g620 ( .A(n_443), .Y(n_620) );
INVx1_ASAP7_75t_L g609 ( .A(n_444), .Y(n_609) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_453), .Y(n_448) );
INVxp67_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g472 ( .A(n_450), .B(n_462), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_453), .Y(n_473) );
INVx1_ASAP7_75t_L g471 ( .A(n_456), .Y(n_471) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_460), .Y(n_456) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g500 ( .A(n_459), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g648 ( .A1(n_459), .A2(n_649), .B(n_650), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_459), .A2(n_684), .B(n_685), .Y(n_683) );
NAND4xp75_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .C(n_472), .D(n_473), .Y(n_467) );
NOR2x1_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_551), .B1(n_569), .B2(n_575), .Y(n_478) );
INVx1_ASAP7_75t_L g575 ( .A(n_479), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_513), .B1(n_514), .B2(n_550), .Y(n_479) );
INVx2_ASAP7_75t_L g550 ( .A(n_480), .Y(n_550) );
XNOR2x1_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_503), .Y(n_482) );
NAND4xp25_ASAP7_75t_L g483 ( .A(n_484), .B(n_489), .C(n_495), .D(n_499), .Y(n_483) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g644 ( .A(n_488), .Y(n_644) );
INVx3_ASAP7_75t_L g688 ( .A(n_488), .Y(n_688) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g623 ( .A(n_493), .Y(n_623) );
INVx2_ASAP7_75t_L g679 ( .A(n_493), .Y(n_679) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx4_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND4xp25_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .C(n_508), .D(n_509), .Y(n_503) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx3_ASAP7_75t_L g656 ( .A(n_511), .Y(n_656) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NAND2x1_ASAP7_75t_L g516 ( .A(n_517), .B(n_543), .Y(n_516) );
NOR3xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_526), .C(n_530), .Y(n_517) );
OAI22xp33_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_521), .B1(n_522), .B2(n_975), .Y(n_518) );
INVx1_ASAP7_75t_L g548 ( .A(n_519), .Y(n_548) );
NOR2xp67_ASAP7_75t_L g526 ( .A(n_521), .B(n_527), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_521), .A2(n_531), .B1(n_532), .B2(n_976), .Y(n_530) );
INVx1_ASAP7_75t_L g545 ( .A(n_522), .Y(n_545) );
INVx1_ASAP7_75t_L g682 ( .A(n_524), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g543 ( .A(n_527), .B(n_544), .C(n_547), .Y(n_543) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g549 ( .A(n_531), .Y(n_549) );
INVx1_ASAP7_75t_L g546 ( .A(n_532), .Y(n_546) );
NOR2x1_ASAP7_75t_L g532 ( .A(n_533), .B(n_538), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B1(n_536), .B2(n_537), .Y(n_533) );
OAI22xp33_ASAP7_75t_L g939 ( .A1(n_537), .A2(n_540), .B1(n_940), .B2(n_941), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B1(n_541), .B2(n_542), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVxp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_564), .Y(n_555) );
NAND4xp25_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .C(n_560), .D(n_562), .Y(n_556) );
BUFx3_ASAP7_75t_L g615 ( .A(n_558), .Y(n_615) );
NAND4xp25_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .C(n_567), .D(n_568), .Y(n_564) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g702 ( .A(n_577), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_632), .B1(n_691), .B2(n_692), .Y(n_577) );
INVx1_ASAP7_75t_L g691 ( .A(n_578), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_580), .B1(n_602), .B2(n_631), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
BUFx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
XNOR2x1_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_585), .Y(n_584) );
NOR2x1_ASAP7_75t_L g586 ( .A(n_587), .B(n_594), .Y(n_586) );
NAND4xp25_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .C(n_592), .D(n_593), .Y(n_587) );
NAND4xp25_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .C(n_598), .D(n_599), .Y(n_594) );
INVx1_ASAP7_75t_L g631 ( .A(n_602), .Y(n_631) );
INVx4_ASAP7_75t_R g602 ( .A(n_603), .Y(n_602) );
XNOR2x1_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
AND2x4_ASAP7_75t_L g605 ( .A(n_606), .B(n_624), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_612), .C(n_618), .Y(n_606) );
OAI21xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B(n_610), .Y(n_607) );
OAI22xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B1(n_616), .B2(n_617), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B1(n_621), .B2(n_622), .Y(n_618) );
INVxp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND4x1_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .C(n_628), .D(n_630), .Y(n_624) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_627), .Y(n_654) );
INVx1_ASAP7_75t_L g692 ( .A(n_632), .Y(n_692) );
OA22x2_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_667), .B1(n_668), .B2(n_690), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_652), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_641), .C(n_645), .Y(n_636) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
BUFx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND4xp25_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .C(n_659), .D(n_663), .Y(n_652) );
BUFx3_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
BUFx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
XOR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_689), .Y(n_669) );
NOR2x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_677), .Y(n_670) );
NAND4xp25_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .C(n_674), .D(n_675), .Y(n_671) );
NAND3xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_680), .C(n_687), .Y(n_677) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
BUFx3_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_699), .C(n_700), .Y(n_695) );
AND2x2_ASAP7_75t_L g948 ( .A(n_696), .B(n_949), .Y(n_948) );
AND2x2_ASAP7_75t_L g968 ( .A(n_696), .B(n_950), .Y(n_968) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OA21x2_ASAP7_75t_L g970 ( .A1(n_697), .A2(n_734), .B(n_971), .Y(n_970) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g711 ( .A(n_698), .B(n_712), .Y(n_711) );
AND3x4_ASAP7_75t_L g733 ( .A(n_698), .B(n_713), .C(n_734), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g949 ( .A(n_699), .B(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_700), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
OAI221xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_915), .B1(n_917), .B2(n_946), .C(n_951), .Y(n_704) );
AOI211xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_723), .B(n_802), .C(n_911), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI221xp5_ASAP7_75t_SL g832 ( .A1(n_707), .A2(n_831), .B1(n_833), .B2(n_834), .C(n_835), .Y(n_832) );
INVx1_ASAP7_75t_L g875 ( .A(n_707), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_707), .B(n_807), .Y(n_887) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
HB1xp67_ASAP7_75t_L g901 ( .A(n_708), .Y(n_901) );
OAI221xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_715), .B1(n_716), .B2(n_718), .C(n_719), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_709), .A2(n_716), .B1(n_768), .B2(n_769), .Y(n_767) );
INVx3_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_711), .B(n_713), .Y(n_710) );
AND2x4_ASAP7_75t_L g720 ( .A(n_711), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g727 ( .A(n_711), .B(n_721), .Y(n_727) );
AND2x2_ASAP7_75t_L g737 ( .A(n_711), .B(n_721), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_713), .B(n_717), .Y(n_716) );
AND2x4_ASAP7_75t_L g730 ( .A(n_713), .B(n_717), .Y(n_730) );
AND2x4_ASAP7_75t_L g735 ( .A(n_713), .B(n_717), .Y(n_735) );
AND2x4_ASAP7_75t_L g722 ( .A(n_717), .B(n_721), .Y(n_722) );
AND2x2_ASAP7_75t_L g728 ( .A(n_717), .B(n_721), .Y(n_728) );
AND2x2_ASAP7_75t_L g738 ( .A(n_717), .B(n_721), .Y(n_738) );
INVx3_ASAP7_75t_L g771 ( .A(n_720), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g971 ( .A(n_721), .Y(n_971) );
INVx2_ASAP7_75t_L g773 ( .A(n_722), .Y(n_773) );
BUFx2_ASAP7_75t_L g916 ( .A(n_722), .Y(n_916) );
OAI211xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_739), .B(n_752), .C(n_792), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_724), .B(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g795 ( .A(n_724), .Y(n_795) );
OR2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_731), .Y(n_724) );
INVx1_ASAP7_75t_L g808 ( .A(n_725), .Y(n_808) );
INVx1_ASAP7_75t_L g820 ( .A(n_725), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_729), .Y(n_725) );
AND2x2_ASAP7_75t_L g765 ( .A(n_731), .B(n_766), .Y(n_765) );
OR2x2_ASAP7_75t_L g801 ( .A(n_731), .B(n_766), .Y(n_801) );
INVx2_ASAP7_75t_L g827 ( .A(n_731), .Y(n_827) );
OR2x2_ASAP7_75t_L g835 ( .A(n_731), .B(n_820), .Y(n_835) );
AND2x2_ASAP7_75t_L g844 ( .A(n_731), .B(n_820), .Y(n_844) );
OR2x2_ASAP7_75t_L g848 ( .A(n_731), .B(n_780), .Y(n_848) );
AND2x2_ASAP7_75t_L g874 ( .A(n_731), .B(n_819), .Y(n_874) );
HB1xp67_ASAP7_75t_L g882 ( .A(n_731), .Y(n_882) );
AND2x2_ASAP7_75t_L g886 ( .A(n_731), .B(n_780), .Y(n_886) );
AND2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_736), .Y(n_731) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI31xp33_ASAP7_75t_L g792 ( .A1(n_740), .A2(n_761), .A3(n_793), .B(n_799), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_740), .A2(n_797), .B1(n_801), .B2(n_816), .Y(n_815) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_745), .Y(n_740) );
AND2x2_ASAP7_75t_L g822 ( .A(n_741), .B(n_754), .Y(n_822) );
AND2x2_ASAP7_75t_L g845 ( .A(n_741), .B(n_798), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_741), .B(n_749), .Y(n_852) );
AND2x2_ASAP7_75t_L g907 ( .A(n_741), .B(n_760), .Y(n_907) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g753 ( .A(n_742), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g763 ( .A(n_742), .Y(n_763) );
AND2x2_ASAP7_75t_L g797 ( .A(n_742), .B(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_742), .B(n_749), .Y(n_831) );
OR2x2_ASAP7_75t_L g837 ( .A(n_742), .B(n_759), .Y(n_837) );
AOI221xp5_ASAP7_75t_L g842 ( .A1(n_742), .A2(n_843), .B1(n_845), .B2(n_846), .C(n_849), .Y(n_842) );
OR2x2_ASAP7_75t_L g850 ( .A(n_742), .B(n_784), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_742), .B(n_839), .Y(n_879) );
AND2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_745), .B(n_811), .Y(n_833) );
AND2x2_ASAP7_75t_L g872 ( .A(n_745), .B(n_762), .Y(n_872) );
INVx1_ASAP7_75t_L g884 ( .A(n_745), .Y(n_884) );
AND2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_749), .Y(n_745) );
OR2x2_ASAP7_75t_L g759 ( .A(n_746), .B(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g764 ( .A(n_746), .B(n_760), .Y(n_764) );
OR2x2_ASAP7_75t_L g784 ( .A(n_746), .B(n_749), .Y(n_784) );
INVx1_ASAP7_75t_L g798 ( .A(n_746), .Y(n_798) );
OAI221xp5_ASAP7_75t_L g804 ( .A1(n_746), .A2(n_805), .B1(n_815), .B2(n_818), .C(n_821), .Y(n_804) );
AND2x2_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_L g760 ( .A(n_749), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_749), .A2(n_881), .B1(n_883), .B2(n_885), .Y(n_880) );
AND2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
O2A1O1Ixp33_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_761), .B(n_765), .C(n_775), .Y(n_752) );
NOR2x1_ASAP7_75t_L g754 ( .A(n_755), .B(n_759), .Y(n_754) );
AND2x2_ASAP7_75t_L g777 ( .A(n_755), .B(n_766), .Y(n_777) );
AND2x2_ASAP7_75t_L g796 ( .A(n_755), .B(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g800 ( .A(n_755), .Y(n_800) );
INVx2_ASAP7_75t_L g811 ( .A(n_755), .Y(n_811) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_755), .Y(n_813) );
NAND2xp5_ASAP7_75t_SL g829 ( .A(n_755), .B(n_830), .Y(n_829) );
AND2x2_ASAP7_75t_L g839 ( .A(n_755), .B(n_764), .Y(n_839) );
INVx2_ASAP7_75t_L g859 ( .A(n_755), .Y(n_859) );
NOR2xp33_ASAP7_75t_L g908 ( .A(n_755), .B(n_808), .Y(n_908) );
INVx4_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OR2x2_ASAP7_75t_L g791 ( .A(n_756), .B(n_762), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_756), .B(n_780), .Y(n_817) );
AND2x2_ASAP7_75t_L g855 ( .A(n_756), .B(n_766), .Y(n_855) );
AND2x2_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx3_ASAP7_75t_SL g868 ( .A(n_759), .Y(n_868) );
NAND2xp67_ASAP7_75t_L g904 ( .A(n_761), .B(n_811), .Y(n_904) );
AND2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_764), .Y(n_761) );
AND2x4_ASAP7_75t_L g782 ( .A(n_762), .B(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g790 ( .A(n_764), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_764), .B(n_854), .Y(n_853) );
OAI21xp5_ASAP7_75t_L g906 ( .A1(n_764), .A2(n_907), .B(n_908), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_765), .B(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g834 ( .A(n_765), .Y(n_834) );
AOI221xp5_ASAP7_75t_L g902 ( .A1(n_765), .A2(n_830), .B1(n_846), .B2(n_903), .C(n_905), .Y(n_902) );
INVx2_ASAP7_75t_L g780 ( .A(n_766), .Y(n_780) );
INVx1_ASAP7_75t_L g787 ( .A(n_766), .Y(n_787) );
AND2x2_ASAP7_75t_L g843 ( .A(n_766), .B(n_844), .Y(n_843) );
OR2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_770), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_770) );
A2O1A1Ixp33_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_778), .B(n_781), .C(n_785), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_777), .B(n_807), .Y(n_851) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AND2x2_ASAP7_75t_L g841 ( .A(n_780), .B(n_808), .Y(n_841) );
INVx2_ASAP7_75t_L g857 ( .A(n_780), .Y(n_857) );
INVx2_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_782), .B(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_784), .B(n_884), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_786), .B(n_818), .Y(n_898) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_787), .B(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_789), .B(n_834), .Y(n_910) );
OR2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
INVx1_ASAP7_75t_L g867 ( .A(n_791), .Y(n_867) );
INVxp33_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
O2A1O1Ixp33_ASAP7_75t_L g909 ( .A1(n_796), .A2(n_847), .B(n_872), .C(n_910), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_800), .B(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g814 ( .A(n_801), .Y(n_814) );
OAI221xp5_ASAP7_75t_L g849 ( .A1(n_801), .A2(n_850), .B1(n_851), .B2(n_852), .C(n_853), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_801), .A2(n_829), .B1(n_835), .B2(n_906), .Y(n_905) );
NAND5xp2_ASAP7_75t_L g802 ( .A(n_803), .B(n_876), .C(n_896), .D(n_902), .E(n_909), .Y(n_802) );
OAI21xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_823), .B(n_861), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_809), .B1(n_812), .B2(n_814), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
AND2x2_ASAP7_75t_L g846 ( .A(n_807), .B(n_847), .Y(n_846) );
AOI21xp33_ASAP7_75t_L g911 ( .A1(n_807), .A2(n_912), .B(n_914), .Y(n_911) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
BUFx3_ASAP7_75t_L g893 ( .A(n_808), .Y(n_893) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_812), .B(n_886), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_812), .B(n_890), .Y(n_889) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_813), .B(n_871), .Y(n_870) );
OAI21xp33_ASAP7_75t_SL g877 ( .A1(n_813), .A2(n_878), .B(n_879), .Y(n_877) );
AND2x2_ASAP7_75t_L g892 ( .A(n_814), .B(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g914 ( .A(n_822), .Y(n_914) );
NAND3xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_842), .C(n_856), .Y(n_823) );
AOI211xp5_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_828), .B(n_832), .C(n_836), .Y(n_824) );
CKINVDCx14_ASAP7_75t_R g825 ( .A(n_826), .Y(n_825) );
CKINVDCx14_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
AND2x2_ASAP7_75t_L g854 ( .A(n_827), .B(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
AOI21xp33_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B(n_840), .Y(n_836) );
INVx1_ASAP7_75t_L g895 ( .A(n_837), .Y(n_895) );
A2O1A1Ixp33_ASAP7_75t_L g888 ( .A1(n_838), .A2(n_889), .B(n_891), .C(n_894), .Y(n_888) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_843), .B(n_895), .Y(n_894) );
AOI221xp5_ASAP7_75t_L g876 ( .A1(n_844), .A2(n_877), .B1(n_880), .B2(n_887), .C(n_888), .Y(n_876) );
INVx1_ASAP7_75t_L g878 ( .A(n_845), .Y(n_878) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g860 ( .A(n_850), .Y(n_860) );
INVx1_ASAP7_75t_L g890 ( .A(n_852), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_857), .B(n_858), .Y(n_856) );
INVx2_ASAP7_75t_L g869 ( .A(n_857), .Y(n_869) );
AND2x2_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
INVx1_ASAP7_75t_L g863 ( .A(n_859), .Y(n_863) );
A2O1A1Ixp33_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_864), .B(n_873), .C(n_875), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_863), .B(n_872), .Y(n_900) );
AOI21xp5_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_869), .B(n_870), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
NOR2xp33_ASAP7_75t_L g913 ( .A(n_869), .B(n_904), .Y(n_913) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
OAI211xp5_ASAP7_75t_L g896 ( .A1(n_886), .A2(n_897), .B(n_899), .C(n_901), .Y(n_896) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVxp67_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_916), .Y(n_915) );
INVxp67_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
HB1xp67_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
XNOR2x1_ASAP7_75t_L g922 ( .A(n_923), .B(n_924), .Y(n_922) );
AND2x2_ASAP7_75t_L g924 ( .A(n_925), .B(n_932), .Y(n_924) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_926), .B(n_929), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_927), .B(n_928), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_930), .B(n_931), .Y(n_929) );
NOR3xp33_ASAP7_75t_L g932 ( .A(n_933), .B(n_939), .C(n_942), .Y(n_932) );
OAI21xp33_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_935), .B(n_936), .Y(n_933) );
OAI21xp5_ASAP7_75t_SL g942 ( .A1(n_943), .A2(n_944), .B(n_945), .Y(n_942) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
HB1xp67_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g966 ( .A(n_954), .Y(n_966) );
HB1xp67_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
OR2x2_ASAP7_75t_L g955 ( .A(n_956), .B(n_961), .Y(n_955) );
NAND4xp25_ASAP7_75t_L g956 ( .A(n_957), .B(n_958), .C(n_959), .D(n_960), .Y(n_956) );
NAND4xp25_ASAP7_75t_L g961 ( .A(n_962), .B(n_963), .C(n_964), .D(n_965), .Y(n_961) );
HB1xp67_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
endmodule