module fake_jpeg_12022_n_470 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_470);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_470;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_7),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_90),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_16),
.B(n_7),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_53),
.B(n_13),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g122 ( 
.A(n_77),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_87),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_7),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_91),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_41),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_93),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_28),
.Y(n_106)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_96),
.Y(n_100)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_106),
.B(n_58),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_56),
.B(n_21),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_113),
.B(n_126),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_80),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_116),
.B(n_147),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_57),
.A2(n_28),
.B1(n_39),
.B2(n_48),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_119),
.A2(n_133),
.B(n_151),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_61),
.A2(n_39),
.B1(n_46),
.B2(n_26),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_92),
.A2(n_41),
.B(n_24),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_135),
.B(n_20),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_50),
.A2(n_39),
.B1(n_30),
.B2(n_43),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_146),
.A2(n_150),
.B1(n_36),
.B2(n_30),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_69),
.B(n_19),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_82),
.B(n_38),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_37),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_64),
.A2(n_38),
.B1(n_36),
.B2(n_43),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_70),
.A2(n_32),
.B1(n_46),
.B2(n_27),
.Y(n_151)
);

INVx4_ASAP7_75t_SL g152 ( 
.A(n_117),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_152),
.B(n_161),
.Y(n_219)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_153),
.Y(n_202)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_112),
.A2(n_52),
.B1(n_58),
.B2(n_72),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_159),
.A2(n_188),
.B1(n_197),
.B2(n_198),
.Y(n_239)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_117),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_170),
.Y(n_207)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_98),
.A2(n_133),
.B1(n_119),
.B2(n_106),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_166),
.A2(n_176),
.B1(n_184),
.B2(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_167),
.Y(n_228)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_105),
.A2(n_94),
.B1(n_89),
.B2(n_54),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g225 ( 
.A1(n_169),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.Y(n_225)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_99),
.B(n_85),
.CI(n_72),
.CON(n_170),
.SN(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_171),
.Y(n_235)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_173),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_174),
.B(n_191),
.Y(n_231)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_175),
.Y(n_236)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_178),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_186),
.Y(n_208)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_183),
.Y(n_227)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_101),
.A2(n_68),
.B1(n_83),
.B2(n_87),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_110),
.A2(n_75),
.B1(n_73),
.B2(n_62),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_130),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_189),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

BUFx12_ASAP7_75t_L g190 ( 
.A(n_130),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_40),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_112),
.B(n_40),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_194),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_120),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_101),
.B(n_23),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_196),
.Y(n_237)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_141),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_136),
.B(n_88),
.Y(n_199)
);

NOR2xp67_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_200),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_37),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_213),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_20),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_161),
.B(n_142),
.C(n_110),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_217),
.C(n_199),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_152),
.B(n_23),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_139),
.B1(n_115),
.B2(n_114),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_218),
.A2(n_220),
.B1(n_188),
.B2(n_179),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_164),
.A2(n_114),
.B1(n_115),
.B2(n_137),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_35),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_221),
.B(n_233),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_169),
.A2(n_78),
.B1(n_79),
.B2(n_91),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_224),
.A2(n_226),
.B1(n_186),
.B2(n_216),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_225),
.A2(n_132),
.B1(n_177),
.B2(n_32),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_169),
.A2(n_159),
.B1(n_137),
.B2(n_140),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_182),
.B(n_35),
.Y(n_233)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_201),
.Y(n_241)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_241),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_242),
.A2(n_266),
.B1(n_225),
.B2(n_215),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_237),
.B(n_183),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_243),
.B(n_246),
.Y(n_288)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_213),
.B(n_193),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_247),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_208),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_219),
.A2(n_170),
.B1(n_194),
.B2(n_198),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_249),
.A2(n_251),
.B(n_273),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_231),
.B(n_160),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_268),
.Y(n_293)
);

NOR2x1_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_86),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_253),
.A2(n_254),
.B1(n_259),
.B2(n_261),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_230),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_258),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_204),
.B(n_24),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_256),
.B(n_274),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_207),
.A2(n_219),
.B(n_239),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_267),
.B(n_223),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_230),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_224),
.A2(n_81),
.B1(n_131),
.B2(n_138),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_210),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_260),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_205),
.A2(n_131),
.B1(n_138),
.B2(n_29),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_211),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_262),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_205),
.A2(n_27),
.B1(n_46),
.B2(n_29),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_264),
.A2(n_265),
.B1(n_209),
.B2(n_234),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_220),
.A2(n_27),
.B1(n_46),
.B2(n_29),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_225),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_240),
.A2(n_132),
.B(n_178),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_221),
.B(n_0),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_222),
.B(n_233),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_269),
.B(n_271),
.Y(n_304)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_211),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_244),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_1),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_206),
.B(n_86),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_275),
.C(n_276),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_225),
.A2(n_32),
.B1(n_122),
.B2(n_41),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_204),
.B(n_10),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_190),
.C(n_122),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_228),
.B(n_190),
.C(n_47),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_279),
.A2(n_296),
.B(n_252),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_281),
.A2(n_214),
.B1(n_202),
.B2(n_229),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_257),
.A2(n_249),
.B(n_267),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_283),
.A2(n_306),
.B(n_214),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_256),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_284),
.B(n_285),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_251),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_292),
.C(n_305),
.Y(n_315)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_248),
.B(n_230),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_250),
.B(n_243),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_242),
.A2(n_255),
.B1(n_258),
.B2(n_269),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_246),
.B(n_215),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_309),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_299),
.A2(n_265),
.B1(n_245),
.B2(n_262),
.Y(n_323)
);

BUFx8_ASAP7_75t_L g301 ( 
.A(n_251),
.Y(n_301)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_254),
.A2(n_209),
.B1(n_234),
.B2(n_238),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_302),
.A2(n_235),
.B1(n_202),
.B2(n_212),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_260),
.Y(n_303)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_227),
.C(n_238),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_273),
.A2(n_227),
.B(n_210),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_241),
.Y(n_307)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_274),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_263),
.B(n_268),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_252),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_296),
.A2(n_264),
.B1(n_261),
.B2(n_253),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_311),
.A2(n_323),
.B1(n_328),
.B2(n_335),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_283),
.A2(n_275),
.B(n_263),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_318),
.A2(n_339),
.B(n_313),
.Y(n_341)
);

AOI22x1_ASAP7_75t_L g320 ( 
.A1(n_286),
.A2(n_266),
.B1(n_259),
.B2(n_270),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_320),
.A2(n_330),
.B1(n_340),
.B2(n_287),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_321),
.B(n_322),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_247),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_327),
.Y(n_358)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_290),
.Y(n_325)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_325),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_278),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_278),
.A2(n_276),
.B1(n_271),
.B2(n_232),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_227),
.Y(n_329)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_329),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_288),
.Y(n_331)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_331),
.Y(n_357)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_297),
.Y(n_332)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_332),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_288),
.B(n_203),
.Y(n_333)
);

NAND2xp33_ASAP7_75t_SL g346 ( 
.A(n_333),
.B(n_334),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_277),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_286),
.A2(n_232),
.B1(n_203),
.B2(n_212),
.Y(n_335)
);

OAI21x1_ASAP7_75t_R g336 ( 
.A1(n_301),
.A2(n_308),
.B(n_300),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_336),
.A2(n_339),
.B(n_301),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_289),
.B(n_235),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_338),
.B(n_305),
.C(n_282),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_341),
.A2(n_366),
.B(n_346),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_348),
.C(n_350),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_327),
.A2(n_295),
.B1(n_284),
.B2(n_293),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_345),
.A2(n_332),
.B1(n_336),
.B2(n_319),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_312),
.Y(n_347)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_347),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_315),
.B(n_292),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_282),
.C(n_293),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_311),
.A2(n_302),
.B1(n_281),
.B2(n_277),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_352),
.A2(n_356),
.B1(n_325),
.B2(n_337),
.Y(n_376)
);

BUFx5_ASAP7_75t_L g353 ( 
.A(n_312),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_353),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_304),
.C(n_291),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_354),
.B(n_360),
.C(n_361),
.Y(n_378)
);

INVxp33_ASAP7_75t_L g381 ( 
.A(n_355),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_335),
.A2(n_291),
.B1(n_280),
.B2(n_308),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_304),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_300),
.C(n_297),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_322),
.B(n_298),
.Y(n_362)
);

XOR2x2_ASAP7_75t_L g372 ( 
.A(n_362),
.B(n_360),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_306),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_326),
.C(n_329),
.Y(n_379)
);

INVxp33_ASAP7_75t_L g382 ( 
.A(n_365),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_321),
.A2(n_301),
.B(n_280),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_314),
.Y(n_367)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_367),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_361),
.B(n_316),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_369),
.B(n_385),
.Y(n_408)
);

A2O1A1Ixp33_ASAP7_75t_SL g371 ( 
.A1(n_341),
.A2(n_336),
.B(n_337),
.C(n_320),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_371),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_372),
.B(n_373),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_317),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_374),
.A2(n_366),
.B(n_355),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_376),
.A2(n_386),
.B1(n_387),
.B2(n_349),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_317),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_377),
.B(n_351),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_379),
.B(n_345),
.Y(n_396)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_358),
.Y(n_380)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_380),
.Y(n_393)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_343),
.Y(n_383)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_357),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_349),
.A2(n_333),
.B1(n_330),
.B2(n_320),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_364),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_342),
.B(n_334),
.C(n_333),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_388),
.B(n_389),
.C(n_359),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_354),
.B(n_359),
.C(n_363),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_390),
.A2(n_367),
.B1(n_307),
.B2(n_287),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_391),
.A2(n_381),
.B(n_371),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_392),
.B(n_395),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_396),
.B(n_389),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_368),
.B(n_362),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_404),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_374),
.A2(n_356),
.B(n_344),
.Y(n_398)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_398),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_399),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_382),
.A2(n_352),
.B1(n_353),
.B2(n_319),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_400),
.A2(n_409),
.B1(n_384),
.B2(n_370),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_401),
.A2(n_384),
.B1(n_375),
.B2(n_379),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_390),
.A2(n_314),
.B1(n_294),
.B2(n_303),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_403),
.B(n_405),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_368),
.B(n_229),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_373),
.B(n_294),
.C(n_47),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_294),
.C(n_2),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_406),
.B(n_388),
.C(n_384),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_382),
.A2(n_8),
.B1(n_13),
.B2(n_3),
.Y(n_409)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_410),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_395),
.B(n_377),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_420),
.Y(n_425)
);

OA21x2_ASAP7_75t_L g413 ( 
.A1(n_407),
.A2(n_381),
.B(n_371),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_413),
.B(n_1),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_417),
.Y(n_426)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_402),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_421),
.A2(n_400),
.B(n_409),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_422),
.A2(n_423),
.B1(n_6),
.B2(n_12),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_391),
.A2(n_371),
.B1(n_372),
.B2(n_378),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_393),
.A2(n_8),
.B1(n_12),
.B2(n_3),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_424),
.B(n_408),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_423),
.A2(n_392),
.B(n_406),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_427),
.B(n_428),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_404),
.C(n_397),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_429),
.B(n_433),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_416),
.A2(n_396),
.B1(n_405),
.B2(n_394),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_430),
.B(n_420),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_431),
.B(n_432),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_418),
.B(n_394),
.C(n_2),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_8),
.Y(n_434)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_434),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_436),
.A2(n_413),
.B1(n_9),
.B2(n_3),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_6),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_437),
.B(n_422),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_426),
.A2(n_415),
.B(n_421),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_439),
.A2(n_429),
.B(n_6),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_445),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_441),
.B(n_446),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_411),
.Y(n_442)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_442),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_419),
.C(n_413),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_435),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_447),
.B(n_425),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_444),
.A2(n_436),
.B1(n_433),
.B2(n_432),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_449),
.B(n_451),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_448),
.B(n_419),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_452),
.B(n_453),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_442),
.B(n_430),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_456),
.A2(n_438),
.B(n_6),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_450),
.A2(n_443),
.B(n_441),
.Y(n_458)
);

AOI21x1_ASAP7_75t_L g463 ( 
.A1(n_458),
.A2(n_452),
.B(n_3),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_459),
.B(n_4),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_455),
.A2(n_438),
.B(n_10),
.Y(n_460)
);

AOI21xp33_ASAP7_75t_L g462 ( 
.A1(n_460),
.A2(n_454),
.B(n_461),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_462),
.Y(n_465)
);

O2A1O1Ixp33_ASAP7_75t_SL g466 ( 
.A1(n_463),
.A2(n_464),
.B(n_4),
.C(n_12),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_466),
.B(n_465),
.C(n_457),
.Y(n_467)
);

BUFx24_ASAP7_75t_SL g468 ( 
.A(n_467),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_468),
.A2(n_14),
.B(n_1),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_469),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_470)
);


endmodule