module fake_jpeg_11887_n_510 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_510);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_510;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_51),
.Y(n_133)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_20),
.B(n_9),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_58),
.B(n_63),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_8),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_70),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_75),
.Y(n_156)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_29),
.B(n_8),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_79),
.B(n_88),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_29),
.B(n_11),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_84),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_37),
.B(n_39),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_85),
.Y(n_155)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_91),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_95),
.Y(n_107)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_96),
.Y(n_102)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_51),
.A2(n_56),
.B1(n_55),
.B2(n_53),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_97),
.A2(n_145),
.B1(n_148),
.B2(n_22),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_66),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_103),
.A2(n_116),
.B1(n_121),
.B2(n_128),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_37),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_108),
.B(n_114),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_39),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_59),
.A2(n_31),
.B1(n_27),
.B2(n_33),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_77),
.A2(n_32),
.B1(n_27),
.B2(n_28),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_42),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_130),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_67),
.A2(n_32),
.B1(n_27),
.B2(n_28),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_42),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_61),
.B(n_40),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_134),
.B(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_69),
.B(n_40),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_136),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_48),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_74),
.A2(n_32),
.B1(n_25),
.B2(n_28),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_75),
.A2(n_33),
.B1(n_25),
.B2(n_31),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_82),
.B(n_48),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_157),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_83),
.B(n_26),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_85),
.B(n_38),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_17),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_87),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_45),
.B1(n_44),
.B2(n_35),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_91),
.B(n_38),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_158),
.Y(n_221)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_160),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_116),
.A2(n_92),
.B1(n_31),
.B2(n_33),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_161),
.A2(n_168),
.B1(n_173),
.B2(n_195),
.Y(n_240)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_163),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_164),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_165),
.A2(n_213),
.B1(n_214),
.B2(n_129),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_132),
.A2(n_45),
.B1(n_44),
.B2(n_35),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_166),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_167),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_98),
.A2(n_45),
.B1(n_44),
.B2(n_35),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_99),
.B(n_119),
.C(n_101),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_169),
.B(n_175),
.C(n_194),
.Y(n_222)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_170),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_171),
.B(n_177),
.Y(n_234)
);

NAND2xp33_ASAP7_75t_SL g172 ( 
.A(n_149),
.B(n_64),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_172),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_154),
.B1(n_128),
.B2(n_103),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_22),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_176),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_111),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_179),
.Y(n_259)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_102),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_182),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_155),
.Y(n_182)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_185),
.Y(n_241)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_140),
.Y(n_186)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_142),
.A2(n_22),
.B1(n_60),
.B2(n_12),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_188),
.A2(n_207),
.B1(n_146),
.B2(n_139),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_105),
.B(n_0),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_191),
.Y(n_220)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_190),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_105),
.B(n_0),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_192),
.Y(n_252)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_126),
.Y(n_193)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_118),
.B(n_0),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_121),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_111),
.Y(n_196)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_97),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_197)
);

AO22x1_ASAP7_75t_L g227 ( 
.A1(n_197),
.A2(n_143),
.B1(n_113),
.B2(n_156),
.Y(n_227)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_198),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_206),
.Y(n_236)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_200),
.Y(n_260)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_201),
.Y(n_265)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_203),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_118),
.B(n_11),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_204),
.B(n_205),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_142),
.B(n_11),
.CI(n_16),
.CON(n_205),
.SN(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_141),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_127),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_125),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_208),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_115),
.A2(n_7),
.B(n_15),
.C(n_14),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_210),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_109),
.B(n_1),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_211),
.B(n_200),
.Y(n_263)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_131),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_215),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_109),
.A2(n_12),
.B1(n_15),
.B2(n_4),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_129),
.A2(n_12),
.B1(n_14),
.B2(n_4),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_120),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_127),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_216),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_172),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_217),
.B(n_228),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_223),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_195),
.A2(n_139),
.B1(n_146),
.B2(n_138),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_226),
.A2(n_164),
.B1(n_167),
.B2(n_178),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_227),
.A2(n_242),
.B(n_196),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_158),
.A2(n_150),
.B1(n_156),
.B2(n_143),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_229),
.A2(n_239),
.B1(n_255),
.B2(n_234),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_237),
.A2(n_247),
.B1(n_191),
.B2(n_189),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_175),
.B(n_138),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_258),
.C(n_169),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_160),
.A2(n_113),
.B1(n_115),
.B2(n_120),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_162),
.A2(n_122),
.B1(n_141),
.B2(n_5),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_122),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_246),
.B(n_262),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_161),
.A2(n_5),
.B1(n_13),
.B2(n_17),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_187),
.B(n_2),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_183),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_187),
.B(n_5),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_194),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_263),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_184),
.B(n_5),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_267),
.B(n_3),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_240),
.A2(n_171),
.B1(n_183),
.B2(n_174),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_268),
.A2(n_275),
.B1(n_277),
.B2(n_297),
.Y(n_315)
);

AO22x1_ASAP7_75t_L g269 ( 
.A1(n_230),
.A2(n_197),
.B1(n_205),
.B2(n_209),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_269),
.A2(n_278),
.B(n_294),
.Y(n_334)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_271),
.B(n_274),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_253),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_272),
.B(n_290),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_220),
.B(n_210),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_276),
.B(n_258),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_240),
.A2(n_174),
.B1(n_197),
.B2(n_192),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_230),
.A2(n_196),
.B(n_177),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_222),
.B(n_185),
.C(n_202),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_279),
.B(n_282),
.C(n_292),
.Y(n_318)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_235),
.Y(n_280)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_280),
.Y(n_322)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_222),
.B(n_238),
.Y(n_282)
);

INVx11_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

BUFx5_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_264),
.Y(n_284)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_284),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_220),
.B(n_233),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_286),
.B(n_288),
.Y(n_345)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_289),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_231),
.Y(n_290)
);

AO21x2_ASAP7_75t_L g291 ( 
.A1(n_227),
.A2(n_197),
.B(n_186),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_291),
.A2(n_255),
.B1(n_259),
.B2(n_232),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_238),
.B(n_163),
.C(n_170),
.Y(n_292)
);

NOR2x1_ASAP7_75t_L g293 ( 
.A(n_219),
.B(n_201),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_293),
.B(n_295),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_249),
.A2(n_190),
.B(n_179),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_233),
.B(n_159),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_251),
.Y(n_296)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_296),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_237),
.A2(n_208),
.B1(n_180),
.B2(n_203),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_221),
.A2(n_224),
.B1(n_242),
.B2(n_246),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_298),
.A2(n_304),
.B1(n_313),
.B2(n_261),
.Y(n_337)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_252),
.Y(n_299)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_299),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_300),
.A2(n_301),
.B1(n_302),
.B2(n_311),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_234),
.A2(n_211),
.B1(n_13),
.B2(n_17),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_234),
.A2(n_3),
.B1(n_13),
.B2(n_249),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_252),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_303),
.B(n_305),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_221),
.A2(n_224),
.B1(n_262),
.B2(n_219),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_218),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_306),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_256),
.B(n_3),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_254),
.Y(n_339)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_218),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_308),
.Y(n_350)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_309),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_236),
.B(n_3),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_310),
.A2(n_260),
.B(n_257),
.Y(n_324)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_248),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_312),
.A2(n_294),
.B(n_278),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_227),
.A2(n_244),
.B1(n_250),
.B2(n_243),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_316),
.B(n_323),
.C(n_327),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_291),
.A2(n_250),
.B1(n_244),
.B2(n_243),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_319),
.A2(n_321),
.B1(n_329),
.B2(n_331),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_282),
.B(n_263),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_320),
.B(n_332),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_279),
.B(n_257),
.C(n_263),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_324),
.B(n_350),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_276),
.B(n_241),
.C(n_260),
.Y(n_327)
);

OAI32xp33_ASAP7_75t_L g328 ( 
.A1(n_286),
.A2(n_232),
.A3(n_225),
.B1(n_241),
.B2(n_265),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_303),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_291),
.A2(n_295),
.B1(n_268),
.B2(n_277),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_291),
.A2(n_245),
.B1(n_254),
.B2(n_259),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_274),
.B(n_225),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_265),
.C(n_254),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_352),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_336),
.B(n_341),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_337),
.A2(n_341),
.B1(n_346),
.B2(n_351),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_287),
.A2(n_261),
.B(n_245),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_338),
.A2(n_283),
.B(n_281),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_309),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_313),
.A2(n_297),
.B1(n_314),
.B2(n_291),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_314),
.A2(n_288),
.B1(n_271),
.B2(n_269),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_312),
.A2(n_273),
.B1(n_269),
.B2(n_285),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_349),
.A2(n_352),
.B1(n_319),
.B2(n_345),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_285),
.A2(n_270),
.B1(n_280),
.B2(n_290),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_293),
.B(n_307),
.Y(n_352)
);

OAI32xp33_ASAP7_75t_L g357 ( 
.A1(n_347),
.A2(n_345),
.A3(n_349),
.B1(n_330),
.B2(n_329),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_357),
.B(n_358),
.Y(n_410)
);

A2O1A1Ixp33_ASAP7_75t_L g358 ( 
.A1(n_334),
.A2(n_289),
.B(n_284),
.C(n_310),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_318),
.B(n_285),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_359),
.B(n_361),
.C(n_362),
.Y(n_399)
);

AO21x1_ASAP7_75t_L g394 ( 
.A1(n_360),
.A2(n_381),
.B(n_382),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_318),
.B(n_272),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_308),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_317),
.Y(n_363)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_363),
.Y(n_400)
);

BUFx4f_ASAP7_75t_SL g364 ( 
.A(n_326),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_364),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_299),
.Y(n_365)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_353),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_366),
.B(n_376),
.Y(n_413)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_317),
.Y(n_367)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_355),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_334),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_371),
.B(n_388),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_320),
.B(n_306),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_383),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_311),
.Y(n_374)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_346),
.A2(n_296),
.B1(n_305),
.B2(n_315),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_375),
.A2(n_324),
.B1(n_340),
.B2(n_350),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_354),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_377),
.A2(n_360),
.B1(n_372),
.B2(n_357),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_321),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_378),
.B(n_386),
.Y(n_417)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_322),
.Y(n_380)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_380),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_323),
.B(n_327),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_336),
.A2(n_338),
.B(n_347),
.Y(n_384)
);

AO21x1_ASAP7_75t_L g390 ( 
.A1(n_384),
.A2(n_382),
.B(n_371),
.Y(n_390)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_322),
.Y(n_385)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_332),
.B(n_337),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_328),
.B(n_340),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_315),
.B(n_333),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_348),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_390),
.A2(n_406),
.B(n_410),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_377),
.A2(n_331),
.B1(n_342),
.B2(n_343),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_392),
.A2(n_393),
.B1(n_405),
.B2(n_407),
.Y(n_420)
);

OAI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_370),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_395),
.B(n_397),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_365),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_398),
.A2(n_414),
.B1(n_409),
.B2(n_394),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_374),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_402),
.B(n_404),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_384),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g427 ( 
.A(n_403),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_388),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_370),
.A2(n_355),
.B1(n_325),
.B2(n_335),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_361),
.B(n_335),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_412),
.B(n_356),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_375),
.A2(n_325),
.B1(n_348),
.B2(n_326),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_416),
.B(n_359),
.C(n_356),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_419),
.B(n_422),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_421),
.B(n_422),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_396),
.B(n_362),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_399),
.B(n_383),
.C(n_387),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_429),
.C(n_430),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_418),
.A2(n_382),
.B(n_369),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_425),
.B(n_433),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_387),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_424),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_389),
.C(n_373),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_396),
.B(n_412),
.C(n_379),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_397),
.B(n_358),
.Y(n_431)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_431),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_418),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_436),
.Y(n_456)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_417),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_404),
.A2(n_364),
.B1(n_379),
.B2(n_398),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_434),
.A2(n_391),
.B1(n_400),
.B2(n_408),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_395),
.B(n_364),
.C(n_413),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_442),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_405),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_394),
.B(n_410),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_437),
.B(n_400),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_438),
.B(n_440),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_392),
.A2(n_402),
.B1(n_409),
.B2(n_406),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_439),
.A2(n_408),
.B1(n_411),
.B2(n_415),
.Y(n_448)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_401),
.Y(n_441)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_441),
.Y(n_457)
);

FAx1_ASAP7_75t_SL g442 ( 
.A(n_390),
.B(n_401),
.CI(n_414),
.CON(n_442),
.SN(n_442)
);

OAI21x1_ASAP7_75t_L g445 ( 
.A1(n_423),
.A2(n_390),
.B(n_391),
.Y(n_445)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_445),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_446),
.B(n_458),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_447),
.A2(n_448),
.B1(n_449),
.B2(n_440),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_420),
.A2(n_411),
.B1(n_415),
.B2(n_432),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_454),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_426),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_453),
.B(n_461),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_421),
.Y(n_454)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_441),
.Y(n_459)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_459),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_419),
.B(n_429),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_423),
.B(n_426),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_462),
.B(n_431),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_463),
.A2(n_472),
.B(n_460),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_464),
.A2(n_469),
.B1(n_472),
.B2(n_463),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_452),
.B(n_435),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_465),
.B(n_456),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_430),
.C(n_434),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_468),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_462),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_449),
.A2(n_437),
.B1(n_436),
.B2(n_427),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_461),
.C(n_451),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_476),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_443),
.A2(n_438),
.B(n_439),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_450),
.A2(n_420),
.B1(n_425),
.B2(n_442),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_473),
.A2(n_460),
.B1(n_442),
.B2(n_456),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_446),
.B(n_425),
.Y(n_476)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_478),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_475),
.B(n_469),
.Y(n_479)
);

OAI21x1_ASAP7_75t_SL g490 ( 
.A1(n_479),
.A2(n_485),
.B(n_464),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_480),
.B(n_488),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_466),
.B(n_444),
.C(n_451),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_481),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_470),
.B(n_455),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_484),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_474),
.A2(n_457),
.B(n_448),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_466),
.B(n_458),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_467),
.Y(n_494)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_490),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_494),
.B(n_495),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_483),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_488),
.B(n_473),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_496),
.A2(n_486),
.B(n_479),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_497),
.B(n_489),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_491),
.A2(n_480),
.B(n_481),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_500),
.A2(n_493),
.B(n_492),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_501),
.B(n_502),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_498),
.B(n_489),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_503),
.B(n_499),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_504),
.A2(n_492),
.B(n_478),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_506),
.A2(n_505),
.B(n_477),
.Y(n_507)
);

BUFx24_ASAP7_75t_SL g508 ( 
.A(n_507),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_476),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_509),
.A2(n_471),
.B(n_494),
.Y(n_510)
);


endmodule