module fake_jpeg_1018_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_41),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_50),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_15),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

CKINVDCx9p33_ASAP7_75t_R g55 ( 
.A(n_32),
.Y(n_55)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_62),
.B1(n_27),
.B2(n_25),
.Y(n_95)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_22),
.B(n_0),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_20),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_20),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_64),
.B(n_72),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_38),
.A2(n_26),
.B1(n_37),
.B2(n_30),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_90),
.B1(n_91),
.B2(n_55),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_44),
.B(n_36),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_19),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_19),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_41),
.B(n_24),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_40),
.B(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_93),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_42),
.A2(n_28),
.B1(n_34),
.B2(n_30),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_59),
.A2(n_37),
.B1(n_34),
.B2(n_28),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_29),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_29),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_45),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_122),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_103),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_57),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_104),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_96),
.A2(n_58),
.B1(n_23),
.B2(n_25),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_43),
.C(n_46),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_94),
.C(n_76),
.Y(n_131)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_23),
.B1(n_27),
.B2(n_39),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_110),
.A2(n_113),
.B(n_115),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_78),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_74),
.A2(n_48),
.B1(n_61),
.B2(n_2),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_12),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_127),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_86),
.A2(n_48),
.B1(n_1),
.B2(n_4),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_7),
.B(n_8),
.Y(n_145)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_68),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_83),
.B1(n_77),
.B2(n_87),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_83),
.B1(n_77),
.B2(n_76),
.Y(n_132)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_125),
.Y(n_135)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_92),
.Y(n_130)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_64),
.B(n_11),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_67),
.B(n_94),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_145),
.B(n_120),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_141),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_108),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_133),
.B1(n_136),
.B2(n_147),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_100),
.A2(n_70),
.B1(n_87),
.B2(n_84),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_9),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_84),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_109),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_111),
.B(n_5),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_144),
.B(n_151),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_104),
.A2(n_8),
.B1(n_84),
.B2(n_126),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_104),
.A2(n_126),
.B1(n_117),
.B2(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_147),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_99),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_156),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_167),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_134),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_129),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_166),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_169),
.C(n_171),
.Y(n_174)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_151),
.B(n_111),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_163),
.B(n_165),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_144),
.B(n_112),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_148),
.A2(n_125),
.B1(n_123),
.B2(n_107),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_148),
.A2(n_112),
.B1(n_106),
.B2(n_114),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_122),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_140),
.B(n_124),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_170),
.B(n_146),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_131),
.C(n_150),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_139),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_173),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_138),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_162),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_177),
.Y(n_197)
);

OAI32xp33_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_142),
.A3(n_135),
.B1(n_136),
.B2(n_146),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_181),
.B(n_182),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_154),
.B(n_140),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_157),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_183),
.B(n_187),
.Y(n_196)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_167),
.B1(n_155),
.B2(n_159),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_190),
.A2(n_186),
.B1(n_180),
.B2(n_137),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_171),
.C(n_160),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_193),
.C(n_195),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_169),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_173),
.C(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_128),
.C(n_129),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_200),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_168),
.C(n_142),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_178),
.A2(n_168),
.B1(n_133),
.B2(n_132),
.Y(n_201)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

OA21x2_ASAP7_75t_SL g202 ( 
.A1(n_197),
.A2(n_185),
.B(n_178),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_203),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_SL g203 ( 
.A(n_192),
.B(n_175),
.C(n_189),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_200),
.A2(n_185),
.B(n_177),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_206),
.Y(n_215)
);

OAI322xp33_ASAP7_75t_L g205 ( 
.A1(n_195),
.A2(n_184),
.A3(n_186),
.B1(n_180),
.B2(n_145),
.C1(n_137),
.C2(n_133),
.Y(n_205)
);

NOR4xp25_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_196),
.C(n_199),
.D(n_204),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_194),
.Y(n_212)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_208),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_213),
.A2(n_210),
.B(n_206),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_191),
.C(n_193),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_209),
.Y(n_222)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_217),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_221),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_207),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_215),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_211),
.B1(n_210),
.B2(n_212),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_225),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_219),
.A2(n_203),
.B(n_222),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_226),
.B(n_219),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_223),
.B(n_227),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_221),
.Y(n_231)
);


endmodule