module fake_jpeg_13230_n_620 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_620);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_620;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_14),
.B(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_18),
.Y(n_60)
);

INVx5_ASAP7_75t_SL g202 ( 
.A(n_60),
.Y(n_202)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_62),
.B(n_69),
.Y(n_151)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_17),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_70),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_71),
.B(n_82),
.Y(n_129)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_72),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_74),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_75),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_76),
.Y(n_190)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_79),
.Y(n_191)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_80),
.Y(n_183)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_8),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_83),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g171 ( 
.A(n_85),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_18),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_87),
.B(n_88),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_17),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_28),
.B(n_31),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_89),
.B(n_92),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_91),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_28),
.B(n_31),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_95),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_35),
.Y(n_96)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_97),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_38),
.B(n_8),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_100),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_23),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_101),
.Y(n_178)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_102),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_23),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_112),
.Y(n_159)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_104),
.Y(n_140)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

BUFx10_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_107),
.Y(n_179)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_108),
.Y(n_205)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_109),
.Y(n_187)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

BUFx4f_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_38),
.B(n_8),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_115),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_49),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_114),
.A2(n_19),
.B1(n_54),
.B2(n_42),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_45),
.B(n_6),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_20),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_116),
.B(n_117),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_39),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_45),
.B(n_9),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g198 ( 
.A1(n_118),
.A2(n_13),
.B(n_11),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_35),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g199 ( 
.A(n_119),
.B(n_123),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_39),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_120),
.B(n_121),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_37),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_39),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_122),
.B(n_124),
.Y(n_181)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_37),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_70),
.A2(n_34),
.B1(n_47),
.B2(n_41),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_127),
.A2(n_162),
.B1(n_164),
.B2(n_192),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_66),
.A2(n_59),
.B1(n_49),
.B2(n_34),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_130),
.A2(n_147),
.B1(n_157),
.B2(n_203),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_79),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_133),
.B(n_154),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_65),
.A2(n_34),
.B1(n_47),
.B2(n_41),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_134),
.A2(n_156),
.B1(n_167),
.B2(n_170),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_68),
.B(n_24),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_136),
.B(n_152),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_80),
.A2(n_59),
.B1(n_49),
.B2(n_47),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_73),
.B(n_29),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_105),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_74),
.A2(n_47),
.B1(n_41),
.B2(n_37),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_64),
.A2(n_59),
.B1(n_41),
.B2(n_26),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_161),
.A2(n_177),
.B1(n_180),
.B2(n_188),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_75),
.A2(n_25),
.B1(n_29),
.B2(n_24),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_83),
.A2(n_25),
.B1(n_30),
.B2(n_46),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_84),
.B(n_30),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_165),
.B(n_168),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_90),
.A2(n_51),
.B1(n_50),
.B2(n_42),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_85),
.B(n_46),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_97),
.A2(n_50),
.B1(n_51),
.B2(n_19),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_98),
.A2(n_36),
.B1(n_44),
.B2(n_43),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_101),
.A2(n_44),
.B1(n_43),
.B2(n_32),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_117),
.B(n_26),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_186),
.B(n_196),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_111),
.A2(n_44),
.B1(n_43),
.B2(n_32),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_114),
.A2(n_32),
.B1(n_26),
.B2(n_54),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_107),
.A2(n_54),
.B1(n_58),
.B2(n_10),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_195),
.A2(n_4),
.B(n_199),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_117),
.B(n_15),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_120),
.B(n_14),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_197),
.B(n_126),
.Y(n_265)
);

OR2x2_ASAP7_75t_SL g222 ( 
.A(n_198),
.B(n_0),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_94),
.A2(n_58),
.B1(n_1),
.B2(n_2),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_201),
.A2(n_171),
.B1(n_182),
.B2(n_141),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_91),
.A2(n_58),
.B1(n_1),
.B2(n_2),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_93),
.A2(n_58),
.B1(n_1),
.B2(n_2),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_204),
.A2(n_86),
.B1(n_76),
.B2(n_119),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_151),
.B(n_96),
.C(n_122),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_206),
.B(n_219),
.C(n_242),
.Y(n_283)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_207),
.Y(n_306)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_128),
.Y(n_209)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_209),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_210),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_159),
.B(n_122),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_211),
.B(n_228),
.Y(n_299)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

INVx13_ASAP7_75t_L g335 ( 
.A(n_212),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_131),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_213),
.Y(n_320)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_215),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_143),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_216),
.B(n_236),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_144),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_217),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_150),
.B(n_87),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_220),
.Y(n_288)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_144),
.Y(n_221)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_221),
.Y(n_294)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_222),
.A2(n_265),
.B(n_266),
.Y(n_305)
);

OR2x4_ASAP7_75t_L g223 ( 
.A(n_150),
.B(n_202),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_223),
.B(n_245),
.Y(n_334)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_138),
.Y(n_225)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_225),
.Y(n_292)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_226),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_227),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_132),
.B(n_120),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_155),
.B(n_123),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_229),
.B(n_240),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_144),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_230),
.Y(n_329)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_231),
.Y(n_319)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_232),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_129),
.A2(n_60),
.B1(n_86),
.B2(n_76),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_233),
.A2(n_277),
.B1(n_278),
.B2(n_137),
.Y(n_289)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_235),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_144),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_237),
.Y(n_307)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_136),
.Y(n_239)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_239),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_173),
.B(n_0),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_150),
.B(n_0),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_241),
.B(n_244),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_158),
.B(n_1),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_176),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_243),
.B(n_256),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_152),
.B(n_165),
.Y(n_244)
);

OR2x4_ASAP7_75t_L g245 ( 
.A(n_155),
.B(n_5),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_125),
.Y(n_246)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_246),
.Y(n_313)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_146),
.Y(n_247)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_247),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_168),
.B(n_3),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_250),
.Y(n_298)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_187),
.Y(n_249)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_249),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_155),
.B(n_3),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_162),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_251),
.A2(n_171),
.B1(n_194),
.B2(n_172),
.Y(n_280)
);

OA22x2_ASAP7_75t_L g252 ( 
.A1(n_164),
.A2(n_3),
.B1(n_4),
.B2(n_127),
.Y(n_252)
);

AO22x1_ASAP7_75t_L g340 ( 
.A1(n_252),
.A2(n_264),
.B1(n_223),
.B2(n_236),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_253),
.A2(n_190),
.B(n_126),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_189),
.B(n_125),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_255),
.B(n_272),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_181),
.B(n_175),
.Y(n_256)
);

BUFx4f_ASAP7_75t_SL g257 ( 
.A(n_191),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_257),
.B(n_262),
.Y(n_337)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_146),
.Y(n_258)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_258),
.Y(n_318)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_189),
.Y(n_259)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_148),
.Y(n_260)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_260),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_160),
.B(n_179),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_261),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_148),
.B(n_163),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_160),
.B(n_179),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_263),
.Y(n_324)
);

OA22x2_ASAP7_75t_L g264 ( 
.A1(n_199),
.A2(n_201),
.B1(n_192),
.B2(n_163),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_139),
.B(n_140),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_139),
.B(n_140),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_267),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_131),
.Y(n_269)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_269),
.Y(n_331)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_200),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_270),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_177),
.A2(n_188),
.B1(n_134),
.B2(n_156),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_271),
.A2(n_274),
.B1(n_275),
.B2(n_279),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_195),
.B(n_169),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_139),
.B(n_140),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_273),
.Y(n_327)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_184),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_142),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_145),
.B(n_183),
.C(n_200),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_183),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_149),
.A2(n_194),
.B1(n_172),
.B2(n_135),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_142),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_L g351 ( 
.A1(n_280),
.A2(n_289),
.B1(n_274),
.B2(n_212),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_149),
.B1(n_135),
.B2(n_153),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_281),
.A2(n_303),
.B1(n_308),
.B2(n_336),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_285),
.A2(n_311),
.B(n_276),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_253),
.A2(n_137),
.B(n_145),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_286),
.A2(n_340),
.B(n_221),
.Y(n_363)
);

AND2x2_ASAP7_75t_SL g354 ( 
.A(n_296),
.B(n_237),
.Y(n_354)
);

OAI32xp33_ASAP7_75t_L g302 ( 
.A1(n_214),
.A2(n_141),
.A3(n_182),
.B1(n_174),
.B2(n_169),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_302),
.B(n_279),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_268),
.A2(n_153),
.B1(n_174),
.B2(n_184),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_214),
.B(n_184),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_304),
.B(n_325),
.C(n_298),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_239),
.A2(n_254),
.B1(n_224),
.B2(n_244),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_272),
.A2(n_224),
.B(n_219),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_206),
.B(n_241),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_234),
.A2(n_277),
.B1(n_264),
.B2(n_219),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_328),
.A2(n_333),
.B1(n_312),
.B2(n_324),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_248),
.B(n_250),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_338),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_234),
.A2(n_264),
.B1(n_254),
.B2(n_252),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_229),
.A2(n_208),
.B1(n_218),
.B2(n_264),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_242),
.B(n_255),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_242),
.B(n_222),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_259),
.Y(n_358)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_288),
.Y(n_341)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_341),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_308),
.B(n_262),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_342),
.B(n_350),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_343),
.A2(n_356),
.B(n_369),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_333),
.A2(n_252),
.B1(n_226),
.B2(n_220),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_344),
.A2(n_368),
.B1(n_295),
.B2(n_319),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_296),
.B(n_252),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_345),
.B(n_363),
.Y(n_422)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_288),
.Y(n_346)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_346),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_337),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_348),
.B(n_352),
.Y(n_405)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_349),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_297),
.B(n_238),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_351),
.A2(n_353),
.B1(n_359),
.B2(n_366),
.Y(n_394)
);

BUFx24_ASAP7_75t_SL g352 ( 
.A(n_290),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_328),
.A2(n_245),
.B1(n_270),
.B2(n_207),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_354),
.B(n_358),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_355),
.A2(n_357),
.B(n_329),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_323),
.A2(n_275),
.B(n_217),
.Y(n_356)
);

A2O1A1O1Ixp25_ASAP7_75t_L g357 ( 
.A1(n_311),
.A2(n_230),
.B(n_257),
.C(n_247),
.D(n_258),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_323),
.A2(n_231),
.B1(n_235),
.B2(n_215),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_293),
.Y(n_360)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_360),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_284),
.B(n_257),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_361),
.B(n_370),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_297),
.B(n_249),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_364),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_213),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_340),
.A2(n_309),
.B1(n_286),
.B2(n_289),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_317),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_367),
.B(n_373),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_309),
.A2(n_210),
.B1(n_269),
.B2(n_340),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_210),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_291),
.B(n_327),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_325),
.B(n_283),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_292),
.C(n_313),
.Y(n_389)
);

INVx6_ASAP7_75t_L g372 ( 
.A(n_320),
.Y(n_372)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_372),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_315),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_291),
.B(n_327),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_374),
.B(n_378),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_304),
.B(n_332),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_377),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_334),
.A2(n_326),
.B1(n_283),
.B2(n_280),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_376),
.A2(n_382),
.B1(n_386),
.B2(n_387),
.Y(n_424)
);

NOR3xp33_ASAP7_75t_SL g377 ( 
.A(n_339),
.B(n_298),
.C(n_305),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_299),
.B(n_300),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_335),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_379),
.B(n_295),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_314),
.B(n_324),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_380),
.B(n_383),
.Y(n_403)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_306),
.Y(n_381)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_381),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_287),
.B(n_300),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_306),
.Y(n_384)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_384),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_322),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_312),
.A2(n_302),
.B1(n_314),
.B2(n_285),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_287),
.A2(n_292),
.B1(n_330),
.B2(n_313),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_388),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_389),
.B(n_402),
.C(n_407),
.Y(n_445)
);

XOR2x2_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_330),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_390),
.B(n_414),
.Y(n_439)
);

AOI322xp5_ASAP7_75t_L g392 ( 
.A1(n_382),
.A2(n_321),
.A3(n_335),
.B1(n_320),
.B2(n_318),
.C1(n_331),
.C2(n_282),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_392),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_344),
.A2(n_331),
.B1(n_321),
.B2(n_318),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_393),
.A2(n_413),
.B1(n_341),
.B2(n_346),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_363),
.A2(n_307),
.B(n_316),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_399),
.A2(n_426),
.B(n_357),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_369),
.A2(n_307),
.B(n_316),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_401),
.A2(n_408),
.B(n_427),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_404),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_371),
.B(n_322),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_369),
.A2(n_301),
.B(n_310),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_347),
.B(n_301),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_411),
.B(n_415),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_383),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_406),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_385),
.B(n_375),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_347),
.B(n_310),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_350),
.B(n_319),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_416),
.B(n_370),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_362),
.B(n_294),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_367),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_343),
.A2(n_282),
.B(n_294),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_357),
.A2(n_345),
.B(n_355),
.Y(n_427)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_428),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_406),
.B(n_374),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_429),
.B(n_438),
.Y(n_464)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_430),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_404),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_432),
.B(n_446),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_379),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_433),
.B(n_435),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_373),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_395),
.Y(n_436)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_436),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_437),
.A2(n_449),
.B1(n_450),
.B2(n_460),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_380),
.Y(n_438)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_395),
.Y(n_440)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_440),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_414),
.B(n_354),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_461),
.C(n_445),
.Y(n_466)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_444),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_420),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_410),
.Y(n_447)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_447),
.Y(n_488)
);

CKINVDCx14_ASAP7_75t_R g448 ( 
.A(n_403),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_448),
.B(n_452),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_424),
.A2(n_365),
.B1(n_394),
.B2(n_399),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_424),
.A2(n_365),
.B1(n_368),
.B2(n_342),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_420),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_422),
.A2(n_356),
.B(n_345),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_453),
.B(n_454),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_396),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_455),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_425),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_458),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_393),
.A2(n_366),
.B1(n_386),
.B2(n_376),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_457),
.A2(n_463),
.B1(n_398),
.B2(n_426),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_403),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_417),
.Y(n_459)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_459),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_394),
.A2(n_345),
.B1(n_364),
.B2(n_348),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_407),
.B(n_354),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_391),
.B(n_361),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_391),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_451),
.A2(n_396),
.B1(n_411),
.B2(n_400),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_465),
.A2(n_472),
.B1(n_478),
.B2(n_485),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_466),
.B(n_468),
.C(n_469),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_439),
.B(n_445),
.C(n_441),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_445),
.B(n_402),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_436),
.Y(n_470)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_470),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_433),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_471),
.B(n_481),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_457),
.A2(n_400),
.B1(n_415),
.B2(n_427),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_439),
.B(n_390),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_483),
.C(n_487),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_439),
.B(n_390),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_434),
.A2(n_398),
.B1(n_388),
.B2(n_422),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_441),
.B(n_389),
.C(n_354),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_450),
.A2(n_413),
.B1(n_422),
.B2(n_353),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_491),
.A2(n_473),
.B1(n_463),
.B2(n_443),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_443),
.A2(n_422),
.B1(n_416),
.B2(n_392),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_492),
.A2(n_449),
.B1(n_460),
.B2(n_431),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_461),
.B(n_397),
.C(n_358),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_446),
.C(n_452),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_440),
.Y(n_495)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_495),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_494),
.B(n_437),
.Y(n_497)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_497),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_469),
.B(n_461),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_499),
.B(n_504),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_486),
.B(n_458),
.Y(n_501)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_501),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_502),
.A2(n_505),
.B1(n_512),
.B2(n_519),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_464),
.A2(n_435),
.B1(n_438),
.B2(n_448),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_503),
.A2(n_467),
.B1(n_477),
.B2(n_470),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_473),
.A2(n_437),
.B1(n_456),
.B2(n_463),
.Y(n_505)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_475),
.Y(n_509)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_509),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_510),
.A2(n_511),
.B1(n_477),
.B2(n_493),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_492),
.A2(n_449),
.B1(n_431),
.B2(n_432),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_491),
.A2(n_453),
.B1(n_430),
.B2(n_442),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_444),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_513),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_475),
.B(n_429),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_514),
.B(n_521),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_466),
.B(n_397),
.C(n_442),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_515),
.B(n_518),
.C(n_522),
.Y(n_532)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_474),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_516),
.B(n_520),
.Y(n_531)
);

A2O1A1Ixp33_ASAP7_75t_SL g517 ( 
.A1(n_484),
.A2(n_408),
.B(n_401),
.C(n_455),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_517),
.A2(n_485),
.B(n_495),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_468),
.B(n_397),
.C(n_459),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_484),
.A2(n_428),
.B1(n_462),
.B2(n_447),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_476),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_467),
.B(n_405),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_487),
.B(n_418),
.C(n_417),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_476),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_523),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_524),
.A2(n_512),
.B1(n_505),
.B2(n_502),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_499),
.B(n_479),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_526),
.B(n_498),
.Y(n_553)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_527),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_529),
.A2(n_497),
.B(n_513),
.Y(n_549)
);

BUFx12_ASAP7_75t_L g530 ( 
.A(n_511),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g559 ( 
.A(n_530),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_496),
.B(n_483),
.C(n_465),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_533),
.B(n_534),
.C(n_535),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_496),
.B(n_478),
.C(n_489),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_522),
.B(n_490),
.C(n_489),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_515),
.B(n_490),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_537),
.B(n_545),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_518),
.B(n_488),
.C(n_482),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_540),
.B(n_508),
.C(n_506),
.Y(n_566)
);

BUFx12f_ASAP7_75t_SL g541 ( 
.A(n_500),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_541),
.A2(n_544),
.B(n_510),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_SL g542 ( 
.A(n_519),
.B(n_488),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_542),
.B(n_513),
.Y(n_551)
);

BUFx12f_ASAP7_75t_SL g544 ( 
.A(n_497),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_504),
.B(n_482),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_549),
.A2(n_558),
.B(n_536),
.Y(n_578)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_550),
.Y(n_571)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_551),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_553),
.B(n_565),
.Y(n_576)
);

CKINVDCx16_ASAP7_75t_R g554 ( 
.A(n_531),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_554),
.B(n_555),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_540),
.B(n_405),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_538),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_556),
.B(n_562),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_543),
.B(n_378),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_557),
.B(n_560),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_547),
.B(n_507),
.Y(n_560)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_538),
.Y(n_562)
);

NOR2xp67_ASAP7_75t_SL g563 ( 
.A(n_528),
.B(n_498),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_563),
.A2(n_537),
.B(n_526),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_527),
.A2(n_546),
.B1(n_525),
.B2(n_539),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_564),
.A2(n_530),
.B1(n_517),
.B2(n_541),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_528),
.B(n_507),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_566),
.B(n_529),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_561),
.B(n_532),
.C(n_534),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_567),
.B(n_568),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_561),
.B(n_532),
.C(n_545),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_552),
.A2(n_525),
.B1(n_544),
.B2(n_533),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_570),
.A2(n_564),
.B1(n_550),
.B2(n_559),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_572),
.A2(n_566),
.B(n_549),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_565),
.B(n_535),
.C(n_536),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_573),
.B(n_577),
.C(n_581),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_575),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_548),
.B(n_553),
.C(n_552),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_SL g587 ( 
.A1(n_578),
.A2(n_517),
.B(n_556),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_548),
.B(n_517),
.C(n_530),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_558),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_582),
.A2(n_583),
.B1(n_581),
.B2(n_571),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_585),
.A2(n_589),
.B(n_590),
.Y(n_605)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_586),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_587),
.A2(n_592),
.B(n_359),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_582),
.A2(n_562),
.B(n_480),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_570),
.A2(n_480),
.B(n_419),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_SL g592 ( 
.A1(n_578),
.A2(n_418),
.B(n_349),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_567),
.B(n_419),
.C(n_421),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_593),
.B(n_595),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_594),
.B(n_596),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_574),
.A2(n_579),
.B1(n_580),
.B2(n_569),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_568),
.B(n_423),
.C(n_421),
.Y(n_596)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_598),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_588),
.A2(n_577),
.B(n_573),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_601),
.A2(n_587),
.B(n_592),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_591),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_602),
.B(n_603),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_584),
.B(n_576),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_591),
.B(n_576),
.Y(n_604)
);

AOI21xp33_ASAP7_75t_L g611 ( 
.A1(n_604),
.A2(n_377),
.B(n_372),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_606),
.A2(n_600),
.B(n_377),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_597),
.A2(n_599),
.B1(n_605),
.B2(n_604),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_608),
.B(n_611),
.Y(n_612)
);

AO21x1_ASAP7_75t_L g609 ( 
.A1(n_599),
.A2(n_423),
.B(n_360),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_609),
.Y(n_613)
);

NAND4xp25_ASAP7_75t_L g617 ( 
.A(n_614),
.B(n_615),
.C(n_387),
.D(n_372),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_607),
.B(n_610),
.Y(n_615)
);

BUFx24_ASAP7_75t_SL g616 ( 
.A(n_612),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_616),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_618),
.A2(n_613),
.B1(n_617),
.B2(n_381),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_619),
.B(n_384),
.Y(n_620)
);


endmodule