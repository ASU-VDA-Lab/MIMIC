module fake_ariane_1189_n_1107 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1107);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1107;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_1016;
wire n_346;
wire n_940;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_945;
wire n_702;
wire n_958;
wire n_905;
wire n_207;
wire n_898;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_779;
wire n_754;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_928;
wire n_839;
wire n_1099;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_658;
wire n_617;
wire n_616;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_772;
wire n_741;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_1081;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_664;
wire n_629;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_931;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1102;
wire n_975;
wire n_1101;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_484;
wire n_411;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_767;
wire n_736;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g206 ( 
.A(n_27),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_63),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_46),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_85),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_188),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_28),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_86),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_22),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_81),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_8),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_181),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_66),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_194),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_116),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_41),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_94),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_78),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_120),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_162),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_26),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_64),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_34),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_163),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_59),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_192),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_117),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_189),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_51),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_137),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_150),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_10),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_53),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_195),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_112),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_104),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_76),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_191),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_7),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_21),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_61),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_12),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_168),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_160),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_184),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_106),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_23),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_147),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_165),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_89),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_176),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_67),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_68),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_45),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_29),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_190),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_21),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_152),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_202),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_91),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_44),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_50),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_37),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_186),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_107),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_183),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_153),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_128),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_113),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_206),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_212),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_213),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_215),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_214),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_208),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_212),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_217),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_217),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_256),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_233),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_218),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_233),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_246),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_256),
.Y(n_292)
);

INVxp33_ASAP7_75t_SL g293 ( 
.A(n_253),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_254),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_224),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_230),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_234),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_235),
.Y(n_299)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_211),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_236),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_254),
.Y(n_303)
);

INVxp33_ASAP7_75t_SL g304 ( 
.A(n_269),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_237),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_241),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_258),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_258),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_264),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_242),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_226),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_247),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_251),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_260),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_271),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_257),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_273),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_275),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_257),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_264),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_207),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_209),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_210),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_285),
.Y(n_326)
);

AND2x6_ASAP7_75t_L g327 ( 
.A(n_289),
.B(n_216),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_289),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_219),
.Y(n_329)
);

OA21x2_ASAP7_75t_L g330 ( 
.A1(n_285),
.A2(n_287),
.B(n_286),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_277),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_286),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_301),
.B(n_226),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_293),
.A2(n_238),
.B1(n_248),
.B2(n_263),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_302),
.B(n_220),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_280),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_287),
.Y(n_337)
);

OAI21x1_ASAP7_75t_L g338 ( 
.A1(n_283),
.A2(n_222),
.B(n_221),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_325),
.B(n_268),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_293),
.A2(n_238),
.B1(n_248),
.B2(n_263),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_292),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_276),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_296),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_297),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_298),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_276),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_299),
.Y(n_349)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_324),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_279),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_304),
.A2(n_274),
.B1(n_267),
.B2(n_266),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_310),
.B(n_223),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_291),
.Y(n_355)
);

INVxp33_ASAP7_75t_SL g356 ( 
.A(n_324),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_304),
.B(n_225),
.Y(n_357)
);

OA21x2_ASAP7_75t_L g358 ( 
.A1(n_305),
.A2(n_228),
.B(n_227),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_306),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_295),
.B(n_323),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_281),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_312),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_313),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_314),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_300),
.B(n_229),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_316),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_323),
.B(n_231),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_320),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_317),
.B(n_232),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_321),
.Y(n_372)
);

INVxp33_ASAP7_75t_SL g373 ( 
.A(n_322),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_282),
.B(n_239),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_291),
.B(n_240),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_278),
.B(n_243),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_311),
.Y(n_377)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_278),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_290),
.B(n_244),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_290),
.Y(n_380)
);

NOR3xp33_ASAP7_75t_L g381 ( 
.A(n_378),
.B(n_288),
.C(n_284),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_330),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_330),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_330),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_326),
.Y(n_385)
);

INVx8_ASAP7_75t_L g386 ( 
.A(n_327),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_328),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_326),
.Y(n_388)
);

AO21x2_ASAP7_75t_L g389 ( 
.A1(n_338),
.A2(n_250),
.B(n_249),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_329),
.B(n_252),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_332),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_332),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_342),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

OR2x6_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_303),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_328),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_328),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_339),
.Y(n_398)
);

INVxp33_ASAP7_75t_SL g399 ( 
.A(n_369),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_342),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_329),
.B(n_255),
.Y(n_401)
);

NOR2x1p5_ASAP7_75t_L g402 ( 
.A(n_350),
.B(n_294),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_337),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_343),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_335),
.B(n_308),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_348),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_351),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_369),
.B(n_294),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_348),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_348),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_363),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_344),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_373),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_365),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_339),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

AND3x2_ASAP7_75t_L g418 ( 
.A(n_333),
.B(n_309),
.C(n_307),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_335),
.B(n_0),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_361),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_361),
.Y(n_423)
);

OAI22xp33_ASAP7_75t_L g424 ( 
.A1(n_334),
.A2(n_322),
.B1(n_309),
.B2(n_307),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_363),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_363),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_363),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_370),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_375),
.B(n_259),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_370),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_362),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_370),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_362),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_370),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_366),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_366),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_345),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_367),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_367),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_346),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_347),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_349),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_359),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_375),
.B(n_262),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_364),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_368),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_372),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_331),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_336),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_358),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_358),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_358),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_340),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_335),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_327),
.Y(n_455)
);

NOR2xp67_ASAP7_75t_L g456 ( 
.A(n_408),
.B(n_350),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_414),
.B(n_373),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_388),
.Y(n_458)
);

INVx4_ASAP7_75t_SL g459 ( 
.A(n_455),
.Y(n_459)
);

INVx4_ASAP7_75t_SL g460 ( 
.A(n_455),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_388),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_L g462 ( 
.A(n_454),
.B(n_360),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_387),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_406),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_392),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_406),
.B(n_355),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_393),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_395),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_393),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_419),
.Y(n_471)
);

BUFx5_ASAP7_75t_L g472 ( 
.A(n_451),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_419),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_442),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_442),
.Y(n_475)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_382),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_399),
.B(n_356),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_413),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_448),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_424),
.B(n_356),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_448),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_404),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_360),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_420),
.Y(n_484)
);

AND2x2_ASAP7_75t_SL g485 ( 
.A(n_420),
.B(n_341),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_395),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_404),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_395),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_418),
.B(n_379),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_405),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_453),
.B(n_377),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_405),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_415),
.B(n_329),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_435),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_435),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_436),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_409),
.B(n_380),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_413),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_436),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_386),
.B(n_327),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_438),
.Y(n_501)
);

INVxp33_ASAP7_75t_L g502 ( 
.A(n_420),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_395),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_438),
.Y(n_504)
);

AND2x2_ASAP7_75t_SL g505 ( 
.A(n_420),
.B(n_381),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_417),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_447),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_447),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_454),
.B(n_377),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_398),
.B(n_376),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_431),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_431),
.Y(n_512)
);

INVxp33_ASAP7_75t_L g513 ( 
.A(n_390),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_433),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_401),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_443),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_443),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_443),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_449),
.Y(n_520)
);

XOR2x2_ASAP7_75t_L g521 ( 
.A(n_429),
.B(n_379),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_417),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_449),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_449),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_440),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_382),
.B(n_327),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_440),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_395),
.B(n_379),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_441),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_417),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_386),
.B(n_327),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_444),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_385),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_451),
.B(n_353),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_385),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_437),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_445),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_445),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_483),
.A2(n_357),
.B1(n_371),
.B2(n_398),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_477),
.B(n_357),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_480),
.A2(n_374),
.B1(n_354),
.B2(n_371),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_474),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_483),
.B(n_416),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_462),
.B(n_456),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_516),
.B(n_484),
.Y(n_546)
);

NAND2x1p5_ASAP7_75t_L g547 ( 
.A(n_503),
.B(n_427),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_516),
.B(n_416),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_513),
.B(n_437),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_510),
.B(n_437),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_475),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_510),
.B(n_446),
.Y(n_552)
);

NOR3xp33_ASAP7_75t_L g553 ( 
.A(n_467),
.B(n_374),
.C(n_354),
.Y(n_553)
);

AND2x6_ASAP7_75t_L g554 ( 
.A(n_526),
.B(n_382),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_479),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_478),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_493),
.B(n_374),
.Y(n_557)
);

AOI221xp5_ASAP7_75t_L g558 ( 
.A1(n_457),
.A2(n_354),
.B1(n_446),
.B2(n_439),
.C(n_412),
.Y(n_558)
);

AND2x2_ASAP7_75t_SL g559 ( 
.A(n_485),
.B(n_386),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_L g560 ( 
.A(n_463),
.B(n_402),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_491),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_498),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_537),
.B(n_402),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_481),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_493),
.B(n_439),
.Y(n_565)
);

INVxp67_ASAP7_75t_SL g566 ( 
.A(n_476),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_509),
.B(n_439),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_502),
.B(n_427),
.Y(n_568)
);

NOR2x1p5_ASAP7_75t_L g569 ( 
.A(n_528),
.B(n_486),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_532),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_507),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_508),
.B(n_439),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_497),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_482),
.B(n_391),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_506),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_487),
.B(n_391),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_469),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_490),
.Y(n_578)
);

O2A1O1Ixp5_ASAP7_75t_L g579 ( 
.A1(n_492),
.A2(n_427),
.B(n_428),
.C(n_412),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_489),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_464),
.B(n_386),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_476),
.B(n_383),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_534),
.A2(n_452),
.B1(n_450),
.B2(n_386),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_488),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_502),
.B(n_427),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_511),
.B(n_383),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_464),
.B(n_428),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_525),
.A2(n_452),
.B1(n_450),
.B2(n_400),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_512),
.B(n_384),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_527),
.B(n_428),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_522),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_505),
.B(n_428),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_529),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_530),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_535),
.B(n_400),
.Y(n_595)
);

CKINVDCx11_ASAP7_75t_R g596 ( 
.A(n_463),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_538),
.B(n_421),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_539),
.B(n_421),
.Y(n_598)
);

INVx8_ASAP7_75t_L g599 ( 
.A(n_463),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_521),
.A2(n_412),
.B1(n_411),
.B2(n_434),
.Y(n_600)
);

A2O1A1Ixp33_ASAP7_75t_L g601 ( 
.A1(n_514),
.A2(n_452),
.B(n_450),
.C(n_412),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_515),
.B(n_411),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_458),
.B(n_384),
.Y(n_603)
);

INVx8_ASAP7_75t_L g604 ( 
.A(n_459),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_461),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_541),
.A2(n_465),
.B1(n_468),
.B2(n_466),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_586),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_544),
.B(n_470),
.Y(n_608)
);

A2O1A1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_540),
.A2(n_518),
.B(n_519),
.C(n_517),
.Y(n_609)
);

OR2x6_ASAP7_75t_L g610 ( 
.A(n_604),
.B(n_471),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_543),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_542),
.B(n_473),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_557),
.B(n_520),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_551),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_596),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_569),
.B(n_459),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_570),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_556),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_549),
.B(n_472),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_555),
.Y(n_620)
);

NOR2xp67_ASAP7_75t_L g621 ( 
.A(n_573),
.B(n_523),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_564),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_584),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_553),
.A2(n_524),
.B1(n_531),
.B2(n_500),
.Y(n_624)
);

NOR3xp33_ASAP7_75t_SL g625 ( 
.A(n_545),
.B(n_265),
.C(n_389),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_604),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_587),
.A2(n_531),
.B1(n_500),
.B2(n_432),
.Y(n_627)
);

BUFx12f_ASAP7_75t_L g628 ( 
.A(n_563),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_561),
.B(n_422),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_604),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_563),
.B(n_422),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_599),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_599),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_571),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_599),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_586),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_577),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_587),
.B(n_459),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_590),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_578),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_581),
.B(n_460),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_581),
.B(n_460),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_552),
.B(n_494),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_580),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_605),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_548),
.B(n_423),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_593),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_546),
.B(n_495),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_558),
.B(n_423),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g650 ( 
.A(n_566),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_559),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_574),
.Y(n_652)
);

OR2x6_ASAP7_75t_L g653 ( 
.A(n_581),
.B(n_425),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_550),
.B(n_496),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_547),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_590),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_562),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_600),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_565),
.B(n_499),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_575),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_576),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_SL g662 ( 
.A(n_592),
.B(n_389),
.C(n_501),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_590),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_589),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_568),
.B(n_460),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_591),
.Y(n_666)
);

AO21x1_ASAP7_75t_L g667 ( 
.A1(n_612),
.A2(n_602),
.B(n_589),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_609),
.A2(n_601),
.B(n_579),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_641),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_611),
.Y(n_670)
);

A2O1A1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_606),
.A2(n_560),
.B(n_567),
.C(n_572),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_658),
.B(n_582),
.Y(n_672)
);

AOI21x1_ASAP7_75t_L g673 ( 
.A1(n_619),
.A2(n_597),
.B(n_595),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_654),
.A2(n_603),
.B(n_598),
.Y(n_674)
);

OAI21x1_ASAP7_75t_L g675 ( 
.A1(n_624),
.A2(n_603),
.B(n_582),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_608),
.B(n_547),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g677 ( 
.A1(n_659),
.A2(n_613),
.B(n_643),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_631),
.B(n_594),
.Y(n_678)
);

AO31x2_ASAP7_75t_L g679 ( 
.A1(n_607),
.A2(n_526),
.A3(n_504),
.B(n_533),
.Y(n_679)
);

NOR2xp67_ASAP7_75t_SL g680 ( 
.A(n_626),
.B(n_628),
.Y(n_680)
);

OAI21x1_ASAP7_75t_L g681 ( 
.A1(n_607),
.A2(n_588),
.B(n_536),
.Y(n_681)
);

OAI22x1_ASAP7_75t_L g682 ( 
.A1(n_663),
.A2(n_585),
.B1(n_426),
.B2(n_425),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_650),
.A2(n_583),
.B(n_389),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_652),
.B(n_426),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_626),
.Y(n_685)
);

AND2x6_ASAP7_75t_SL g686 ( 
.A(n_610),
.B(n_0),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_636),
.A2(n_472),
.B(n_410),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_641),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_636),
.A2(n_664),
.B(n_627),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_614),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_661),
.B(n_430),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_642),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_620),
.B(n_430),
.Y(n_693)
);

OAI21x1_ASAP7_75t_L g694 ( 
.A1(n_664),
.A2(n_434),
.B(n_397),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_610),
.A2(n_410),
.B1(n_407),
.B2(n_403),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_656),
.B(n_472),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_632),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_622),
.B(n_407),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_618),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_634),
.Y(n_700)
);

AO31x2_ASAP7_75t_L g701 ( 
.A1(n_657),
.A2(n_397),
.A3(n_403),
.B(n_410),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_638),
.A2(n_472),
.B(n_407),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_648),
.A2(n_397),
.B(n_432),
.C(n_396),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_638),
.A2(n_653),
.B(n_656),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_644),
.B(n_432),
.Y(n_705)
);

OAI21x1_ASAP7_75t_L g706 ( 
.A1(n_647),
.A2(n_472),
.B(n_554),
.Y(n_706)
);

AOI21x1_ASAP7_75t_SL g707 ( 
.A1(n_665),
.A2(n_1),
.B(n_2),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_640),
.B(n_645),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_615),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_666),
.Y(n_710)
);

OAI21x1_ASAP7_75t_L g711 ( 
.A1(n_630),
.A2(n_646),
.B(n_649),
.Y(n_711)
);

OAI21x1_ASAP7_75t_SL g712 ( 
.A1(n_639),
.A2(n_554),
.B(n_432),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_623),
.B(n_554),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_617),
.Y(n_714)
);

AOI21xp33_ASAP7_75t_L g715 ( 
.A1(n_629),
.A2(n_432),
.B(n_394),
.Y(n_715)
);

A2O1A1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_625),
.A2(n_432),
.B(n_396),
.C(n_394),
.Y(n_716)
);

OAI21x1_ASAP7_75t_L g717 ( 
.A1(n_630),
.A2(n_554),
.B(n_394),
.Y(n_717)
);

OAI21x1_ASAP7_75t_L g718 ( 
.A1(n_660),
.A2(n_394),
.B(n_387),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_662),
.A2(n_396),
.B(n_394),
.C(n_387),
.Y(n_719)
);

AOI221xp5_ASAP7_75t_L g720 ( 
.A1(n_637),
.A2(n_396),
.B1(n_394),
.B2(n_387),
.C(n_4),
.Y(n_720)
);

OAI21xp5_ASAP7_75t_L g721 ( 
.A1(n_665),
.A2(n_396),
.B(n_387),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_621),
.B(n_387),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_655),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_616),
.B(n_1),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_714),
.Y(n_725)
);

A2O1A1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_683),
.A2(n_651),
.B(n_616),
.C(n_642),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_677),
.A2(n_656),
.B(n_653),
.Y(n_727)
);

OAI22x1_ASAP7_75t_L g728 ( 
.A1(n_670),
.A2(n_639),
.B1(n_626),
.B2(n_635),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_672),
.B(n_655),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_708),
.B(n_655),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_705),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_677),
.B(n_632),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_674),
.A2(n_635),
.B(n_396),
.Y(n_733)
);

A2O1A1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_720),
.A2(n_633),
.B(n_632),
.C(n_4),
.Y(n_734)
);

AO31x2_ASAP7_75t_L g735 ( 
.A1(n_667),
.A2(n_111),
.A3(n_205),
.B(n_204),
.Y(n_735)
);

OAI22xp33_ASAP7_75t_L g736 ( 
.A1(n_713),
.A2(n_633),
.B1(n_3),
.B2(n_5),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_686),
.B(n_633),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_706),
.A2(n_35),
.B(n_33),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_674),
.A2(n_2),
.B(n_3),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_697),
.Y(n_740)
);

O2A1O1Ixp33_ASAP7_75t_SL g741 ( 
.A1(n_671),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_676),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_687),
.A2(n_668),
.B(n_719),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_690),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_716),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_668),
.A2(n_11),
.B(n_12),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_700),
.Y(n_747)
);

O2A1O1Ixp33_ASAP7_75t_SL g748 ( 
.A1(n_696),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_678),
.Y(n_749)
);

AO31x2_ASAP7_75t_L g750 ( 
.A1(n_682),
.A2(n_121),
.A3(n_203),
.B(n_201),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_689),
.A2(n_13),
.B(n_14),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_697),
.Y(n_752)
);

O2A1O1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_703),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_753)
);

AO31x2_ASAP7_75t_L g754 ( 
.A1(n_710),
.A2(n_122),
.A3(n_200),
.B(n_199),
.Y(n_754)
);

AO31x2_ASAP7_75t_L g755 ( 
.A1(n_699),
.A2(n_118),
.A3(n_198),
.B(n_197),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_702),
.A2(n_16),
.B(n_17),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_675),
.A2(n_18),
.B(n_19),
.Y(n_757)
);

NAND3x1_ASAP7_75t_L g758 ( 
.A(n_724),
.B(n_18),
.C(n_19),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_723),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_L g760 ( 
.A(n_697),
.B(n_20),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_L g761 ( 
.A(n_685),
.B(n_36),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_721),
.A2(n_20),
.B(n_22),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_686),
.B(n_23),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_695),
.B(n_24),
.Y(n_764)
);

OAI21xp5_ASAP7_75t_L g765 ( 
.A1(n_711),
.A2(n_24),
.B(n_25),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_698),
.Y(n_766)
);

O2A1O1Ixp33_ASAP7_75t_SL g767 ( 
.A1(n_722),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_693),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_721),
.A2(n_28),
.B(n_29),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_669),
.B(n_30),
.Y(n_770)
);

OA21x2_ASAP7_75t_L g771 ( 
.A1(n_694),
.A2(n_130),
.B(n_196),
.Y(n_771)
);

AOI211x1_ASAP7_75t_L g772 ( 
.A1(n_680),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_717),
.A2(n_31),
.B(n_32),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_SL g774 ( 
.A1(n_684),
.A2(n_691),
.B(n_704),
.C(n_715),
.Y(n_774)
);

OAI22xp33_ASAP7_75t_L g775 ( 
.A1(n_669),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_775)
);

AOI221x1_ASAP7_75t_L g776 ( 
.A1(n_712),
.A2(n_42),
.B1(n_43),
.B2(n_47),
.C(n_48),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_718),
.A2(n_681),
.B(n_688),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_673),
.A2(n_49),
.B(n_52),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_688),
.A2(n_692),
.B(n_685),
.Y(n_779)
);

O2A1O1Ixp33_ASAP7_75t_SL g780 ( 
.A1(n_707),
.A2(n_54),
.B(n_55),
.C(n_56),
.Y(n_780)
);

AO31x2_ASAP7_75t_L g781 ( 
.A1(n_679),
.A2(n_57),
.A3(n_58),
.B(n_60),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_692),
.A2(n_62),
.B(n_65),
.C(n_69),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_SL g783 ( 
.A1(n_709),
.A2(n_70),
.B(n_71),
.C(n_72),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_679),
.A2(n_73),
.B(n_74),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_679),
.A2(n_75),
.B(n_77),
.Y(n_785)
);

OAI21x1_ASAP7_75t_L g786 ( 
.A1(n_701),
.A2(n_79),
.B(n_80),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_701),
.A2(n_82),
.B(n_83),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_744),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_763),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_789)
);

BUFx12f_ASAP7_75t_L g790 ( 
.A(n_740),
.Y(n_790)
);

INVx6_ASAP7_75t_L g791 ( 
.A(n_740),
.Y(n_791)
);

OAI22xp33_ASAP7_75t_L g792 ( 
.A1(n_742),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_731),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_746),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_752),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_759),
.Y(n_796)
);

CKINVDCx11_ASAP7_75t_R g797 ( 
.A(n_752),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_749),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_747),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_739),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_725),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_734),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_768),
.Y(n_803)
);

CKINVDCx11_ASAP7_75t_R g804 ( 
.A(n_766),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_729),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_730),
.Y(n_806)
);

BUFx2_ASAP7_75t_SL g807 ( 
.A(n_761),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_737),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_L g809 ( 
.A1(n_732),
.A2(n_110),
.B1(n_114),
.B2(n_115),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_SL g810 ( 
.A1(n_772),
.A2(n_119),
.B1(n_124),
.B2(n_125),
.Y(n_810)
);

OAI22xp33_ASAP7_75t_L g811 ( 
.A1(n_762),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_811)
);

CKINVDCx6p67_ASAP7_75t_R g812 ( 
.A(n_728),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_727),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_770),
.B(n_131),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_SL g815 ( 
.A1(n_778),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_815)
);

NAND2x1p5_ASAP7_75t_L g816 ( 
.A(n_779),
.B(n_135),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_781),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_781),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_754),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_SL g820 ( 
.A1(n_765),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_820)
);

INVx6_ASAP7_75t_L g821 ( 
.A(n_760),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_738),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_733),
.Y(n_823)
);

BUFx10_ASAP7_75t_L g824 ( 
.A(n_758),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_767),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_745),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_SL g827 ( 
.A1(n_751),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_777),
.Y(n_828)
);

BUFx2_ASAP7_75t_SL g829 ( 
.A(n_764),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_755),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_771),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_735),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_726),
.B(n_146),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_769),
.Y(n_834)
);

CKINVDCx6p67_ASAP7_75t_R g835 ( 
.A(n_783),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_735),
.B(n_148),
.Y(n_836)
);

INVx4_ASAP7_75t_L g837 ( 
.A(n_771),
.Y(n_837)
);

CKINVDCx11_ASAP7_75t_R g838 ( 
.A(n_736),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_756),
.A2(n_149),
.B1(n_151),
.B2(n_154),
.Y(n_839)
);

CKINVDCx11_ASAP7_75t_R g840 ( 
.A(n_741),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_755),
.Y(n_841)
);

BUFx2_ASAP7_75t_L g842 ( 
.A(n_750),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_774),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_750),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_757),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_797),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_799),
.Y(n_847)
);

BUFx2_ASAP7_75t_SL g848 ( 
.A(n_834),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_788),
.B(n_743),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_801),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_796),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_812),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_793),
.B(n_748),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_803),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_817),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_818),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_806),
.B(n_785),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_828),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_805),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_844),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_831),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_830),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_819),
.Y(n_863)
);

AOI222xp33_ASAP7_75t_L g864 ( 
.A1(n_838),
.A2(n_775),
.B1(n_782),
.B2(n_753),
.C1(n_786),
.C2(n_780),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_831),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_845),
.Y(n_866)
);

OAI21x1_ASAP7_75t_L g867 ( 
.A1(n_843),
.A2(n_784),
.B(n_787),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_823),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_823),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_813),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_813),
.B(n_776),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_791),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_816),
.A2(n_773),
.B(n_156),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_837),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_842),
.Y(n_875)
);

NAND2x1p5_ASAP7_75t_L g876 ( 
.A(n_841),
.B(n_155),
.Y(n_876)
);

BUFx2_ASAP7_75t_SL g877 ( 
.A(n_795),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_832),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_837),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_822),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_822),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_822),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_816),
.A2(n_157),
.B(n_158),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_836),
.Y(n_884)
);

INVx4_ASAP7_75t_L g885 ( 
.A(n_835),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_825),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_795),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_804),
.B(n_159),
.Y(n_888)
);

INVxp67_ASAP7_75t_SL g889 ( 
.A(n_833),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_795),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_847),
.Y(n_891)
);

OA21x2_ASAP7_75t_L g892 ( 
.A1(n_879),
.A2(n_865),
.B(n_870),
.Y(n_892)
);

OR2x6_ASAP7_75t_L g893 ( 
.A(n_884),
.B(n_807),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_868),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_861),
.Y(n_895)
);

AO21x1_ASAP7_75t_SL g896 ( 
.A1(n_879),
.A2(n_794),
.B(n_814),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_851),
.B(n_868),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_851),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_858),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_887),
.Y(n_900)
);

AOI221xp5_ASAP7_75t_L g901 ( 
.A1(n_870),
.A2(n_810),
.B1(n_800),
.B2(n_820),
.C(n_826),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_849),
.B(n_808),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_858),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_847),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_858),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_862),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_869),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_869),
.B(n_849),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_862),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_866),
.B(n_791),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_850),
.Y(n_911)
);

OR2x6_ASAP7_75t_L g912 ( 
.A(n_884),
.B(n_821),
.Y(n_912)
);

AO21x2_ASAP7_75t_L g913 ( 
.A1(n_871),
.A2(n_800),
.B(n_811),
.Y(n_913)
);

AO21x2_ASAP7_75t_L g914 ( 
.A1(n_871),
.A2(n_826),
.B(n_792),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_854),
.B(n_829),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_855),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_861),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_854),
.B(n_810),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_859),
.B(n_821),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_859),
.B(n_820),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_907),
.B(n_889),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_R g922 ( 
.A(n_911),
.B(n_846),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_894),
.Y(n_923)
);

NAND3xp33_ASAP7_75t_SL g924 ( 
.A(n_901),
.B(n_920),
.C(n_918),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_893),
.B(n_861),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_894),
.B(n_848),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_897),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_906),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_902),
.B(n_848),
.Y(n_929)
);

AOI21xp33_ASAP7_75t_L g930 ( 
.A1(n_914),
.A2(n_853),
.B(n_886),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_SL g931 ( 
.A1(n_914),
.A2(n_824),
.B1(n_884),
.B2(n_871),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_906),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_902),
.B(n_865),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_908),
.B(n_865),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_906),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_897),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_909),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_908),
.B(n_871),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_898),
.B(n_861),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_898),
.B(n_874),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_899),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_914),
.A2(n_840),
.B1(n_864),
.B2(n_824),
.Y(n_942)
);

AO21x2_ASAP7_75t_L g943 ( 
.A1(n_913),
.A2(n_882),
.B(n_863),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_941),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_923),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_941),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_926),
.B(n_910),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_926),
.B(n_910),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_928),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_934),
.B(n_915),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_928),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_924),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_934),
.B(n_915),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_929),
.B(n_913),
.Y(n_954)
);

NAND2x1p5_ASAP7_75t_SL g955 ( 
.A(n_927),
.B(n_888),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_927),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_941),
.Y(n_957)
);

AO21x2_ASAP7_75t_L g958 ( 
.A1(n_930),
.A2(n_914),
.B(n_913),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_932),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_950),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_954),
.B(n_930),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_945),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_955),
.B(n_936),
.Y(n_963)
);

OR2x2_ASAP7_75t_L g964 ( 
.A(n_955),
.B(n_936),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_947),
.B(n_929),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_950),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_951),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_953),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_947),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_953),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_956),
.B(n_938),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_948),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_965),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_962),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_972),
.B(n_960),
.Y(n_975)
);

INVxp67_ASAP7_75t_L g976 ( 
.A(n_962),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_969),
.B(n_948),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_971),
.B(n_952),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_967),
.Y(n_979)
);

OR2x6_ASAP7_75t_L g980 ( 
.A(n_963),
.B(n_888),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_978),
.B(n_954),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_974),
.B(n_966),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_976),
.B(n_968),
.Y(n_983)
);

OAI221xp5_ASAP7_75t_L g984 ( 
.A1(n_980),
.A2(n_961),
.B1(n_942),
.B2(n_931),
.C(n_964),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_973),
.B(n_970),
.Y(n_985)
);

NOR2x1_ASAP7_75t_L g986 ( 
.A(n_980),
.B(n_945),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_977),
.B(n_956),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_982),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_983),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_986),
.B(n_975),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_987),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_981),
.B(n_979),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_SL g993 ( 
.A1(n_984),
.A2(n_961),
.B1(n_958),
.B2(n_913),
.Y(n_993)
);

CKINVDCx16_ASAP7_75t_R g994 ( 
.A(n_985),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_982),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_986),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_982),
.B(n_967),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_982),
.Y(n_998)
);

INVx1_ASAP7_75t_SL g999 ( 
.A(n_994),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_997),
.Y(n_1000)
);

INVxp67_ASAP7_75t_L g1001 ( 
.A(n_996),
.Y(n_1001)
);

OAI211xp5_ASAP7_75t_SL g1002 ( 
.A1(n_995),
.A2(n_918),
.B(n_921),
.C(n_920),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_990),
.B(n_922),
.Y(n_1003)
);

INVxp67_ASAP7_75t_SL g1004 ( 
.A(n_990),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_993),
.A2(n_919),
.B(n_885),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_988),
.A2(n_958),
.B1(n_896),
.B2(n_943),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_991),
.A2(n_885),
.B1(n_852),
.B2(n_951),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_1005),
.A2(n_992),
.B(n_997),
.C(n_998),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_999),
.B(n_989),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_1004),
.B(n_958),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_1001),
.A2(n_919),
.B(n_885),
.Y(n_1011)
);

OAI32xp33_ASAP7_75t_L g1012 ( 
.A1(n_1002),
.A2(n_885),
.A3(n_852),
.B1(n_949),
.B2(n_959),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_1003),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_R g1014 ( 
.A(n_1000),
.B(n_852),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1007),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1006),
.Y(n_1016)
);

AOI221x1_ASAP7_75t_L g1017 ( 
.A1(n_1013),
.A2(n_802),
.B1(n_946),
.B2(n_944),
.C(n_957),
.Y(n_1017)
);

AOI221xp5_ASAP7_75t_L g1018 ( 
.A1(n_1016),
.A2(n_1008),
.B1(n_1012),
.B2(n_1010),
.C(n_1014),
.Y(n_1018)
);

AOI222xp33_ASAP7_75t_L g1019 ( 
.A1(n_1015),
.A2(n_957),
.B1(n_946),
.B2(n_944),
.C1(n_875),
.C2(n_878),
.Y(n_1019)
);

OAI221xp5_ASAP7_75t_L g1020 ( 
.A1(n_1009),
.A2(n_876),
.B1(n_815),
.B2(n_827),
.C(n_893),
.Y(n_1020)
);

OAI311xp33_ASAP7_75t_L g1021 ( 
.A1(n_1011),
.A2(n_789),
.A3(n_798),
.B1(n_839),
.C1(n_933),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_1008),
.A2(n_943),
.B(n_872),
.Y(n_1022)
);

OAI221xp5_ASAP7_75t_L g1023 ( 
.A1(n_1016),
.A2(n_876),
.B1(n_893),
.B2(n_896),
.C(n_872),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1013),
.B(n_943),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1024),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1019),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1017),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_1023),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_1018),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1020),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1021),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1022),
.Y(n_1032)
);

NAND2x1_ASAP7_75t_SL g1033 ( 
.A(n_1027),
.B(n_939),
.Y(n_1033)
);

NAND3xp33_ASAP7_75t_L g1034 ( 
.A(n_1029),
.B(n_809),
.C(n_886),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_1029),
.A2(n_883),
.B(n_873),
.Y(n_1035)
);

NAND3xp33_ASAP7_75t_SL g1036 ( 
.A(n_1031),
.B(n_876),
.C(n_933),
.Y(n_1036)
);

NAND4xp25_ASAP7_75t_L g1037 ( 
.A(n_1030),
.B(n_925),
.C(n_940),
.D(n_939),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_1032),
.B(n_925),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1026),
.Y(n_1039)
);

NOR4xp25_ASAP7_75t_L g1040 ( 
.A(n_1039),
.B(n_1025),
.C(n_1028),
.D(n_937),
.Y(n_1040)
);

NAND3xp33_ASAP7_75t_L g1041 ( 
.A(n_1034),
.B(n_892),
.C(n_937),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1033),
.B(n_932),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_1035),
.B(n_790),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_1038),
.A2(n_893),
.B(n_935),
.C(n_892),
.Y(n_1044)
);

OAI221xp5_ASAP7_75t_L g1045 ( 
.A1(n_1037),
.A2(n_893),
.B1(n_892),
.B2(n_935),
.C(n_882),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_1043),
.Y(n_1046)
);

NOR2x1_ASAP7_75t_L g1047 ( 
.A(n_1042),
.B(n_1036),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_L g1048 ( 
.A(n_1040),
.B(n_892),
.C(n_904),
.Y(n_1048)
);

NOR2x1_ASAP7_75t_L g1049 ( 
.A(n_1041),
.B(n_1045),
.Y(n_1049)
);

NAND5xp2_ASAP7_75t_L g1050 ( 
.A(n_1044),
.B(n_940),
.C(n_878),
.D(n_875),
.E(n_883),
.Y(n_1050)
);

NOR4xp25_ASAP7_75t_L g1051 ( 
.A(n_1043),
.B(n_916),
.C(n_891),
.D(n_904),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_1043),
.B(n_887),
.Y(n_1052)
);

NAND4xp25_ASAP7_75t_L g1053 ( 
.A(n_1043),
.B(n_925),
.C(n_917),
.D(n_895),
.Y(n_1053)
);

NAND4xp25_ASAP7_75t_L g1054 ( 
.A(n_1043),
.B(n_925),
.C(n_917),
.D(n_895),
.Y(n_1054)
);

NAND4xp75_ASAP7_75t_L g1055 ( 
.A(n_1047),
.B(n_900),
.C(n_891),
.D(n_887),
.Y(n_1055)
);

NOR3xp33_ASAP7_75t_L g1056 ( 
.A(n_1046),
.B(n_1049),
.C(n_1052),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1048),
.Y(n_1057)
);

AND3x4_ASAP7_75t_L g1058 ( 
.A(n_1051),
.B(n_890),
.C(n_877),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1054),
.B(n_900),
.Y(n_1059)
);

NOR4xp75_ASAP7_75t_SL g1060 ( 
.A(n_1053),
.B(n_917),
.C(n_895),
.D(n_874),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_1050),
.B(n_916),
.Y(n_1061)
);

NOR4xp25_ASAP7_75t_L g1062 ( 
.A(n_1046),
.B(n_890),
.C(n_909),
.D(n_881),
.Y(n_1062)
);

OAI211xp5_ASAP7_75t_SL g1063 ( 
.A1(n_1046),
.A2(n_874),
.B(n_895),
.C(n_917),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_1056),
.B(n_874),
.Y(n_1064)
);

NOR2xp67_ASAP7_75t_L g1065 ( 
.A(n_1057),
.B(n_161),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1058),
.Y(n_1066)
);

OAI221xp5_ASAP7_75t_L g1067 ( 
.A1(n_1061),
.A2(n_877),
.B1(n_912),
.B2(n_881),
.C(n_880),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_1055),
.B(n_880),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1059),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_1063),
.B(n_873),
.Y(n_1070)
);

NOR3xp33_ASAP7_75t_L g1071 ( 
.A(n_1060),
.B(n_867),
.C(n_166),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_1062),
.B(n_912),
.Y(n_1072)
);

NOR2xp67_ASAP7_75t_L g1073 ( 
.A(n_1057),
.B(n_164),
.Y(n_1073)
);

AND3x4_ASAP7_75t_L g1074 ( 
.A(n_1056),
.B(n_909),
.C(n_905),
.Y(n_1074)
);

NOR3xp33_ASAP7_75t_L g1075 ( 
.A(n_1056),
.B(n_867),
.C(n_169),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_SL g1076 ( 
.A(n_1055),
.B(n_167),
.C(n_170),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1066),
.A2(n_912),
.B1(n_857),
.B2(n_903),
.Y(n_1077)
);

XNOR2x1_ASAP7_75t_L g1078 ( 
.A(n_1065),
.B(n_1073),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_1069),
.Y(n_1079)
);

NAND2xp33_ASAP7_75t_SL g1080 ( 
.A(n_1076),
.B(n_1064),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1074),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_1072),
.B(n_171),
.Y(n_1082)
);

NOR2xp67_ASAP7_75t_L g1083 ( 
.A(n_1067),
.B(n_172),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1068),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1079),
.A2(n_1075),
.B1(n_1071),
.B2(n_1070),
.Y(n_1085)
);

OAI22x1_ASAP7_75t_L g1086 ( 
.A1(n_1084),
.A2(n_863),
.B1(n_860),
.B2(n_899),
.Y(n_1086)
);

AO22x2_ASAP7_75t_L g1087 ( 
.A1(n_1078),
.A2(n_860),
.B1(n_903),
.B2(n_899),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1082),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1081),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1080),
.Y(n_1090)
);

NAND2xp33_ASAP7_75t_SL g1091 ( 
.A(n_1090),
.B(n_1083),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1088),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1085),
.B(n_1077),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1092),
.B(n_1089),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1094),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1095),
.A2(n_1093),
.B1(n_1091),
.B2(n_1087),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1095),
.A2(n_1086),
.B1(n_905),
.B2(n_903),
.Y(n_1097)
);

OA22x2_ASAP7_75t_L g1098 ( 
.A1(n_1096),
.A2(n_912),
.B1(n_174),
.B2(n_175),
.Y(n_1098)
);

OAI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1097),
.A2(n_912),
.B1(n_857),
.B2(n_905),
.Y(n_1099)
);

OAI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_1096),
.A2(n_856),
.B1(n_855),
.B2(n_178),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1100),
.B(n_173),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1098),
.B(n_177),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1099),
.Y(n_1103)
);

OA21x2_ASAP7_75t_L g1104 ( 
.A1(n_1103),
.A2(n_1102),
.B(n_1101),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1102),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1105),
.A2(n_179),
.B1(n_180),
.B2(n_182),
.Y(n_1106)
);

AOI211xp5_ASAP7_75t_L g1107 ( 
.A1(n_1106),
.A2(n_1104),
.B(n_185),
.C(n_187),
.Y(n_1107)
);


endmodule