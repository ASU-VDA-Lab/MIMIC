module fake_jpeg_1431_n_217 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_217);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_10),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_31),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_82),
.Y(n_95)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_84),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_91),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_56),
.B1(n_64),
.B2(n_66),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_90),
.B1(n_85),
.B2(n_78),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_64),
.B1(n_56),
.B2(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_84),
.B(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_57),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_53),
.B1(n_54),
.B2(n_72),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_54),
.B1(n_80),
.B2(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_73),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_4),
.Y(n_136)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_94),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_63),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_68),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_95),
.A2(n_80),
.B1(n_84),
.B2(n_71),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_109),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_110),
.B(n_116),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_75),
.B(n_61),
.C(n_69),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_112),
.B(n_3),
.C(n_4),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_85),
.B(n_61),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_119),
.B1(n_98),
.B2(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_70),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_104),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_92),
.A2(n_59),
.B1(n_72),
.B2(n_55),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_86),
.B1(n_94),
.B2(n_99),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_138),
.B1(n_8),
.B2(n_9),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_16),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_135),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_98),
.B1(n_1),
.B2(n_2),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_130),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_27),
.B(n_50),
.C(n_47),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_139),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_141),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_6),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_135),
.B(n_107),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_142),
.B(n_159),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_112),
.B(n_111),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_153),
.B(n_35),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_136),
.A2(n_105),
.B1(n_103),
.B2(n_10),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_164),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_26),
.C(n_46),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_150),
.C(n_155),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_25),
.C(n_45),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_152),
.B(n_29),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_11),
.B(n_12),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_11),
.Y(n_154)
);

AO21x1_ASAP7_75t_L g178 ( 
.A1(n_154),
.A2(n_160),
.B(n_33),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_32),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_24),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_136),
.A2(n_34),
.B1(n_44),
.B2(n_43),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_17),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_162),
.B(n_163),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_139),
.B(n_17),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_130),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_18),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_39),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_23),
.Y(n_166)
);

NOR3xp33_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_155),
.C(n_38),
.Y(n_181)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_171),
.C(n_172),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_184),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_143),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_176),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_127),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_174),
.B(n_175),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_124),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_180),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_161),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_182),
.C(n_160),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_37),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_41),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_185),
.A2(n_164),
.B1(n_157),
.B2(n_149),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_149),
.B1(n_157),
.B2(n_146),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_196),
.Y(n_199)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_191),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_197),
.B(n_198),
.Y(n_206)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_179),
.C(n_167),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_203),
.C(n_182),
.Y(n_204)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_201),
.A2(n_180),
.B(n_192),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_189),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_207),
.C(n_208),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_178),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_186),
.C(n_195),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_186),
.C(n_196),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_210),
.A2(n_194),
.B1(n_170),
.B2(n_183),
.Y(n_213)
);

O2A1O1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_202),
.B(n_169),
.C(n_190),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_202),
.B(n_187),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

OAI21x1_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_209),
.B(n_177),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_51),
.Y(n_217)
);


endmodule