module fake_jpeg_13474_n_200 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_200);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_11),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_18),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_3),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_49),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_30),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_17),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_77),
.B(n_1),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_79),
.Y(n_97)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_24),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_67),
.C(n_69),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g93 ( 
.A(n_89),
.B(n_67),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_103),
.B(n_1),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_66),
.B1(n_67),
.B2(n_65),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_80),
.B1(n_75),
.B2(n_60),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_84),
.B1(n_85),
.B2(n_65),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_109),
.A2(n_111),
.B1(n_125),
.B2(n_28),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_104),
.A2(n_86),
.B1(n_80),
.B2(n_62),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_73),
.B(n_58),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_100),
.A2(n_91),
.B1(n_62),
.B2(n_75),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_127),
.Y(n_130)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_120),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_95),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_68),
.B1(n_60),
.B2(n_61),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_128),
.B1(n_2),
.B2(n_4),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_68),
.B1(n_63),
.B2(n_64),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_95),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_126),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_82),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_122),
.B(n_76),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_134),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_125),
.B(n_78),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_81),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_140),
.B1(n_150),
.B2(n_6),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_119),
.B(n_111),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_151),
.C(n_148),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_54),
.C(n_26),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_31),
.C(n_52),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_5),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_130),
.B1(n_144),
.B2(n_143),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_161),
.B1(n_163),
.B2(n_169),
.Y(n_173)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_155),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_160),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_147),
.C(n_142),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_136),
.B(n_33),
.Y(n_164)
);

NOR4xp25_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_14),
.C(n_156),
.D(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_167),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_168),
.Y(n_177)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_162),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_179),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_159),
.A2(n_36),
.B(n_51),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_175),
.C(n_176),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_SL g175 ( 
.A(n_153),
.B(n_29),
.C(n_50),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_10),
.B(n_12),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_152),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_158),
.C(n_19),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_15),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_22),
.Y(n_186)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_178),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_183),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_16),
.C(n_21),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_186),
.C(n_188),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_154),
.B1(n_39),
.B2(n_40),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_190),
.C(n_189),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_187),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_176),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_195),
.A2(n_173),
.B1(n_187),
.B2(n_175),
.Y(n_196)
);

AO21x1_ASAP7_75t_SL g197 ( 
.A1(n_196),
.A2(n_173),
.B(n_191),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_197),
.A2(n_23),
.B(n_41),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_198),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);


endmodule