module fake_jpeg_7155_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_12),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_61),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_26),
.B(n_16),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_59),
.Y(n_78)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_33),
.B(n_15),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_41),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_21),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_15),
.B1(n_31),
.B2(n_23),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_70),
.B1(n_71),
.B2(n_75),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_15),
.B1(n_31),
.B2(n_23),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_31),
.B1(n_23),
.B2(n_20),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_20),
.B1(n_19),
.B2(n_17),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_20),
.B1(n_19),
.B2(n_17),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_22),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_63),
.C(n_26),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_25),
.B1(n_28),
.B2(n_24),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_60),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_97),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_105),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_90),
.Y(n_131)
);

OAI21x1_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_49),
.B(n_48),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_83),
.B1(n_84),
.B2(n_67),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_43),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_93),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_44),
.C(n_18),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_99),
.C(n_95),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_55),
.B(n_62),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_102),
.C(n_18),
.Y(n_121)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_86),
.B(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_53),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_100),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_44),
.C(n_54),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_18),
.B(n_29),
.Y(n_102)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_45),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_18),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_70),
.B(n_10),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_79),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_118),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_88),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_77),
.B1(n_73),
.B2(n_67),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_113),
.A2(n_116),
.B1(n_118),
.B2(n_131),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_104),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_114),
.B(n_107),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_73),
.B1(n_83),
.B2(n_79),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_80),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_108),
.B1(n_103),
.B2(n_97),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_123),
.B1(n_126),
.B2(n_89),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_94),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_80),
.B1(n_42),
.B2(n_47),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_42),
.B1(n_47),
.B2(n_85),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_127),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_0),
.Y(n_157)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_30),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_29),
.B(n_30),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_100),
.Y(n_135)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_93),
.Y(n_138)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_141),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_157),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_119),
.B(n_101),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_152),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_102),
.B(n_96),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_146),
.B1(n_147),
.B2(n_156),
.Y(n_166)
);

NAND2x1p5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_99),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_148),
.B(n_150),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_106),
.B1(n_99),
.B2(n_109),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_90),
.B(n_1),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_133),
.B1(n_120),
.B2(n_137),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_106),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_122),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_154),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_85),
.B1(n_30),
.B2(n_69),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_159),
.C(n_112),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_113),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_162),
.B1(n_176),
.B2(n_3),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_123),
.B1(n_133),
.B2(n_126),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_169),
.C(n_177),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_115),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_164),
.B(n_9),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_167),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_144),
.A2(n_153),
.B1(n_158),
.B2(n_150),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_170),
.B(n_147),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_116),
.C(n_125),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_111),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_111),
.B1(n_119),
.B2(n_134),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_122),
.C(n_127),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_135),
.B(n_8),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_179),
.B(n_148),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_0),
.C(n_1),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_169),
.C(n_163),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_188),
.B(n_198),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_175),
.B(n_156),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_196),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_157),
.B(n_154),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_192),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_174),
.A2(n_145),
.B(n_149),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_145),
.Y(n_193)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

OAI22x1_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_149),
.B1(n_2),
.B2(n_3),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_200),
.B1(n_166),
.B2(n_173),
.Y(n_211)
);

NAND2x1_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_0),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_178),
.B(n_2),
.Y(n_197)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_183),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_201),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_181),
.C(n_177),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_3),
.Y(n_203)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_211),
.A2(n_195),
.B1(n_184),
.B2(n_196),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_187),
.B(n_184),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_162),
.B1(n_168),
.B2(n_170),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_217),
.A2(n_192),
.B1(n_187),
.B2(n_204),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_160),
.C(n_167),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_221),
.C(n_201),
.Y(n_227)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_222),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_160),
.C(n_6),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_223),
.A2(n_232),
.B1(n_205),
.B2(n_212),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_185),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_224),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_228),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_212),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_231),
.Y(n_249)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_214),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_230),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_191),
.C(n_190),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_235),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_199),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_234),
.B(n_236),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_202),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_185),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_208),
.A2(n_194),
.B1(n_196),
.B2(n_189),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_228),
.B(n_217),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_235),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_225),
.A2(n_207),
.B1(n_210),
.B2(n_213),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_243),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_237),
.B(n_216),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_242),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g243 ( 
.A(n_226),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_246),
.A2(n_5),
.B(n_7),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_223),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_251),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_248),
.A2(n_233),
.B(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_255),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_9),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_188),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_248),
.A2(n_209),
.B1(n_221),
.B2(n_8),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_256),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_247),
.B1(n_249),
.B2(n_238),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_258),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_5),
.Y(n_258)
);

FAx1_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_10),
.CI(n_11),
.CON(n_266),
.SN(n_266)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_260),
.A2(n_266),
.B1(n_257),
.B2(n_259),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_7),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_264),
.Y(n_267)
);

AOI21xp33_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_254),
.B(n_250),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_268),
.A2(n_269),
.B(n_270),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_263),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_264),
.Y(n_270)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

A2O1A1O1Ixp25_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_256),
.B(n_266),
.C(n_13),
.D(n_14),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_274),
.A2(n_270),
.B(n_11),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_272),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_275),
.Y(n_277)
);

AO21x1_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_273),
.B(n_276),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_11),
.Y(n_279)
);


endmodule