module fake_jpeg_3301_n_114 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

NAND2xp33_ASAP7_75t_SL g43 ( 
.A(n_42),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_49),
.Y(n_56)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_49),
.B(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_50),
.B(n_2),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_54),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_40),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_33),
.B1(n_47),
.B2(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_44),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_57),
.A2(n_51),
.B1(n_55),
.B2(n_52),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_68),
.B1(n_61),
.B2(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_34),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_41),
.B1(n_36),
.B2(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_80),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_82),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_41),
.C(n_17),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

OAI22x1_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_3),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_89),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_5),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_91),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_73),
.B(n_81),
.C(n_80),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_5),
.B(n_6),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_6),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_23),
.Y(n_101)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_89),
.B1(n_85),
.B2(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_98),
.B(n_100),
.Y(n_104)
);

NOR2xp67_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_22),
.Y(n_99)
);

OAI321xp33_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_101),
.A3(n_24),
.B1(n_31),
.B2(n_30),
.C(n_11),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_103),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_85),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_104),
.A2(n_95),
.B(n_101),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_103),
.B1(n_106),
.B2(n_105),
.Y(n_109)
);

OAI31xp33_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_107),
.A3(n_8),
.B(n_9),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_7),
.B(n_13),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_14),
.C(n_15),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_27),
.Y(n_114)
);


endmodule