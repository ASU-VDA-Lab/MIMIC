module fake_jpeg_17409_n_184 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_SL g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_33),
.B(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_2),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_47),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_4),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_17),
.Y(n_68)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_18),
.A2(n_4),
.B(n_5),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_4),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_54),
.Y(n_85)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_62),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_24),
.B1(n_22),
.B2(n_20),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_20),
.B1(n_17),
.B2(n_32),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_7),
.B(n_9),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_46),
.B(n_27),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_73),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_18),
.B1(n_15),
.B2(n_22),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_15),
.B1(n_31),
.B2(n_29),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_27),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_72),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_7),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_32),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_86),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_71),
.B1(n_49),
.B2(n_50),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_78),
.B(n_92),
.Y(n_114)
);

OR2x2_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_26),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_SL g117 ( 
.A(n_79),
.B(n_83),
.C(n_95),
.Y(n_117)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_44),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_29),
.C(n_31),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_59),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_91),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_31),
.B1(n_29),
.B2(n_28),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_59),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_94),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_38),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_97),
.Y(n_113)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_89),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_115),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_63),
.B1(n_70),
.B2(n_66),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_97),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_105),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_85),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_72),
.B1(n_66),
.B2(n_51),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_89),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_87),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_56),
.B1(n_30),
.B2(n_28),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_60),
.B1(n_61),
.B2(n_12),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_118),
.B1(n_113),
.B2(n_100),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_127),
.B(n_128),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_88),
.C(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_93),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_115),
.Y(n_140)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_93),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_137),
.B(n_117),
.Y(n_156)
);

AO221x1_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_112),
.B1(n_107),
.B2(n_99),
.C(n_80),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_148),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_96),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_126),
.A2(n_100),
.B(n_118),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_77),
.B(n_82),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_107),
.B(n_102),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_97),
.B(n_131),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_129),
.B1(n_135),
.B2(n_120),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_144),
.B1(n_129),
.B2(n_120),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_102),
.B1(n_119),
.B2(n_117),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_149),
.A2(n_134),
.B1(n_126),
.B2(n_102),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_127),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_158),
.Y(n_161)
);

AOI21x1_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_95),
.B(n_112),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_148),
.B1(n_145),
.B2(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_77),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_160),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_159),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_151),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_152),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_141),
.C(n_140),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_11),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_168),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_160),
.B(n_82),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_169),
.B(n_164),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_166),
.B(n_165),
.C(n_163),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_10),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_171),
.B(n_11),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_162),
.C(n_164),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_174),
.B(n_175),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_176),
.B(n_177),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_178),
.Y(n_181)
);

NAND3xp33_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_173),
.C(n_172),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_179),
.B1(n_12),
.B2(n_13),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_181),
.Y(n_184)
);


endmodule