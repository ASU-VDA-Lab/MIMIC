module real_jpeg_28699_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_242;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_244;
wire n_213;
wire n_128;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_0),
.A2(n_40),
.B1(n_49),
.B2(n_50),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_0),
.A2(n_26),
.B1(n_28),
.B2(n_40),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_0),
.A2(n_40),
.B1(n_58),
.B2(n_59),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_1),
.B(n_58),
.Y(n_57)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_1),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_2),
.A2(n_49),
.B1(n_50),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_2),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_2),
.A2(n_58),
.B1(n_59),
.B2(n_77),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_77),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_3),
.A2(n_26),
.B1(n_28),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_3),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g162 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_99),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_3),
.A2(n_49),
.B1(n_50),
.B2(n_99),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_3),
.A2(n_58),
.B1(n_59),
.B2(n_99),
.Y(n_219)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_5),
.A2(n_26),
.B1(n_28),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_5),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_136),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_5),
.A2(n_49),
.B1(n_50),
.B2(n_136),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_136),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_6),
.A2(n_58),
.B1(n_59),
.B2(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_63),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_8),
.A2(n_26),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_8),
.A2(n_37),
.B1(n_49),
.B2(n_50),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_8),
.A2(n_37),
.B1(n_58),
.B2(n_59),
.Y(n_214)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_10),
.A2(n_25),
.B1(n_33),
.B2(n_34),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_10),
.A2(n_25),
.B1(n_58),
.B2(n_59),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_10),
.A2(n_25),
.B1(n_49),
.B2(n_50),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_11),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_73),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_15),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_SL g141 ( 
.A1(n_15),
.A2(n_30),
.B(n_34),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_15),
.A2(n_26),
.B1(n_28),
.B2(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_15),
.B(n_32),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_15),
.A2(n_49),
.B(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_15),
.B(n_49),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_15),
.B(n_53),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_15),
.A2(n_56),
.B1(n_66),
.B2(n_225),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_15),
.A2(n_33),
.B(n_241),
.Y(n_240)
);

INVx11_ASAP7_75t_SL g61 ( 
.A(n_16),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_17),
.A2(n_58),
.B1(n_59),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_17),
.A2(n_49),
.B1(n_50),
.B2(n_68),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_127),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_125),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_102),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_21),
.B(n_102),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_78),
.C(n_89),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_22),
.B(n_78),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_22),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_38),
.CI(n_54),
.CON(n_22),
.SN(n_22)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_23),
.B(n_38),
.C(n_54),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_24),
.A2(n_29),
.B1(n_32),
.B2(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_26),
.A2(n_35),
.B(n_140),
.C(n_141),
.Y(n_139)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_30),
.Y(n_31)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_29),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_29),
.A2(n_32),
.B1(n_135),
.B2(n_164),
.Y(n_163)
);

AO22x1_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_32),
.Y(n_119)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_43),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g249 ( 
.A1(n_33),
.A2(n_47),
.A3(n_50),
.B1(n_242),
.B2(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_34),
.B(n_140),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_36),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_51),
.B2(n_53),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_39),
.A2(n_41),
.B1(n_53),
.B2(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_41),
.A2(n_53),
.B1(n_162),
.B2(n_181),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_42),
.A2(n_46),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_42),
.A2(n_46),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_42),
.A2(n_46),
.B1(n_145),
.B2(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_42),
.A2(n_46),
.B1(n_182),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_47),
.Y(n_251)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_50),
.B1(n_73),
.B2(n_75),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_49),
.A2(n_59),
.A3(n_75),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_49),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_69),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_55),
.B(n_69),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_67),
.B(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_56),
.A2(n_62),
.B1(n_64),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_56),
.A2(n_88),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_56),
.A2(n_66),
.B1(n_219),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_56),
.A2(n_88),
.B1(n_214),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_57),
.A2(n_65),
.B1(n_93),
.B2(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_57),
.A2(n_65),
.B1(n_143),
.B2(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_57),
.A2(n_65),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_58),
.B(n_73),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_58),
.B(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_SL g88 ( 
.A(n_65),
.Y(n_88)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_76),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_72),
.B1(n_84),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_71),
.A2(n_72),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_71),
.A2(n_72),
.B1(n_200),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_71),
.A2(n_72),
.B1(n_167),
.B2(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_72),
.B(n_140),
.Y(n_226)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_76),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_86),
.B2(n_87),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_79),
.B(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_82),
.A2(n_85),
.B1(n_96),
.B2(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_82),
.A2(n_85),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_87),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_89),
.B(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_97),
.C(n_100),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_90),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_91),
.B(n_94),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_100),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_98),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_101),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_123),
.B2(n_124),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_112),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B(n_111),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_109),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_117),
.A2(n_119),
.B1(n_134),
.B2(n_137),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_123),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_150),
.B(n_277),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_148),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_129),
.B(n_148),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_147),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_147),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.C(n_144),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_144),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_138),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_142),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_140),
.B(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_187),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_170),
.B(n_186),
.Y(n_152)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_168),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_154),
.B(n_168),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.C(n_158),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_158),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.C(n_165),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_159),
.A2(n_160),
.B1(n_165),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_173),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.C(n_178),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_174),
.B(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_275),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_177),
.Y(n_275)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.C(n_185),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_180),
.B(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_183),
.B(n_185),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_184),
.Y(n_253)
);

NOR3xp33_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_189),
.C(n_190),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_271),
.B(n_276),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_257),
.B(n_270),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_235),
.B(n_256),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_215),
.B(n_234),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_205),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_195),
.B(n_205),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_197),
.B1(n_201),
.B2(n_202),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_199),
.Y(n_203)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_210),
.C(n_212),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_211),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_213),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_222),
.B(n_233),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_217),
.B(n_221),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_227),
.B(n_232),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_226),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_236),
.B(n_237),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_248),
.B1(n_254),
.B2(n_255),
.Y(n_237)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_243),
.B1(n_246),
.B2(n_247),
.Y(n_238)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_247),
.C(n_255),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_245),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_248),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_252),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_258),
.B(n_259),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_266),
.C(n_268),
.Y(n_272)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);


endmodule