module fake_jpeg_3977_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_2),
.B(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_8),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_57),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_19),
.B1(n_23),
.B2(n_26),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_48),
.A2(n_54),
.B1(n_55),
.B2(n_68),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_19),
.B1(n_23),
.B2(n_26),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_19),
.B1(n_23),
.B2(n_26),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_56),
.Y(n_85)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_19),
.B1(n_26),
.B2(n_31),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_38),
.B1(n_64),
.B2(n_33),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_29),
.B1(n_17),
.B2(n_28),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_29),
.B1(n_33),
.B2(n_24),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_36),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_30),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_72),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_30),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_41),
.B(n_37),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_73),
.A2(n_93),
.B(n_97),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_21),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_40),
.B(n_32),
.C(n_31),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_77),
.B(n_90),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_44),
.B1(n_38),
.B2(n_45),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_79),
.A2(n_61),
.B1(n_66),
.B2(n_21),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_44),
.B1(n_38),
.B2(n_22),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_83),
.B1(n_92),
.B2(n_31),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_64),
.B1(n_49),
.B2(n_63),
.Y(n_83)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_53),
.B(n_31),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_51),
.B(n_18),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_96),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_58),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_64),
.A2(n_40),
.B1(n_30),
.B2(n_35),
.Y(n_92)
);

NAND2x1_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_46),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_49),
.A2(n_28),
.B1(n_25),
.B2(n_22),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_25),
.B1(n_18),
.B2(n_35),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_51),
.B(n_24),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_58),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

OAI32xp33_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_18),
.A3(n_35),
.B1(n_33),
.B2(n_24),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_100),
.B(n_102),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_101),
.A2(n_119),
.B1(n_76),
.B2(n_80),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_78),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_104),
.B(n_111),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_71),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_106),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_107),
.A2(n_124),
.B1(n_90),
.B2(n_94),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_79),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_84),
.B(n_98),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_0),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_121),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_65),
.B1(n_60),
.B2(n_57),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_52),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_78),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_116),
.B(n_122),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_99),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_89),
.A2(n_47),
.B1(n_61),
.B2(n_46),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_58),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_52),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_77),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_79),
.Y(n_127)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_73),
.C(n_79),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_149),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_86),
.C(n_79),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_130),
.A2(n_27),
.B(n_20),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_126),
.A2(n_81),
.B1(n_83),
.B2(n_82),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_133),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_127),
.B1(n_107),
.B2(n_125),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_115),
.B(n_104),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_91),
.B1(n_84),
.B2(n_80),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_140),
.Y(n_168)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_142),
.Y(n_182)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_143),
.A2(n_124),
.B1(n_101),
.B2(n_108),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_145),
.B(n_148),
.Y(n_183)
);

INVx2_ASAP7_75t_R g147 ( 
.A(n_127),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_122),
.C(n_109),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_87),
.C(n_94),
.Y(n_149)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_153),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_87),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_154),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_100),
.A2(n_91),
.B1(n_58),
.B2(n_66),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_105),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_161),
.B(n_162),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_152),
.B(n_117),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_131),
.B(n_154),
.Y(n_197)
);

AND2x6_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_100),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_132),
.Y(n_198)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_174),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_155),
.B(n_135),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_170),
.A2(n_191),
.B(n_21),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_102),
.B1(n_113),
.B2(n_105),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_171),
.A2(n_175),
.B1(n_176),
.B2(n_180),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_145),
.B(n_120),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_178),
.C(n_128),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_120),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_177),
.A2(n_181),
.B1(n_190),
.B2(n_146),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_143),
.B(n_119),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_147),
.A2(n_103),
.B1(n_46),
.B2(n_52),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_158),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_185),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_50),
.Y(n_187)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_189),
.A2(n_27),
.B(n_20),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_147),
.A2(n_50),
.B1(n_21),
.B2(n_75),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_198),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_149),
.C(n_142),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_203),
.C(n_204),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_197),
.B(n_159),
.Y(n_234)
);

OAI21x1_ASAP7_75t_SL g199 ( 
.A1(n_167),
.A2(n_130),
.B(n_137),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_199),
.A2(n_200),
.B1(n_176),
.B2(n_169),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_137),
.B1(n_129),
.B2(n_50),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_201),
.A2(n_213),
.B1(n_215),
.B2(n_191),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_75),
.C(n_27),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_27),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_190),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_27),
.C(n_20),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_209),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_165),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_208),
.B(n_214),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_170),
.A2(n_27),
.B(n_20),
.Y(n_209)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_163),
.A2(n_27),
.B1(n_20),
.B2(n_0),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_217),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_177),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_160),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_166),
.A2(n_1),
.B(n_3),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_15),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_220),
.C(n_175),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_183),
.A2(n_159),
.B(n_168),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_196),
.B(n_192),
.Y(n_221)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_221),
.B(n_15),
.C(n_7),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_194),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_223),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_206),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_210),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_161),
.Y(n_236)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_240),
.B1(n_243),
.B2(n_244),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_202),
.B(n_184),
.Y(n_241)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_195),
.B(n_164),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_219),
.A2(n_186),
.B1(n_182),
.B2(n_178),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_197),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_193),
.C(n_205),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_187),
.Y(n_246)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_216),
.B(n_215),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_247),
.B(n_256),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_233),
.B(n_200),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_262),
.C(n_237),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_203),
.C(n_204),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_258),
.C(n_254),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_256),
.B(n_235),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_207),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_255),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_211),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_232),
.A2(n_209),
.B1(n_181),
.B2(n_180),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_4),
.C(n_5),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_239),
.B1(n_228),
.B2(n_229),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_237),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_269),
.C(n_280),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_248),
.C(n_255),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_249),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_272),
.Y(n_287)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_225),
.B1(n_238),
.B2(n_226),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_274),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_297)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

BUFx24_ASAP7_75t_SL g295 ( 
.A(n_276),
.Y(n_295)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_6),
.Y(n_292)
);

AOI21xp33_ASAP7_75t_L g278 ( 
.A1(n_267),
.A2(n_236),
.B(n_246),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_278),
.A2(n_251),
.B(n_266),
.Y(n_291)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

AND2x2_ASAP7_75t_SL g281 ( 
.A(n_261),
.B(n_225),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_282),
.B(n_264),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_231),
.C(n_7),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_265),
.C(n_247),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_291),
.B(n_292),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_298),
.C(n_279),
.Y(n_304)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_297),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_268),
.C(n_270),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_301),
.Y(n_317)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_282),
.B(n_281),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_SL g315 ( 
.A1(n_302),
.A2(n_285),
.B(n_289),
.C(n_286),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_281),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_305),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_298),
.C(n_286),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_270),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_307),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_10),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_11),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_309),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_295),
.B(n_280),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_296),
.B(n_11),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_12),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_291),
.Y(n_312)
);

AOI321xp33_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_315),
.C(n_311),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_301),
.Y(n_320)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_315),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_12),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_321),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_302),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_323),
.A2(n_324),
.B(n_14),
.Y(n_327)
);

OAI21x1_ASAP7_75t_SL g324 ( 
.A1(n_317),
.A2(n_14),
.B(n_314),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_323),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_326),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_325),
.B1(n_328),
.B2(n_316),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_327),
.B(n_322),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);


endmodule