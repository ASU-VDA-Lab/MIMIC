module fake_jpeg_30508_n_118 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_17),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_3),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_3),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_57),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_4),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_5),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_6),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_59),
.Y(n_72)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_SL g61 ( 
.A(n_55),
.B(n_46),
.C(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_69),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_41),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_68),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_41),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_76),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_38),
.B1(n_47),
.B2(n_40),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_24),
.B(n_27),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_38),
.B1(n_22),
.B2(n_9),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_7),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_7),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_8),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_8),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_12),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_94),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_16),
.B(n_18),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_102),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_83),
.C(n_34),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_106),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_32),
.C(n_35),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_91),
.B(n_96),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_103),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_109),
.B(n_92),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_107),
.C(n_111),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_112),
.Y(n_116)
);

FAx1_ASAP7_75t_SL g117 ( 
.A(n_116),
.B(n_102),
.CI(n_90),
.CON(n_117),
.SN(n_117)
);

AOI221xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_95),
.B1(n_110),
.B2(n_97),
.C(n_94),
.Y(n_118)
);


endmodule