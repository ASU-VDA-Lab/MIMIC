module fake_jpeg_23166_n_133 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_133);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx2_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_31),
.Y(n_44)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_17),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_37),
.B1(n_17),
.B2(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_17),
.A2(n_3),
.B1(n_13),
.B2(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_41),
.Y(n_52)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_4),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_18),
.Y(n_54)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx2_ASAP7_75t_SL g81 ( 
.A(n_47),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_16),
.C(n_19),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_62),
.C(n_23),
.Y(n_73)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_60),
.B1(n_23),
.B2(n_22),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_32),
.A2(n_18),
.B1(n_38),
.B2(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_28),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_20),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_33),
.B(n_26),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_27),
.B1(n_21),
.B2(n_25),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_69),
.B1(n_75),
.B2(n_78),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_27),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_61),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_62),
.A2(n_30),
.B1(n_26),
.B2(n_25),
.Y(n_68)
);

OAI22x1_ASAP7_75t_SL g94 ( 
.A1(n_68),
.A2(n_53),
.B1(n_22),
.B2(n_57),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_55),
.B1(n_14),
.B2(n_48),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_82),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_23),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_47),
.B(n_58),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_79),
.B(n_43),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_40),
.B1(n_33),
.B2(n_29),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_33),
.B1(n_22),
.B2(n_23),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_83),
.B(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_65),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_95),
.B1(n_77),
.B2(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_51),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_75),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_68),
.B1(n_78),
.B2(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_4),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_99),
.B1(n_90),
.B2(n_82),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_94),
.B1(n_85),
.B2(n_86),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_73),
.C(n_43),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_84),
.C(n_83),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_103),
.B(n_65),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_71),
.B(n_70),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_100),
.B(n_97),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_102),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_109),
.B(n_110),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_105),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_101),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_114),
.B(n_104),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_115),
.B1(n_99),
.B2(n_82),
.Y(n_119)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_117),
.B(n_118),
.CI(n_119),
.CON(n_123),
.SN(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_114),
.A2(n_106),
.B(n_107),
.C(n_101),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_9),
.Y(n_125)
);

AO22x1_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_112),
.B1(n_108),
.B2(n_59),
.Y(n_122)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_6),
.C(n_7),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_126),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_12),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_9),
.C(n_10),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_128),
.A2(n_125),
.B1(n_90),
.B2(n_123),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_131),
.Y(n_132)
);

OAI21x1_ASAP7_75t_SL g131 ( 
.A1(n_129),
.A2(n_123),
.B(n_67),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_127),
.Y(n_133)
);


endmodule