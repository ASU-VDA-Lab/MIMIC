module real_jpeg_4109_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_0),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_0),
.B(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_0),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_0),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_0),
.B(n_284),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_0),
.B(n_326),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_0),
.B(n_305),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_0),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_1),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_1),
.B(n_95),
.Y(n_162)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_1),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_1),
.B(n_291),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_1),
.B(n_326),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_1),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_1),
.B(n_407),
.Y(n_406)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_2),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_2),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_2),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_3),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_3),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_3),
.Y(n_233)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_3),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_4),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_5),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_5),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_5),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_5),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_5),
.B(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_5),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_5),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_5),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_6),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_6),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_6),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_6),
.B(n_335),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_6),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_6),
.B(n_382),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_6),
.B(n_397),
.Y(n_396)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_7),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_7),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_9),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_9),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_9),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_9),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_9),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_9),
.B(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_10),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_10),
.Y(n_204)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_10),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_10),
.Y(n_311)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_12),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_12),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_12),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_13),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_13),
.B(n_44),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_13),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_13),
.B(n_309),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_13),
.B(n_324),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_13),
.B(n_281),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_13),
.B(n_377),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_13),
.B(n_100),
.Y(n_403)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_15),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_15),
.B(n_50),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_15),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_15),
.B(n_34),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_15),
.B(n_218),
.Y(n_217)
);

AND2x2_ASAP7_75t_SL g280 ( 
.A(n_15),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_15),
.B(n_326),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_15),
.B(n_173),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_16),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_16),
.B(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_16),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_16),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_16),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_16),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_16),
.B(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_16),
.B(n_176),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_17),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_17),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_17),
.B(n_305),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_17),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_17),
.B(n_348),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_17),
.B(n_384),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_17),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_18),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_18),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_18),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_18),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_18),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_18),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_18),
.B(n_256),
.Y(n_255)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B(n_525),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx13_ASAP7_75t_L g526 ( 
.A(n_22),
.Y(n_526)
);

O2A1O1Ixp33_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_40),
.B(n_78),
.C(n_524),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_45),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_26),
.B(n_45),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_38),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.C(n_36),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_28),
.A2(n_31),
.B1(n_39),
.B2(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_29),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_49),
.C(n_57),
.Y(n_75)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_35),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_35),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_36),
.B(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_74),
.C(n_76),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_46),
.B(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_61),
.C(n_64),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_47),
.B(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_57),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_49),
.A2(n_56),
.B1(n_70),
.B2(n_113),
.Y(n_117)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_51),
.B(n_270),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_53),
.Y(n_147)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_54),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_54),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_65),
.C(n_70),
.Y(n_64)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_61),
.B(n_64),
.Y(n_120)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_65),
.A2(n_66),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_70),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_70),
.A2(n_108),
.B1(n_109),
.B2(n_113),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_72),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_72),
.Y(n_216)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_72),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_72),
.Y(n_407)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_73),
.Y(n_336)
);

BUFx5_ASAP7_75t_L g349 ( 
.A(n_73),
.Y(n_349)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_73),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_76),
.Y(n_123)
);

AO21x1_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_124),
.B(n_523),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_121),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_80),
.B(n_121),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_118),
.C(n_119),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_81),
.A2(n_82),
.B1(n_519),
.B2(n_520),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_106),
.C(n_114),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_83),
.A2(n_84),
.B1(n_499),
.B2(n_501),
.Y(n_498)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_93),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_89),
.C(n_93),
.Y(n_118)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_88),
.Y(n_265)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_88),
.Y(n_397)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.C(n_101),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_94),
.B(n_489),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_96),
.A2(n_97),
.B1(n_101),
.B2(n_102),
.Y(n_489)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_106),
.A2(n_114),
.B1(n_115),
.B2(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_106),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.C(n_113),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_107),
.B(n_495),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_108),
.A2(n_109),
.B1(n_190),
.B2(n_194),
.Y(n_189)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_109),
.B(n_187),
.C(n_190),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_118),
.B(n_119),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_517),
.B(n_522),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_482),
.B(n_514),
.Y(n_125)
);

OAI21x1_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_293),
.B(n_481),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_241),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_128),
.B(n_241),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_184),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_129),
.B(n_185),
.C(n_219),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_160),
.C(n_167),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_130),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_138),
.C(n_148),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_131),
.B(n_466),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_135),
.C(n_136),
.Y(n_166)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_138),
.A2(n_139),
.B1(n_148),
.B2(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_146),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_140),
.B(n_146),
.Y(n_456)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_143),
.B(n_456),
.Y(n_455)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_148),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_149),
.B(n_151),
.C(n_156),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_155),
.B1(n_156),
.B2(n_159),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_155),
.B(n_190),
.C(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_155),
.A2(n_156),
.B1(n_190),
.B2(n_194),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_158),
.Y(n_256)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_158),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_160),
.B(n_167),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_166),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_162),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_163),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_163),
.B(n_164),
.C(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_163),
.A2(n_165),
.B1(n_230),
.B2(n_234),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_165),
.B(n_224),
.C(n_234),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_178),
.C(n_181),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_168),
.B(n_273),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.C(n_175),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_169),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_172),
.B(n_175),
.Y(n_253)
);

BUFx8_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_174),
.Y(n_268)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_178),
.B(n_181),
.Y(n_273)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_183),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_183),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_219),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_195),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_186),
.B(n_196),
.C(n_208),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_190),
.Y(n_194)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_208),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.C(n_205),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_205),
.Y(n_240)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_200),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_200),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_204),
.Y(n_281)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_217),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_210),
.B(n_213),
.C(n_217),
.Y(n_497)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_235),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_221),
.B(n_223),
.C(n_235),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_225),
.B(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.C(n_239),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_239),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_248),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_243),
.B(n_246),
.Y(n_476)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_248),
.B(n_476),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_271),
.C(n_274),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_250),
.B(n_469),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.C(n_261),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_251),
.A2(n_252),
.B1(n_447),
.B2(n_448),
.Y(n_446)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_254),
.A2(n_255),
.B(n_257),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_254),
.B(n_261),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.C(n_269),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_262),
.A2(n_263),
.B1(n_266),
.B2(n_267),
.Y(n_424)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_269),
.B(n_424),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_270),
.B(n_365),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_274),
.Y(n_470)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_286),
.C(n_290),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_276),
.B(n_458),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.C(n_282),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_277),
.B(n_436),
.Y(n_435)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_280),
.A2(n_282),
.B1(n_283),
.B2(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_280),
.Y(n_437)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_286),
.B(n_290),
.Y(n_458)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx8_ASAP7_75t_L g405 ( 
.A(n_288),
.Y(n_405)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_289),
.Y(n_332)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_291),
.Y(n_395)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_474),
.B(n_480),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_461),
.B(n_473),
.Y(n_294)
);

AOI21x1_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_443),
.B(n_460),
.Y(n_295)
);

OAI21x1_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_417),
.B(n_442),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_388),
.B(n_416),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_357),
.B(n_387),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_338),
.B(n_356),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_318),
.B(n_337),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_312),
.B(n_317),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_310),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_310),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_308),
.Y(n_319)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_307),
.Y(n_343)
);

INVx4_ASAP7_75t_SL g365 ( 
.A(n_311),
.Y(n_365)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_320),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_327),
.B2(n_328),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_321),
.B(n_330),
.C(n_333),
.Y(n_355)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_325),
.Y(n_345)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_329),
.A2(n_330),
.B1(n_333),
.B2(n_334),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_355),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_355),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_346),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_345),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_345),
.C(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_344),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_342),
.B(n_344),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_346),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_350),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_347),
.B(n_373),
.C(n_374),
.Y(n_372)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_351),
.Y(n_373)
);

INVx6_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_354),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_360),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_371),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_361),
.B(n_372),
.C(n_375),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_362),
.B(n_364),
.C(n_366),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_368),
.B1(n_369),
.B2(n_370),
.Y(n_366)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_367),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_368),
.B(n_370),
.Y(n_398)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_375),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_380),
.Y(n_375)
);

MAJx2_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_383),
.C(n_385),
.Y(n_414)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_381),
.A2(n_383),
.B1(n_385),
.B2(n_386),
.Y(n_380)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_381),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_383),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_415),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_415),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_400),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_399),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_391),
.B(n_399),
.C(n_441),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_398),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_396),
.Y(n_392)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_393),
.Y(n_431)
);

INVx5_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_396),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_398),
.B(n_431),
.C(n_432),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_400),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_408),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_401),
.B(n_410),
.C(n_413),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_406),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

MAJx2_ASAP7_75t_L g428 ( 
.A(n_403),
.B(n_404),
.C(n_406),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_410),
.B1(n_413),
.B2(n_414),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_412),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_414),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_440),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_440),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_429),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_420),
.B(n_421),
.C(n_429),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_422),
.A2(n_423),
.B1(n_425),
.B2(n_426),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_422),
.B(n_452),
.C(n_453),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_427),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_428),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_433),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_434),
.C(n_439),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_435),
.B1(n_438),
.B2(n_439),
.Y(n_433)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_434),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_435),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_459),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_459),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_445),
.B(n_450),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_449),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_449),
.C(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_447),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_450),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_454),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_455),
.C(n_457),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_457),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_462),
.B(n_471),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_462),
.B(n_471),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_463),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_468),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_465),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_468),
.B(n_478),
.C(n_479),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_477),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_477),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_510),
.Y(n_482)
);

OAI21xp33_ASAP7_75t_L g514 ( 
.A1(n_483),
.A2(n_515),
.B(n_516),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_484),
.B(n_503),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_484),
.B(n_503),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_486),
.B1(n_492),
.B2(n_502),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_485),
.B(n_493),
.C(n_498),
.Y(n_521)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.C(n_490),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_487),
.B(n_505),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_488),
.A2(n_490),
.B1(n_491),
.B2(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_488),
.Y(n_506)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_492),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_498),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_496),
.C(n_497),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_508),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_496),
.B(n_497),
.Y(n_508)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_499),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_507),
.C(n_509),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_504),
.B(n_507),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_509),
.B(n_512),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_511),
.B(n_513),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_511),
.B(n_513),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_521),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_518),
.B(n_521),
.Y(n_522)
);

CKINVDCx14_ASAP7_75t_R g520 ( 
.A(n_519),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_527),
.Y(n_525)
);


endmodule