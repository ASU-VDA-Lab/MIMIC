module fake_netlist_1_10660_n_38 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_5), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_3), .Y(n_13) );
BUFx6f_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_5), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_8), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_6), .Y(n_17) );
AOI22xp5_ASAP7_75t_L g18 ( .A1(n_13), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
NAND3xp33_ASAP7_75t_SL g20 ( .A(n_12), .B(n_0), .C(n_1), .Y(n_20) );
BUFx6f_ASAP7_75t_L g21 ( .A(n_14), .Y(n_21) );
AOI22xp33_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_22) );
HB1xp67_ASAP7_75t_L g23 ( .A(n_18), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_14), .B1(n_19), .B2(n_21), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
INVx1_ASAP7_75t_SL g28 ( .A(n_26), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
INVx2_ASAP7_75t_SL g30 ( .A(n_28), .Y(n_30) );
AOI22xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_17), .B1(n_21), .B2(n_6), .Y(n_31) );
XNOR2xp5_ASAP7_75t_L g32 ( .A(n_29), .B(n_2), .Y(n_32) );
AOI22xp33_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_21), .B1(n_4), .B2(n_9), .Y(n_33) );
OAI22xp5_ASAP7_75t_L g34 ( .A1(n_30), .A2(n_4), .B1(n_7), .B2(n_10), .Y(n_34) );
HB1xp67_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
INVx2_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_33), .Y(n_37) );
OAI222xp33_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_11), .B1(n_31), .B2(n_35), .C1(n_36), .C2(n_32), .Y(n_38) );
endmodule