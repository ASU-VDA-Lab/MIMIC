module fake_jpeg_31636_n_552 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_552);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_552;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_9),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_6),
.B(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_56),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_11),
.B1(n_17),
.B2(n_16),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_58),
.A2(n_20),
.B1(n_47),
.B2(n_42),
.Y(n_149)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_59),
.Y(n_148)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_61),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_11),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_62),
.B(n_70),
.Y(n_119)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_26),
.B(n_11),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_69),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_25),
.B(n_8),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g71 ( 
.A(n_31),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_71),
.B(n_101),
.Y(n_154)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_78),
.Y(n_133)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_25),
.B(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_85),
.B(n_88),
.Y(n_135)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_86),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_25),
.B(n_8),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_95),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_26),
.B(n_12),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_104),
.B(n_19),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_74),
.A2(n_26),
.B1(n_45),
.B2(n_29),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_107),
.A2(n_153),
.B1(n_38),
.B2(n_40),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_44),
.B1(n_29),
.B2(n_27),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_110),
.A2(n_167),
.B1(n_38),
.B2(n_40),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_70),
.B(n_41),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_112),
.B(n_143),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_85),
.B(n_41),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_120),
.B(n_144),
.C(n_155),
.Y(n_187)
);

NOR2x1_ASAP7_75t_R g130 ( 
.A(n_67),
.B(n_45),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_130),
.B(n_149),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_104),
.B(n_41),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_39),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_59),
.A2(n_45),
.B1(n_44),
.B2(n_39),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_71),
.B(n_39),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_102),
.B(n_32),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_38),
.Y(n_190)
);

NOR2x1_ASAP7_75t_L g163 ( 
.A(n_69),
.B(n_32),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_163),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_52),
.A2(n_44),
.B1(n_51),
.B2(n_24),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_168),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_169),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_94),
.B1(n_93),
.B2(n_91),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_170),
.A2(n_179),
.B1(n_215),
.B2(n_162),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_159),
.A2(n_45),
.B1(n_83),
.B2(n_75),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_171),
.A2(n_181),
.B1(n_184),
.B2(n_122),
.Y(n_235)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_172),
.Y(n_271)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_173),
.Y(n_273)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_174),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_115),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_178),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_84),
.B1(n_80),
.B2(n_78),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_159),
.A2(n_61),
.B1(n_63),
.B2(n_32),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_134),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_182),
.B(n_188),
.Y(n_234)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_134),
.A2(n_20),
.B1(n_51),
.B2(n_47),
.Y(n_184)
);

BUFx4f_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_185),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_135),
.A2(n_119),
.B(n_154),
.C(n_113),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_19),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_189),
.B(n_192),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_190),
.B(n_228),
.Y(n_278)
);

AO22x1_ASAP7_75t_SL g191 ( 
.A1(n_110),
.A2(n_65),
.B1(n_64),
.B2(n_56),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g274 ( 
.A1(n_191),
.A2(n_214),
.B1(n_43),
.B2(n_19),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_132),
.B(n_19),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_37),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_203),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_107),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_195),
.B(n_198),
.Y(n_261)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_199),
.Y(n_260)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_200),
.Y(n_259)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_201),
.Y(n_264)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_147),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_202),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_118),
.B(n_37),
.Y(n_203)
);

AND2x4_ASAP7_75t_L g204 ( 
.A(n_153),
.B(n_43),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_127),
.B(n_37),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_206),
.A2(n_24),
.B1(n_137),
.B2(n_43),
.Y(n_258)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_210),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_211),
.A2(n_216),
.B1(n_219),
.B2(n_227),
.Y(n_244)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_212),
.Y(n_263)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_136),
.Y(n_213)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_150),
.A2(n_33),
.B1(n_51),
.B2(n_47),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_161),
.A2(n_54),
.B1(n_33),
.B2(n_42),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_167),
.A2(n_40),
.B1(n_27),
.B2(n_30),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_146),
.Y(n_217)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_217),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_126),
.B(n_27),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_190),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_123),
.A2(n_42),
.B1(n_33),
.B2(n_30),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_125),
.Y(n_220)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_220),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_160),
.Y(n_221)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_221),
.Y(n_280)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_148),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_224),
.Y(n_276)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_140),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_223),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_109),
.B(n_19),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_115),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_225),
.A2(n_158),
.B1(n_126),
.B2(n_133),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_105),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_226),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_161),
.A2(n_30),
.B1(n_24),
.B2(n_20),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_124),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_137),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_229),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_235),
.B(n_246),
.Y(n_283)
);

OAI22x1_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_137),
.B1(n_105),
.B2(n_122),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g300 ( 
.A1(n_238),
.A2(n_185),
.B(n_226),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_193),
.A2(n_157),
.B1(n_139),
.B2(n_131),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_241),
.A2(n_247),
.B1(n_257),
.B2(n_272),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_245),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_197),
.A2(n_208),
.B1(n_198),
.B2(n_203),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_114),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_248),
.B(n_265),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_SL g250 ( 
.A1(n_205),
.A2(n_158),
.B(n_111),
.Y(n_250)
);

AOI32xp33_ASAP7_75t_L g320 ( 
.A1(n_250),
.A2(n_12),
.A3(n_17),
.B1(n_3),
.B2(n_4),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_204),
.A2(n_111),
.B1(n_162),
.B2(n_125),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_197),
.B(n_128),
.C(n_150),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_270),
.C(n_277),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_258),
.A2(n_244),
.B1(n_265),
.B2(n_248),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_211),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_218),
.B(n_139),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_268),
.B(n_281),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_186),
.B(n_157),
.C(n_131),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_204),
.A2(n_191),
.B1(n_216),
.B2(n_214),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_274),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_187),
.B(n_188),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_186),
.B(n_43),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_238),
.A2(n_191),
.B1(n_178),
.B2(n_183),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_284),
.A2(n_295),
.B1(n_314),
.B2(n_322),
.Y(n_332)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_285),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_236),
.A2(n_228),
.B(n_210),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_286),
.A2(n_324),
.B(n_14),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_264),
.A2(n_221),
.B1(n_282),
.B2(n_201),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_287),
.Y(n_333)
);

AO22x1_ASAP7_75t_SL g288 ( 
.A1(n_236),
.A2(n_173),
.B1(n_172),
.B2(n_196),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_288),
.B(n_311),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_264),
.A2(n_194),
.B1(n_217),
.B2(n_202),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_291),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_292),
.A2(n_293),
.B1(n_296),
.B2(n_298),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_244),
.A2(n_233),
.B1(n_272),
.B2(n_258),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_261),
.A2(n_180),
.B1(n_209),
.B2(n_207),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_233),
.A2(n_176),
.B1(n_199),
.B2(n_168),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_234),
.A2(n_169),
.B(n_212),
.Y(n_297)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_297),
.A2(n_300),
.B(n_320),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_274),
.A2(n_225),
.B1(n_175),
.B2(n_220),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_252),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_299),
.B(n_302),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_254),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_278),
.A2(n_200),
.B1(n_185),
.B2(n_222),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_305),
.A2(n_316),
.B1(n_325),
.B2(n_14),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_239),
.Y(n_306)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_306),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_252),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_307),
.B(n_318),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_246),
.B(n_174),
.C(n_43),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_309),
.C(n_263),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_256),
.B(n_43),
.C(n_19),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_242),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_310),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_281),
.B(n_43),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_312),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_257),
.A2(n_12),
.B1(n_17),
.B2(n_16),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_237),
.B(n_0),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_315),
.B(n_317),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_274),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_230),
.B(n_12),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_276),
.Y(n_318)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_277),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_327),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_268),
.B(n_1),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_328),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_274),
.A2(n_6),
.B1(n_17),
.B2(n_3),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_242),
.Y(n_323)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_270),
.A2(n_13),
.B(n_15),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_275),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_L g326 ( 
.A1(n_262),
.A2(n_13),
.B(n_15),
.C(n_4),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_326),
.A2(n_273),
.B(n_269),
.Y(n_348)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_249),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_263),
.B(n_1),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_231),
.B(n_5),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_329),
.B(n_328),
.Y(n_372)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_271),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_273),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_361),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_289),
.A2(n_275),
.B1(n_280),
.B2(n_243),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_336),
.A2(n_338),
.B1(n_340),
.B2(n_346),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_290),
.B(n_266),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_337),
.B(n_351),
.C(n_355),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_289),
.A2(n_275),
.B1(n_280),
.B2(n_279),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_294),
.A2(n_279),
.B1(n_232),
.B2(n_260),
.Y(n_340)
);

NAND3xp33_ASAP7_75t_L g341 ( 
.A(n_315),
.B(n_267),
.C(n_239),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_341),
.B(n_368),
.Y(n_395)
);

NOR2x1_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_267),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_353),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_345),
.Y(n_374)
);

OAI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_304),
.A2(n_240),
.B1(n_255),
.B2(n_249),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_296),
.B(n_259),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_347),
.B(n_354),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_348),
.A2(n_324),
.B(n_298),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_290),
.B(n_269),
.C(n_259),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_301),
.B(n_251),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_317),
.B(n_240),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_308),
.B(n_251),
.C(n_255),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_283),
.B(n_5),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_367),
.C(n_326),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_283),
.B(n_13),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_294),
.A2(n_2),
.B1(n_14),
.B2(n_18),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_366),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_364),
.A2(n_314),
.B1(n_329),
.B2(n_306),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_365),
.A2(n_286),
.B(n_326),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_293),
.A2(n_18),
.B1(n_322),
.B2(n_301),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_283),
.B(n_18),
.C(n_309),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_312),
.Y(n_368)
);

AO21x2_ASAP7_75t_SL g370 ( 
.A1(n_300),
.A2(n_18),
.B(n_297),
.Y(n_370)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_313),
.B(n_321),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_371),
.B(n_310),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_288),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_376),
.A2(n_388),
.B(n_365),
.Y(n_425)
);

OAI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_370),
.A2(n_333),
.B1(n_339),
.B2(n_334),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_377),
.A2(n_392),
.B1(n_332),
.B2(n_343),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_358),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_378),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_342),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_379),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_381),
.B(n_397),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_337),
.B(n_313),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_382),
.B(n_394),
.C(n_401),
.Y(n_415)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_363),
.Y(n_385)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_385),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_371),
.B(n_288),
.Y(n_386)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_386),
.Y(n_434)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_363),
.Y(n_387)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_387),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_356),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_389),
.B(n_396),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_333),
.A2(n_303),
.B1(n_316),
.B2(n_305),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_390),
.A2(n_405),
.B(n_362),
.Y(n_433)
);

OAI22x1_ASAP7_75t_SL g391 ( 
.A1(n_370),
.A2(n_300),
.B1(n_320),
.B2(n_288),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_391),
.A2(n_402),
.B1(n_390),
.B2(n_405),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_351),
.B(n_335),
.C(n_355),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_357),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_360),
.B(n_311),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_399),
.Y(n_422)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_349),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_400),
.B(n_403),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_367),
.B(n_302),
.C(n_299),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_334),
.A2(n_300),
.B1(n_306),
.B2(n_327),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_331),
.B(n_307),
.C(n_285),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_336),
.C(n_338),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_332),
.A2(n_325),
.B1(n_330),
.B2(n_310),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_406),
.B(n_408),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_356),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_323),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_357),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_409),
.A2(n_427),
.B1(n_398),
.B2(n_376),
.Y(n_443)
);

MAJx2_ASAP7_75t_L g410 ( 
.A(n_380),
.B(n_344),
.C(n_359),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_414),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_384),
.A2(n_331),
.B1(n_350),
.B2(n_364),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_413),
.A2(n_419),
.B1(n_433),
.B2(n_392),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_380),
.B(n_361),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_416),
.B(n_431),
.Y(n_460)
);

BUFx24_ASAP7_75t_SL g417 ( 
.A(n_378),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_417),
.B(n_395),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_394),
.B(n_359),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_421),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_382),
.B(n_353),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_366),
.Y(n_423)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_423),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_425),
.A2(n_370),
.B(n_383),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_375),
.B(n_372),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_438),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_388),
.A2(n_384),
.B1(n_391),
.B2(n_343),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_375),
.B(n_350),
.C(n_340),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_429),
.C(n_430),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_368),
.C(n_348),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_401),
.B(n_352),
.C(n_339),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_373),
.B(n_339),
.Y(n_431)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_373),
.B(n_352),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_381),
.B(n_370),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_439),
.B(n_386),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_420),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_441),
.B(n_448),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_443),
.A2(n_433),
.B1(n_413),
.B2(n_431),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_440),
.B(n_379),
.Y(n_445)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_445),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_435),
.B(n_374),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_449),
.B(n_465),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_420),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_450),
.B(n_452),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_451),
.A2(n_425),
.B1(n_439),
.B2(n_422),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_374),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_453),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_418),
.B(n_393),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_454),
.B(n_426),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_415),
.B(n_404),
.C(n_408),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_455),
.B(n_459),
.C(n_461),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_424),
.B(n_398),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_456),
.B(n_428),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_423),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_457),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_415),
.B(n_396),
.C(n_400),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_424),
.B(n_399),
.C(n_385),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_411),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_463),
.Y(n_473)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_412),
.Y(n_464)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_464),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_434),
.B(n_387),
.Y(n_466)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_466),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_414),
.B(n_383),
.C(n_389),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_467),
.B(n_461),
.C(n_449),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_468),
.B(n_481),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_445),
.A2(n_416),
.B(n_411),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_469),
.A2(n_467),
.B(n_451),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_430),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_483),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_446),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_436),
.Y(n_478)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_478),
.Y(n_495)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_464),
.Y(n_480)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_480),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_458),
.A2(n_409),
.B1(n_427),
.B2(n_421),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_429),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_484),
.B(n_444),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_485),
.B(n_487),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_459),
.B(n_407),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_488),
.B(n_466),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_475),
.B(n_462),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_490),
.B(n_498),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_491),
.B(n_501),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_486),
.B(n_476),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_493),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_497),
.Y(n_522)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_470),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_468),
.A2(n_465),
.B(n_481),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_499),
.A2(n_506),
.B(n_482),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_479),
.B(n_455),
.C(n_444),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_505),
.C(n_483),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_473),
.B(n_462),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_503),
.B(n_504),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_479),
.B(n_456),
.C(n_446),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_472),
.B(n_438),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_484),
.B(n_474),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_507),
.B(n_442),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_501),
.A2(n_485),
.B1(n_472),
.B2(n_482),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_508),
.B(n_513),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_491),
.B(n_477),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_509),
.B(n_516),
.C(n_505),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_500),
.A2(n_475),
.B(n_489),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_510),
.B(n_504),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_512),
.B(n_515),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_499),
.B(n_478),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_469),
.C(n_442),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_518),
.A2(n_494),
.B(n_502),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_493),
.B(n_480),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_519),
.B(n_521),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_495),
.B(n_470),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_523),
.B(n_524),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_511),
.A2(n_502),
.B(n_496),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_526),
.B(n_531),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_529),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_514),
.B(n_506),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_512),
.A2(n_492),
.B(n_471),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_522),
.B(n_492),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_532),
.B(n_533),
.Y(n_537)
);

AOI21x1_ASAP7_75t_SL g533 ( 
.A1(n_513),
.A2(n_518),
.B(n_508),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_525),
.B(n_520),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_536),
.B(n_539),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_523),
.B(n_516),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_527),
.B(n_521),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_540),
.A2(n_533),
.B(n_521),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_534),
.B(n_517),
.C(n_527),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_541),
.B(n_542),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_538),
.B(n_530),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_544),
.B(n_538),
.C(n_535),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_545),
.B(n_517),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_546),
.A2(n_543),
.B(n_537),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_547),
.A2(n_548),
.B(n_369),
.Y(n_549)
);

AO21x1_ASAP7_75t_SL g550 ( 
.A1(n_549),
.A2(n_471),
.B(n_410),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_550),
.A2(n_447),
.B(n_509),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_551),
.A2(n_447),
.B1(n_369),
.B2(n_323),
.Y(n_552)
);


endmodule