module fake_netlist_6_4555_n_1471 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1471);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1471;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_873;
wire n_461;
wire n_383;
wire n_1371;
wire n_1285;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_474;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_934;
wire n_482;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1147;
wire n_763;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_151),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_160),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_248),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_156),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_62),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_110),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_327),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_291),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_54),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_107),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_149),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_77),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_62),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_217),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_315),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_229),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_49),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_16),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_17),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_314),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_9),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_63),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_164),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_48),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_220),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_87),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_312),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_213),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_48),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_297),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_244),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_236),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_93),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_299),
.Y(n_364)
);

BUFx10_ASAP7_75t_L g365 ( 
.A(n_324),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_232),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_61),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_296),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_174),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_185),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_172),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_58),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_72),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_88),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_36),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_198),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_22),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_308),
.Y(n_378)
);

BUFx10_ASAP7_75t_L g379 ( 
.A(n_11),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_233),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_246),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_139),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_306),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_279),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_91),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_219),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_184),
.Y(n_387)
);

BUFx5_ASAP7_75t_L g388 ( 
.A(n_176),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_133),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_228),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_69),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_289),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_128),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_165),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_266),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_147),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_117),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_58),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_209),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_19),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_34),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_240),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_134),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_283),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_158),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_215),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_47),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_225),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_80),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_140),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_43),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_274),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_12),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_138),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_27),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_221),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_86),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_169),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_325),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_54),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_59),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_258),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_326),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_261),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_8),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_92),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_153),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_284),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_115),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_135),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_292),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_241),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_304),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_74),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_317),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_146),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_187),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_309),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_237),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_33),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_59),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_273),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_286),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_145),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_192),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_260),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_76),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_264),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_263),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_269),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_2),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_239),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_242),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_212),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_250),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_216),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_132),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_214),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_210),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_318),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_302),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_17),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_166),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_222),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_159),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_98),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_32),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_114),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_202),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_111),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_63),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_109),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_301),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_226),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_21),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_319),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_25),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_28),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_4),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_254),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_19),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_180),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_265),
.Y(n_483)
);

BUFx8_ASAP7_75t_SL g484 ( 
.A(n_157),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_189),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_257),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_282),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_205),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_124),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_154),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_194),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_295),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_34),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_141),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_256),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_101),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_253),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_230),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_5),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_251),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_227),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_208),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_90),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_290),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_22),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_99),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_293),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_275),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_37),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_79),
.Y(n_510)
);

BUFx5_ASAP7_75t_L g511 ( 
.A(n_16),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_211),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_199),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_44),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_168),
.Y(n_515)
);

BUFx5_ASAP7_75t_L g516 ( 
.A(n_173),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_6),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_50),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_94),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_223),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_60),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_47),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_333),
.Y(n_523)
);

INVxp33_ASAP7_75t_SL g524 ( 
.A(n_352),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_478),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_330),
.Y(n_526)
);

INVxp67_ASAP7_75t_SL g527 ( 
.A(n_437),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_511),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_511),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_427),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_478),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_372),
.Y(n_532)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_427),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_511),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_511),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_511),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_334),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_347),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_511),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_511),
.Y(n_540)
);

INVxp33_ASAP7_75t_L g541 ( 
.A(n_339),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_349),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_379),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_332),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_354),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_354),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_379),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_338),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_340),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_411),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_411),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_379),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_446),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_425),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g555 ( 
.A(n_446),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_382),
.B(n_0),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_341),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_425),
.Y(n_558)
);

INVx4_ASAP7_75t_R g559 ( 
.A(n_488),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_421),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_345),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_356),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_382),
.B(n_0),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_353),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g565 ( 
.A(n_488),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_343),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_416),
.B(n_1),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_485),
.B(n_1),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_485),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_368),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_348),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_357),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_351),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_367),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_377),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_359),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_358),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_413),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_420),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_477),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_388),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_479),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_388),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_363),
.Y(n_584)
);

INVxp67_ASAP7_75t_SL g585 ( 
.A(n_519),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_376),
.B(n_2),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_481),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_493),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_356),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_364),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_509),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_500),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_514),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_521),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_522),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_335),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_337),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_388),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_344),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_350),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_458),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_366),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_355),
.Y(n_603)
);

CKINVDCx16_ASAP7_75t_R g604 ( 
.A(n_458),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_470),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_360),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_369),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_388),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_361),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_362),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_378),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_375),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_371),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_506),
.B(n_3),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_398),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_383),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_470),
.Y(n_617)
);

INVxp67_ASAP7_75t_SL g618 ( 
.A(n_385),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_386),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_513),
.B(n_3),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_387),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_373),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_389),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_400),
.Y(n_624)
);

BUFx6f_ASAP7_75t_SL g625 ( 
.A(n_365),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_512),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_390),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_512),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_391),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_374),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_380),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_394),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_515),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_515),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_401),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_381),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_388),
.Y(n_637)
);

CKINVDCx16_ASAP7_75t_R g638 ( 
.A(n_365),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_596),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_526),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_563),
.B(n_567),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_569),
.B(n_331),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_597),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_599),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_528),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_600),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_544),
.B(n_331),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_548),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_549),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_529),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_557),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_618),
.B(n_342),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_603),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_606),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_545),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_534),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_562),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_609),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_627),
.B(n_342),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_562),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_561),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_537),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_535),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_610),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_R g665 ( 
.A(n_537),
.B(n_407),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_611),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_532),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_564),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_572),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_530),
.B(n_346),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_538),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_616),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_619),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_536),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_615),
.B(n_365),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_577),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_589),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_584),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_621),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_539),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_623),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_589),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_540),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_566),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_581),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_601),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_635),
.B(n_448),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_533),
.B(n_346),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_629),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_553),
.B(n_555),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_632),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_590),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_571),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_581),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_527),
.B(n_448),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_573),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_575),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_579),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_624),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_602),
.B(n_370),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_580),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_607),
.B(n_370),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_565),
.B(n_448),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_613),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_622),
.B(n_418),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_582),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_620),
.B(n_418),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_630),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_524),
.A2(n_440),
.B1(n_441),
.B2(n_415),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_570),
.B(n_336),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_587),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_583),
.Y(n_712)
);

OAI21x1_ASAP7_75t_L g713 ( 
.A1(n_583),
.A2(n_608),
.B(n_598),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_585),
.B(n_444),
.Y(n_714)
);

CKINVDCx16_ASAP7_75t_R g715 ( 
.A(n_604),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_588),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_546),
.B(n_444),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_601),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_605),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_598),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_631),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_605),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_636),
.B(n_452),
.Y(n_723)
);

INVxp33_ASAP7_75t_SL g724 ( 
.A(n_538),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_556),
.B(n_395),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_591),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_617),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_542),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_684),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_713),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_645),
.B(n_650),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_707),
.A2(n_568),
.B1(n_614),
.B2(n_586),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_710),
.B(n_592),
.Y(n_733)
);

AOI22x1_ASAP7_75t_L g734 ( 
.A1(n_707),
.A2(n_523),
.B1(n_576),
.B2(n_542),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_645),
.B(n_608),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_725),
.B(n_638),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_725),
.B(n_576),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_690),
.B(n_612),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_647),
.B(n_612),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_700),
.B(n_524),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_667),
.B(n_543),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_693),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_702),
.B(n_625),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_684),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_696),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_690),
.B(n_547),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_650),
.B(n_637),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_684),
.Y(n_748)
);

CKINVDCx8_ASAP7_75t_R g749 ( 
.A(n_715),
.Y(n_749)
);

CKINVDCx12_ASAP7_75t_R g750 ( 
.A(n_675),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_656),
.B(n_637),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_690),
.B(n_552),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_642),
.B(n_550),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_655),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_R g755 ( 
.A(n_728),
.B(n_551),
.Y(n_755)
);

AND2x2_ASAP7_75t_SL g756 ( 
.A(n_662),
.B(n_452),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_697),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_684),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_705),
.B(n_554),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_698),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_698),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_657),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_656),
.B(n_388),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_663),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_642),
.B(n_558),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_663),
.B(n_674),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_706),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_674),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_723),
.B(n_625),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_680),
.Y(n_770)
);

NAND3xp33_ASAP7_75t_L g771 ( 
.A(n_641),
.B(n_578),
.C(n_574),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_716),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_726),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_703),
.B(n_541),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_SL g775 ( 
.A1(n_727),
.A2(n_626),
.B1(n_628),
.B2(n_617),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_698),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_642),
.B(n_593),
.Y(n_777)
);

INVxp33_ASAP7_75t_SL g778 ( 
.A(n_640),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_680),
.B(n_388),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_639),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_641),
.A2(n_625),
.B1(n_468),
.B2(n_472),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_643),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_687),
.B(n_384),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_648),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_695),
.B(n_541),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_699),
.B(n_594),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_655),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_677),
.Y(n_788)
);

INVxp67_ASAP7_75t_SL g789 ( 
.A(n_685),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_686),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_707),
.B(n_595),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_698),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_644),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_646),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_683),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_714),
.B(n_652),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_671),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_683),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_685),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_694),
.B(n_712),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_670),
.B(n_396),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_670),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_694),
.Y(n_803)
);

NAND3xp33_ASAP7_75t_L g804 ( 
.A(n_665),
.B(n_709),
.C(n_714),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_670),
.Y(n_805)
);

AND2x2_ASAP7_75t_SL g806 ( 
.A(n_714),
.B(n_496),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_653),
.Y(n_807)
);

AND2x2_ASAP7_75t_SL g808 ( 
.A(n_652),
.B(n_496),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_688),
.B(n_429),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_688),
.Y(n_810)
);

INVx5_ASAP7_75t_L g811 ( 
.A(n_712),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_654),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_688),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_652),
.Y(n_814)
);

AND2x6_ASAP7_75t_L g815 ( 
.A(n_659),
.B(n_397),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_720),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_717),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_808),
.B(n_659),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_797),
.B(n_717),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_737),
.B(n_724),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_806),
.B(n_756),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_802),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_814),
.B(n_659),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_733),
.Y(n_824)
);

NOR2xp67_ASAP7_75t_L g825 ( 
.A(n_784),
.B(n_649),
.Y(n_825)
);

OAI22xp33_ASAP7_75t_L g826 ( 
.A1(n_813),
.A2(n_462),
.B1(n_475),
.B2(n_665),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_737),
.B(n_651),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_814),
.B(n_661),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_810),
.B(n_668),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_799),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_799),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_785),
.B(n_669),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_732),
.A2(n_796),
.B1(n_804),
.B2(n_815),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_740),
.B(n_676),
.Y(n_834)
);

AND3x1_ASAP7_75t_L g835 ( 
.A(n_740),
.B(n_739),
.C(n_781),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_805),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_803),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_742),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_817),
.Y(n_839)
);

AND3x1_ASAP7_75t_L g840 ( 
.A(n_739),
.B(n_711),
.C(n_701),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_810),
.B(n_678),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_774),
.B(n_692),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_746),
.B(n_704),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_809),
.B(n_708),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_789),
.A2(n_720),
.B(n_664),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_752),
.B(n_721),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_809),
.B(n_658),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_816),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_789),
.B(n_791),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_788),
.Y(n_850)
);

BUFx5_ASAP7_75t_L g851 ( 
.A(n_815),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_732),
.A2(n_815),
.B1(n_801),
.B2(n_791),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_786),
.B(n_717),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_736),
.B(n_666),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_815),
.A2(n_414),
.B1(n_417),
.B2(n_403),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_817),
.B(n_672),
.Y(n_856)
);

NAND2xp33_ASAP7_75t_L g857 ( 
.A(n_817),
.B(n_516),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_738),
.B(n_673),
.Y(n_858)
);

AND3x1_ASAP7_75t_L g859 ( 
.A(n_743),
.B(n_711),
.C(n_701),
.Y(n_859)
);

NAND2xp33_ASAP7_75t_SL g860 ( 
.A(n_755),
.B(n_626),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_777),
.B(n_679),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_787),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_777),
.B(n_681),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_743),
.B(n_392),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_745),
.B(n_689),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_757),
.B(n_691),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_759),
.B(n_451),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_769),
.B(n_393),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_767),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_772),
.B(n_419),
.Y(n_870)
);

OAI22xp33_ASAP7_75t_L g871 ( 
.A1(n_771),
.A2(n_471),
.B1(n_499),
.B2(n_467),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_764),
.Y(n_872)
);

O2A1O1Ixp5_ASAP7_75t_L g873 ( 
.A1(n_801),
.A2(n_428),
.B(n_432),
.C(n_422),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_768),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_769),
.B(n_399),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_773),
.B(n_433),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_780),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_770),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_787),
.B(n_628),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_782),
.B(n_436),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_753),
.B(n_765),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_753),
.A2(n_765),
.B1(n_755),
.B2(n_750),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_754),
.B(n_633),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_793),
.B(n_505),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_794),
.B(n_517),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_783),
.A2(n_730),
.B1(n_734),
.B2(n_807),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_812),
.B(n_445),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_729),
.B(n_447),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_795),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_798),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_730),
.A2(n_454),
.B1(n_455),
.B2(n_449),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_729),
.B(n_761),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_800),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_800),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_731),
.Y(n_895)
);

BUFx8_ASAP7_75t_L g896 ( 
.A(n_762),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_741),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_790),
.B(n_633),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_761),
.B(n_792),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_731),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_766),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_730),
.Y(n_902)
);

NAND3xp33_ASAP7_75t_L g903 ( 
.A(n_766),
.B(n_518),
.C(n_404),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_778),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_792),
.B(n_456),
.Y(n_905)
);

NOR2x1p5_ASAP7_75t_L g906 ( 
.A(n_749),
.B(n_402),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_763),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_744),
.B(n_466),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_744),
.B(n_748),
.Y(n_909)
);

NOR2x1p5_ASAP7_75t_L g910 ( 
.A(n_763),
.B(n_405),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_790),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_744),
.B(n_483),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_735),
.A2(n_487),
.B1(n_492),
.B2(n_489),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_895),
.A2(n_747),
.B(n_751),
.C(n_735),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_879),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_867),
.B(n_634),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_900),
.B(n_747),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_837),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_839),
.Y(n_919)
);

AND3x1_ASAP7_75t_L g920 ( 
.A(n_820),
.B(n_560),
.C(n_531),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_839),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_911),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_901),
.B(n_751),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_836),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_836),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_862),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_904),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_867),
.B(n_634),
.Y(n_928)
);

NOR3xp33_ASAP7_75t_SL g929 ( 
.A(n_826),
.B(n_775),
.C(n_408),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_839),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_823),
.A2(n_779),
.B(n_758),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_834),
.B(n_560),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_839),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_893),
.B(n_779),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_838),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_869),
.Y(n_936)
);

INVxp67_ASAP7_75t_SL g937 ( 
.A(n_902),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_848),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_850),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_872),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_894),
.A2(n_516),
.B1(n_503),
.B2(n_508),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_822),
.B(n_748),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_907),
.B(n_748),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_849),
.B(n_852),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_835),
.A2(n_760),
.B1(n_776),
.B2(n_758),
.Y(n_945)
);

NAND2xp33_ASAP7_75t_SL g946 ( 
.A(n_821),
.B(n_719),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_852),
.B(n_758),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_874),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_878),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_881),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_843),
.B(n_846),
.Y(n_951)
);

INVx5_ASAP7_75t_L g952 ( 
.A(n_819),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_877),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_889),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_890),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_898),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_833),
.B(n_760),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_853),
.B(n_760),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_830),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_827),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_862),
.Y(n_961)
);

INVx6_ASAP7_75t_L g962 ( 
.A(n_896),
.Y(n_962)
);

AND3x2_ASAP7_75t_SL g963 ( 
.A(n_826),
.B(n_531),
.C(n_525),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_818),
.A2(n_776),
.B1(n_409),
.B2(n_410),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_883),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_831),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_910),
.B(n_776),
.Y(n_967)
);

BUFx2_ASAP7_75t_SL g968 ( 
.A(n_825),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_833),
.B(n_811),
.Y(n_969)
);

OAI21xp33_ASAP7_75t_L g970 ( 
.A1(n_820),
.A2(n_834),
.B(n_827),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_824),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_856),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_858),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_819),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_847),
.B(n_811),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_882),
.A2(n_525),
.B1(n_412),
.B2(n_423),
.Y(n_976)
);

BUFx8_ASAP7_75t_L g977 ( 
.A(n_832),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_896),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_897),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_861),
.B(n_722),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_863),
.B(n_657),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_858),
.B(n_811),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_909),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_860),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_819),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_865),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_843),
.B(n_846),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_892),
.Y(n_988)
);

OR2x2_ASAP7_75t_SL g989 ( 
.A(n_828),
.B(n_660),
.Y(n_989)
);

INVx4_ASAP7_75t_L g990 ( 
.A(n_851),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_844),
.B(n_660),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_916),
.B(n_842),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_931),
.A2(n_899),
.B(n_886),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_944),
.A2(n_957),
.B(n_947),
.Y(n_994)
);

OR2x4_ASAP7_75t_L g995 ( 
.A(n_991),
.B(n_842),
.Y(n_995)
);

BUFx12f_ASAP7_75t_L g996 ( 
.A(n_962),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_918),
.Y(n_997)
);

BUFx4_ASAP7_75t_SL g998 ( 
.A(n_978),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_944),
.B(n_854),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_970),
.A2(n_854),
.B(n_885),
.C(n_884),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_917),
.B(n_829),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_917),
.B(n_841),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_951),
.B(n_987),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_L g1004 ( 
.A1(n_931),
.A2(n_905),
.B(n_888),
.Y(n_1004)
);

OAI21x1_ASAP7_75t_L g1005 ( 
.A1(n_914),
.A2(n_845),
.B(n_908),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_914),
.A2(n_912),
.B(n_873),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_943),
.A2(n_969),
.B(n_988),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_943),
.A2(n_859),
.B(n_840),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_980),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_928),
.B(n_884),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_969),
.A2(n_947),
.B(n_983),
.Y(n_1011)
);

O2A1O1Ixp5_ASAP7_75t_L g1012 ( 
.A1(n_982),
.A2(n_864),
.B(n_875),
.C(n_868),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_990),
.A2(n_934),
.B(n_923),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_923),
.B(n_866),
.Y(n_1014)
);

O2A1O1Ixp5_ASAP7_75t_L g1015 ( 
.A1(n_982),
.A2(n_891),
.B(n_870),
.C(n_880),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_935),
.Y(n_1016)
);

AO31x2_ASAP7_75t_L g1017 ( 
.A1(n_957),
.A2(n_975),
.A3(n_934),
.B(n_972),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_973),
.B(n_876),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_956),
.B(n_965),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_936),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_973),
.B(n_887),
.Y(n_1021)
);

AOI211x1_ASAP7_75t_L g1022 ( 
.A1(n_986),
.A2(n_871),
.B(n_903),
.C(n_913),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_960),
.A2(n_929),
.B1(n_941),
.B2(n_855),
.Y(n_1023)
);

OA22x2_ASAP7_75t_L g1024 ( 
.A1(n_963),
.A2(n_871),
.B1(n_906),
.B2(n_718),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_953),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_990),
.A2(n_855),
.B(n_857),
.Y(n_1026)
);

NAND2xp33_ASAP7_75t_L g1027 ( 
.A(n_921),
.B(n_851),
.Y(n_1027)
);

O2A1O1Ixp5_ASAP7_75t_L g1028 ( 
.A1(n_975),
.A2(n_885),
.B(n_851),
.C(n_913),
.Y(n_1028)
);

AO21x1_ASAP7_75t_L g1029 ( 
.A1(n_945),
.A2(n_937),
.B(n_946),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_932),
.B(n_682),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_926),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_955),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_958),
.B(n_851),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_926),
.B(n_682),
.Y(n_1034)
);

NAND2x1p5_ASAP7_75t_L g1035 ( 
.A(n_921),
.B(n_811),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_941),
.A2(n_424),
.B(n_406),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_937),
.A2(n_851),
.B(n_430),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_919),
.A2(n_851),
.B(n_516),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_919),
.A2(n_516),
.B(n_70),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_961),
.B(n_718),
.Y(n_1040)
);

NOR2xp67_ASAP7_75t_SL g1041 ( 
.A(n_968),
.B(n_426),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_958),
.A2(n_434),
.B(n_431),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_950),
.B(n_727),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_930),
.A2(n_516),
.B(n_71),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_971),
.B(n_435),
.Y(n_1045)
);

AOI21x1_ASAP7_75t_L g1046 ( 
.A1(n_938),
.A2(n_516),
.B(n_559),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_930),
.A2(n_966),
.B(n_959),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_961),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_959),
.A2(n_966),
.B(n_940),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_940),
.A2(n_516),
.B(n_73),
.Y(n_1050)
);

OAI22x1_ASAP7_75t_L g1051 ( 
.A1(n_963),
.A2(n_439),
.B1(n_442),
.B2(n_438),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_921),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_SL g1053 ( 
.A1(n_974),
.A2(n_75),
.B(n_68),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_950),
.B(n_443),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_971),
.B(n_450),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_948),
.A2(n_81),
.B(n_78),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_949),
.A2(n_83),
.B(n_82),
.Y(n_1057)
);

AOI31xp33_ASAP7_75t_L g1058 ( 
.A1(n_920),
.A2(n_939),
.A3(n_976),
.B(n_981),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_954),
.A2(n_457),
.B(n_453),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_SL g1060 ( 
.A1(n_974),
.A2(n_85),
.B(n_84),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_915),
.B(n_459),
.Y(n_1061)
);

BUFx4f_ASAP7_75t_L g1062 ( 
.A(n_962),
.Y(n_1062)
);

OA21x2_ASAP7_75t_L g1063 ( 
.A1(n_1028),
.A2(n_964),
.B(n_984),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1011),
.Y(n_1064)
);

OA21x2_ASAP7_75t_L g1065 ( 
.A1(n_1006),
.A2(n_942),
.B(n_929),
.Y(n_1065)
);

AO31x2_ASAP7_75t_L g1066 ( 
.A1(n_1000),
.A2(n_925),
.A3(n_924),
.B(n_989),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1016),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_1014),
.A2(n_967),
.B(n_950),
.C(n_981),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1020),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_1014),
.A2(n_952),
.B1(n_933),
.B2(n_980),
.Y(n_1070)
);

OAI221xp5_ASAP7_75t_L g1071 ( 
.A1(n_1030),
.A2(n_922),
.B1(n_979),
.B2(n_927),
.C(n_985),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1025),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1007),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1001),
.B(n_967),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1001),
.B(n_942),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_1019),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1013),
.A2(n_933),
.B(n_952),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_SL g1078 ( 
.A1(n_1029),
.A2(n_952),
.B(n_933),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1032),
.Y(n_1079)
);

OR2x6_ASAP7_75t_L g1080 ( 
.A(n_994),
.B(n_985),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_SL g1081 ( 
.A1(n_1053),
.A2(n_952),
.B(n_977),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_1031),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1002),
.B(n_985),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1049),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_1038),
.A2(n_977),
.B(n_95),
.Y(n_1085)
);

OR2x2_ASAP7_75t_L g1086 ( 
.A(n_992),
.B(n_460),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1017),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_999),
.B(n_962),
.Y(n_1088)
);

BUFx8_ASAP7_75t_SL g1089 ( 
.A(n_996),
.Y(n_1089)
);

BUFx10_ASAP7_75t_L g1090 ( 
.A(n_1034),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_993),
.A2(n_96),
.B(n_89),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_997),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1004),
.A2(n_100),
.B(n_97),
.Y(n_1093)
);

AND2x4_ASAP7_75t_SL g1094 ( 
.A(n_1048),
.B(n_484),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1024),
.A2(n_484),
.B1(n_510),
.B2(n_507),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1024),
.A2(n_520),
.B1(n_504),
.B2(n_502),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_1010),
.B(n_461),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1017),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_998),
.Y(n_1099)
);

CKINVDCx11_ASAP7_75t_R g1100 ( 
.A(n_1043),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_1009),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1017),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1047),
.A2(n_103),
.B(n_102),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_1043),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1005),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1002),
.A2(n_464),
.B(n_463),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1040),
.A2(n_501),
.B1(n_498),
.B2(n_497),
.Y(n_1107)
);

AO31x2_ASAP7_75t_L g1108 ( 
.A1(n_999),
.A2(n_4),
.A3(n_5),
.B(n_6),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1056),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_994),
.B(n_465),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1018),
.Y(n_1111)
);

INVxp67_ASAP7_75t_L g1112 ( 
.A(n_1045),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1018),
.B(n_469),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1021),
.B(n_473),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1021),
.B(n_474),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1003),
.B(n_104),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_995),
.B(n_476),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1033),
.B(n_105),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1052),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1057),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1026),
.A2(n_495),
.B(n_482),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1026),
.A2(n_1027),
.B(n_1037),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1008),
.B(n_480),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_1062),
.Y(n_1124)
);

AOI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1046),
.A2(n_490),
.B(n_486),
.Y(n_1125)
);

BUFx12f_ASAP7_75t_L g1126 ( 
.A(n_1061),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_1062),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1022),
.B(n_995),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1128),
.A2(n_1023),
.B1(n_1051),
.B2(n_1036),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1067),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1067),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1072),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1112),
.A2(n_1058),
.B1(n_1023),
.B2(n_1054),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_SL g1134 ( 
.A1(n_1116),
.A2(n_1058),
.B1(n_1055),
.B2(n_1042),
.Y(n_1134)
);

NAND3xp33_ASAP7_75t_SL g1135 ( 
.A(n_1096),
.B(n_1012),
.C(n_1015),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1115),
.B(n_1042),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1072),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1074),
.A2(n_1036),
.B1(n_1033),
.B2(n_1059),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1118),
.Y(n_1139)
);

OAI221xp5_ASAP7_75t_L g1140 ( 
.A1(n_1095),
.A2(n_1059),
.B1(n_1041),
.B2(n_1037),
.C(n_491),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1115),
.B(n_1052),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_1099),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1116),
.A2(n_1060),
.B1(n_1044),
.B2(n_1039),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1069),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1116),
.A2(n_1050),
.B1(n_494),
.B2(n_1035),
.Y(n_1145)
);

O2A1O1Ixp5_ASAP7_75t_L g1146 ( 
.A1(n_1122),
.A2(n_1035),
.B(n_8),
.C(n_9),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1111),
.B(n_7),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1104),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1088),
.B(n_1097),
.Y(n_1149)
);

AND2x2_ASAP7_75t_SL g1150 ( 
.A(n_1110),
.B(n_7),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1121),
.A2(n_10),
.B(n_11),
.Y(n_1151)
);

AND3x1_ASAP7_75t_L g1152 ( 
.A(n_1117),
.B(n_10),
.C(n_12),
.Y(n_1152)
);

INVxp33_ASAP7_75t_SL g1153 ( 
.A(n_1099),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1076),
.B(n_13),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1071),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_1155)
);

INVxp33_ASAP7_75t_L g1156 ( 
.A(n_1101),
.Y(n_1156)
);

CKINVDCx8_ASAP7_75t_R g1157 ( 
.A(n_1124),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1088),
.B(n_1083),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1092),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1079),
.Y(n_1160)
);

OAI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1075),
.A2(n_14),
.B1(n_15),
.B2(n_18),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_SL g1162 ( 
.A1(n_1068),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1082),
.Y(n_1163)
);

NAND3x1_ASAP7_75t_L g1164 ( 
.A(n_1107),
.B(n_20),
.C(n_23),
.Y(n_1164)
);

CKINVDCx6p67_ASAP7_75t_R g1165 ( 
.A(n_1127),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1082),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_SL g1167 ( 
.A1(n_1110),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1086),
.B(n_24),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1118),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1126),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1068),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1118),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1070),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_1127),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1113),
.B(n_31),
.Y(n_1175)
);

CKINVDCx6p67_ASAP7_75t_R g1176 ( 
.A(n_1126),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1080),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1114),
.B(n_32),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1124),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_SL g1180 ( 
.A1(n_1077),
.A2(n_33),
.B(n_35),
.C(n_36),
.Y(n_1180)
);

OAI221xp5_ASAP7_75t_L g1181 ( 
.A1(n_1106),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.C(n_39),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1090),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1066),
.B(n_40),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1066),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1066),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_1123),
.B(n_41),
.C(n_42),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1090),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1080),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1080),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1066),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1089),
.Y(n_1191)
);

AOI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1125),
.A2(n_190),
.B(n_328),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1089),
.Y(n_1193)
);

INVx6_ASAP7_75t_L g1194 ( 
.A(n_1090),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1150),
.A2(n_1123),
.B1(n_1080),
.B2(n_1100),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1150),
.A2(n_1100),
.B1(n_1081),
.B2(n_1065),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1181),
.A2(n_1065),
.B1(n_1063),
.B2(n_1078),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1158),
.B(n_1108),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1184),
.A2(n_1105),
.A3(n_1073),
.B(n_1064),
.Y(n_1199)
);

CKINVDCx11_ASAP7_75t_R g1200 ( 
.A(n_1142),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1133),
.A2(n_1065),
.B1(n_1063),
.B2(n_1119),
.Y(n_1201)
);

AO21x1_ASAP7_75t_L g1202 ( 
.A1(n_1188),
.A2(n_1087),
.B(n_1102),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1129),
.A2(n_1134),
.B1(n_1182),
.B2(n_1170),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1186),
.A2(n_1063),
.B1(n_1094),
.B2(n_1087),
.Y(n_1204)
);

OAI222xp33_ASAP7_75t_L g1205 ( 
.A1(n_1167),
.A2(n_1182),
.B1(n_1187),
.B2(n_1155),
.C1(n_1171),
.C2(n_1129),
.Y(n_1205)
);

AOI21xp33_ASAP7_75t_L g1206 ( 
.A1(n_1136),
.A2(n_1064),
.B(n_1073),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_SL g1207 ( 
.A1(n_1151),
.A2(n_1094),
.B1(n_1085),
.B2(n_1091),
.Y(n_1207)
);

AOI222xp33_ASAP7_75t_L g1208 ( 
.A1(n_1161),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.C1(n_53),
.C2(n_55),
.Y(n_1208)
);

OAI211xp5_ASAP7_75t_L g1209 ( 
.A1(n_1167),
.A2(n_1102),
.B(n_1098),
.C(n_1105),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1161),
.A2(n_1098),
.B1(n_1084),
.B2(n_1109),
.Y(n_1210)
);

OAI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1188),
.A2(n_1109),
.B1(n_1120),
.B2(n_1084),
.Y(n_1211)
);

OAI33xp33_ASAP7_75t_L g1212 ( 
.A1(n_1147),
.A2(n_1108),
.A3(n_52),
.B1(n_53),
.B2(n_55),
.B3(n_56),
.Y(n_1212)
);

OAI221xp5_ASAP7_75t_L g1213 ( 
.A1(n_1152),
.A2(n_1120),
.B1(n_1108),
.B2(n_1085),
.C(n_60),
.Y(n_1213)
);

OR2x6_ASAP7_75t_L g1214 ( 
.A(n_1177),
.B(n_1093),
.Y(n_1214)
);

BUFx12f_ASAP7_75t_L g1215 ( 
.A(n_1191),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1135),
.A2(n_1091),
.B(n_1093),
.Y(n_1216)
);

OAI222xp33_ASAP7_75t_L g1217 ( 
.A1(n_1189),
.A2(n_1108),
.B1(n_56),
.B2(n_57),
.C1(n_61),
.C2(n_64),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1144),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_SL g1219 ( 
.A1(n_1178),
.A2(n_1103),
.B1(n_57),
.B2(n_64),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1149),
.A2(n_1103),
.B1(n_65),
.B2(n_66),
.Y(n_1220)
);

AOI221xp5_ASAP7_75t_L g1221 ( 
.A1(n_1173),
.A2(n_1154),
.B1(n_1180),
.B2(n_1162),
.C(n_1135),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1141),
.B(n_106),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1156),
.B(n_51),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1168),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1194),
.A2(n_67),
.B1(n_108),
.B2(n_112),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1163),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1194),
.A2(n_1164),
.B1(n_1139),
.B2(n_1175),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1160),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1130),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1177),
.B(n_113),
.Y(n_1230)
);

OAI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1176),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1156),
.B(n_120),
.Y(n_1232)
);

AND2x4_ASAP7_75t_SL g1233 ( 
.A(n_1165),
.B(n_121),
.Y(n_1233)
);

AOI221xp5_ASAP7_75t_L g1234 ( 
.A1(n_1154),
.A2(n_122),
.B1(n_123),
.B2(n_125),
.C(n_126),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1169),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_1235)
);

AOI21xp33_ASAP7_75t_L g1236 ( 
.A1(n_1140),
.A2(n_131),
.B(n_136),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1148),
.B(n_137),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1194),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1159),
.B(n_1131),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1137),
.Y(n_1240)
);

AOI221xp5_ASAP7_75t_L g1241 ( 
.A1(n_1180),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.C(n_148),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_1153),
.Y(n_1242)
);

NAND2x1_ASAP7_75t_L g1243 ( 
.A(n_1139),
.B(n_150),
.Y(n_1243)
);

AOI222xp33_ASAP7_75t_L g1244 ( 
.A1(n_1183),
.A2(n_152),
.B1(n_155),
.B2(n_161),
.C1(n_162),
.C2(n_163),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1172),
.A2(n_167),
.B1(n_170),
.B2(n_171),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1179),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1132),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1166),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1138),
.A2(n_175),
.B1(n_177),
.B2(n_178),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1174),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1145),
.A2(n_183),
.B1(n_186),
.B2(n_188),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1162),
.B(n_1145),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1146),
.A2(n_191),
.B(n_193),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1185),
.B(n_195),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1190),
.B(n_196),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1157),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1198),
.B(n_1146),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1218),
.B(n_1143),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1200),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1199),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1242),
.B(n_1193),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1246),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1226),
.B(n_1143),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1228),
.B(n_1192),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1229),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1232),
.B(n_1237),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1221),
.A2(n_203),
.B(n_204),
.C(n_206),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1240),
.B(n_207),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1248),
.Y(n_1269)
);

INVx4_ASAP7_75t_SL g1270 ( 
.A(n_1254),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1199),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1199),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1238),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1206),
.B(n_218),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1239),
.B(n_224),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1201),
.B(n_231),
.Y(n_1276)
);

AND2x4_ASAP7_75t_SL g1277 ( 
.A(n_1254),
.B(n_234),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1247),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1214),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1197),
.B(n_235),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1214),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1222),
.B(n_238),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1195),
.A2(n_1203),
.B1(n_1196),
.B2(n_1251),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1214),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1223),
.B(n_243),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1202),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1255),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1254),
.B(n_245),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1252),
.Y(n_1289)
);

NAND2x1_ASAP7_75t_L g1290 ( 
.A(n_1204),
.B(n_247),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1227),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1210),
.B(n_249),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1253),
.B(n_252),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1207),
.B(n_255),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1208),
.B(n_259),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1211),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1209),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1219),
.B(n_262),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1230),
.B(n_267),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1230),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1213),
.B(n_268),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1243),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1241),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1225),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1216),
.Y(n_1305)
);

NOR2x1p5_ASAP7_75t_L g1306 ( 
.A(n_1215),
.B(n_270),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1220),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1258),
.B(n_1244),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1289),
.B(n_1244),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1269),
.B(n_1224),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1258),
.B(n_1249),
.Y(n_1311)
);

OAI221xp5_ASAP7_75t_L g1312 ( 
.A1(n_1303),
.A2(n_1234),
.B1(n_1236),
.B2(n_1256),
.C(n_1235),
.Y(n_1312)
);

AOI31xp33_ASAP7_75t_L g1313 ( 
.A1(n_1259),
.A2(n_1212),
.A3(n_1231),
.B(n_1205),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1262),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1265),
.Y(n_1315)
);

NAND2xp33_ASAP7_75t_R g1316 ( 
.A(n_1303),
.B(n_1217),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1260),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1278),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1283),
.A2(n_1250),
.B1(n_1233),
.B2(n_1245),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1260),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1307),
.A2(n_271),
.B1(n_272),
.B2(n_276),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1263),
.B(n_277),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_1273),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1279),
.B(n_278),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1257),
.B(n_280),
.Y(n_1325)
);

OR2x6_ASAP7_75t_SL g1326 ( 
.A(n_1259),
.B(n_281),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1278),
.Y(n_1327)
);

NOR4xp25_ASAP7_75t_SL g1328 ( 
.A(n_1297),
.B(n_285),
.C(n_287),
.D(n_288),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1271),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1257),
.B(n_294),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1279),
.B(n_300),
.Y(n_1331)
);

OAI21xp33_ASAP7_75t_L g1332 ( 
.A1(n_1301),
.A2(n_303),
.B(n_305),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1271),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1281),
.B(n_307),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1262),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_1273),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1286),
.Y(n_1337)
);

AOI221xp5_ASAP7_75t_L g1338 ( 
.A1(n_1295),
.A2(n_329),
.B1(n_311),
.B2(n_313),
.C(n_316),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1329),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1317),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1337),
.B(n_1284),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1335),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1314),
.B(n_1284),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1336),
.B(n_1281),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1333),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1323),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1323),
.B(n_1272),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1315),
.B(n_1296),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_1325),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1318),
.B(n_1305),
.Y(n_1350)
);

HB1xp67_ASAP7_75t_L g1351 ( 
.A(n_1327),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1317),
.B(n_1272),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1320),
.B(n_1270),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1320),
.B(n_1270),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1325),
.B(n_1270),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1310),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1324),
.Y(n_1357)
);

NAND2x1_ASAP7_75t_SL g1358 ( 
.A(n_1330),
.B(n_1297),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1308),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1351),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1340),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1356),
.B(n_1308),
.Y(n_1362)
);

INVxp67_ASAP7_75t_L g1363 ( 
.A(n_1348),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1359),
.B(n_1270),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1345),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1345),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1359),
.B(n_1326),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1346),
.B(n_1343),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1357),
.B(n_1296),
.Y(n_1369)
);

NOR2x1_ASAP7_75t_SL g1370 ( 
.A(n_1350),
.B(n_1355),
.Y(n_1370)
);

INVx4_ASAP7_75t_L g1371 ( 
.A(n_1346),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1343),
.B(n_1330),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1348),
.A2(n_1309),
.B(n_1313),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1357),
.B(n_1322),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1370),
.B(n_1355),
.Y(n_1375)
);

NAND2xp33_ASAP7_75t_R g1376 ( 
.A(n_1367),
.B(n_1328),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1364),
.B(n_1342),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1362),
.B(n_1342),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1365),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1373),
.B(n_1326),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1367),
.B(n_1349),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1363),
.B(n_1358),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1364),
.B(n_1344),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1369),
.B(n_1341),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1368),
.B(n_1372),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1368),
.B(n_1344),
.Y(n_1386)
);

OAI322xp33_ASAP7_75t_L g1387 ( 
.A1(n_1360),
.A2(n_1316),
.A3(n_1301),
.B1(n_1307),
.B2(n_1291),
.C1(n_1350),
.C2(n_1319),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1372),
.B(n_1358),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1371),
.B(n_1334),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1379),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1380),
.B(n_1374),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1384),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1377),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1375),
.B(n_1371),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1385),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1378),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1387),
.A2(n_1298),
.B1(n_1332),
.B2(n_1312),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1386),
.Y(n_1398)
);

AOI221xp5_ASAP7_75t_L g1399 ( 
.A1(n_1387),
.A2(n_1382),
.B1(n_1375),
.B2(n_1381),
.C(n_1388),
.Y(n_1399)
);

NOR2xp67_ASAP7_75t_L g1400 ( 
.A(n_1383),
.B(n_1371),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1390),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1395),
.B(n_1389),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1392),
.Y(n_1403)
);

AOI31xp33_ASAP7_75t_L g1404 ( 
.A1(n_1399),
.A2(n_1376),
.A3(n_1316),
.B(n_1261),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1394),
.Y(n_1405)
);

INVx8_ASAP7_75t_L g1406 ( 
.A(n_1400),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1396),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1391),
.A2(n_1277),
.B1(n_1298),
.B2(n_1294),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1393),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1398),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1398),
.Y(n_1411)
);

NAND2xp33_ASAP7_75t_L g1412 ( 
.A(n_1406),
.B(n_1397),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1406),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_R g1414 ( 
.A(n_1409),
.B(n_1397),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1411),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1405),
.B(n_1389),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1404),
.B(n_1366),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1411),
.B(n_1389),
.Y(n_1418)
);

XOR2xp5_ASAP7_75t_L g1419 ( 
.A(n_1408),
.B(n_1402),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1407),
.A2(n_1267),
.B(n_1338),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1415),
.B(n_1403),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_SL g1422 ( 
.A1(n_1413),
.A2(n_1411),
.B1(n_1401),
.B2(n_1410),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1412),
.A2(n_1401),
.B(n_1321),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1417),
.B(n_1341),
.Y(n_1424)
);

AOI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1414),
.A2(n_1266),
.B1(n_1293),
.B2(n_1321),
.C(n_1294),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_1418),
.B(n_1273),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1419),
.B(n_1361),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1417),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1416),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1420),
.B(n_1285),
.Y(n_1430)
);

AOI221xp5_ASAP7_75t_L g1431 ( 
.A1(n_1428),
.A2(n_1423),
.B1(n_1422),
.B2(n_1429),
.C(n_1430),
.Y(n_1431)
);

AOI322xp5_ASAP7_75t_L g1432 ( 
.A1(n_1425),
.A2(n_1311),
.A3(n_1293),
.B1(n_1288),
.B2(n_1292),
.C1(n_1304),
.C2(n_1290),
.Y(n_1432)
);

NAND2xp33_ASAP7_75t_SL g1433 ( 
.A(n_1427),
.B(n_1306),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1421),
.Y(n_1434)
);

NAND2xp33_ASAP7_75t_R g1435 ( 
.A(n_1424),
.B(n_1288),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1426),
.A2(n_1290),
.B(n_1285),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1423),
.A2(n_1277),
.B(n_1282),
.Y(n_1437)
);

OAI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1423),
.A2(n_1287),
.B1(n_1280),
.B2(n_1276),
.C(n_1304),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1434),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1433),
.A2(n_1334),
.B1(n_1331),
.B2(n_1353),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1435),
.Y(n_1441)
);

NAND2xp33_ASAP7_75t_R g1442 ( 
.A(n_1437),
.B(n_1334),
.Y(n_1442)
);

NOR3xp33_ASAP7_75t_L g1443 ( 
.A(n_1431),
.B(n_1275),
.C(n_1299),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1438),
.Y(n_1444)
);

A2O1A1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1443),
.A2(n_1432),
.B(n_1436),
.C(n_1280),
.Y(n_1445)
);

INVx3_ASAP7_75t_SL g1446 ( 
.A(n_1439),
.Y(n_1446)
);

NAND3xp33_ASAP7_75t_L g1447 ( 
.A(n_1441),
.B(n_1268),
.C(n_1276),
.Y(n_1447)
);

FAx1_ASAP7_75t_SL g1448 ( 
.A(n_1440),
.B(n_1354),
.CI(n_1353),
.CON(n_1448),
.SN(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1444),
.A2(n_1331),
.B(n_1299),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1442),
.A2(n_1292),
.B1(n_1331),
.B2(n_1311),
.C(n_1274),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1439),
.B(n_1361),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1451),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1446),
.B(n_1273),
.Y(n_1453)
);

NAND4xp25_ASAP7_75t_L g1454 ( 
.A(n_1445),
.B(n_1449),
.C(n_1447),
.D(n_1448),
.Y(n_1454)
);

NAND3xp33_ASAP7_75t_SL g1455 ( 
.A(n_1450),
.B(n_1268),
.C(n_1274),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1451),
.B(n_1354),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1452),
.A2(n_1273),
.B1(n_1347),
.B2(n_1339),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1453),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1456),
.Y(n_1459)
);

BUFx8_ASAP7_75t_SL g1460 ( 
.A(n_1454),
.Y(n_1460)
);

NOR2x1_ASAP7_75t_L g1461 ( 
.A(n_1459),
.B(n_1455),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1460),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1461),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1462),
.A2(n_1458),
.B1(n_1457),
.B2(n_1347),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1463),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1464),
.Y(n_1466)
);

OAI21xp33_ASAP7_75t_L g1467 ( 
.A1(n_1466),
.A2(n_1347),
.B(n_1339),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1467),
.A2(n_1465),
.B1(n_1302),
.B2(n_1339),
.Y(n_1468)
);

AOI322xp5_ASAP7_75t_L g1469 ( 
.A1(n_1468),
.A2(n_1347),
.A3(n_1302),
.B1(n_1352),
.B2(n_1340),
.C1(n_1264),
.C2(n_1300),
.Y(n_1469)
);

OAI221xp5_ASAP7_75t_R g1470 ( 
.A1(n_1469),
.A2(n_310),
.B1(n_320),
.B2(n_321),
.C(n_322),
.Y(n_1470)
);

AOI211xp5_ASAP7_75t_L g1471 ( 
.A1(n_1470),
.A2(n_323),
.B(n_1264),
.C(n_1352),
.Y(n_1471)
);


endmodule