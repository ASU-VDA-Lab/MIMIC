module fake_ariane_120_n_1982 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_172, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1982);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1982;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_699;
wire n_590;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_181;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_177;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_SL g173 ( 
.A(n_45),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_11),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_104),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_83),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_103),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_33),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_63),
.Y(n_179)
);

BUFx2_ASAP7_75t_SL g180 ( 
.A(n_24),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_76),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_16),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_95),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_129),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_106),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_45),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_86),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_32),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_112),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_101),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_65),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_25),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_158),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_167),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_115),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_108),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_146),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_90),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_34),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_118),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_53),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_134),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_78),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_114),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_81),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_75),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_80),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_32),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_14),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_73),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_138),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_60),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_28),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_99),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_36),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_44),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_137),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_126),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_87),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_27),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_23),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_142),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_135),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_168),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_155),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_152),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_1),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_144),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_109),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_166),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_21),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_161),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_122),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_162),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_33),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_125),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_107),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_54),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_12),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_92),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_39),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_6),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_11),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_111),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_21),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_25),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_66),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_116),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_98),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_127),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_51),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_100),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_110),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_105),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_139),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_31),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_63),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_10),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_71),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_2),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_121),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_68),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_49),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_36),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_131),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_72),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_13),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_79),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_18),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_117),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_58),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_88),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_102),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_65),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_60),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_67),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_140),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_8),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_47),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_61),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_93),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_149),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_12),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_18),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_28),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_26),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_44),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_51),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_6),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_5),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_3),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_91),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_57),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_15),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_123),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_54),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_74),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_67),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_71),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_30),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_52),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_119),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_13),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_97),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_50),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_53),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_136),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_141),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_153),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_48),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_94),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_159),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_35),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_46),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_96),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_150),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_128),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_156),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_14),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_43),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_89),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_23),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_59),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_113),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_16),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_151),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_124),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_7),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_157),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_10),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_20),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_40),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_20),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_1),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_169),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_41),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_15),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_160),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_37),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_205),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_174),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_240),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_174),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_175),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_174),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_185),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_279),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_174),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_300),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_205),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_174),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_R g357 ( 
.A(n_187),
.B(n_172),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_215),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_174),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_174),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_L g361 ( 
.A(n_173),
.B(n_0),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_307),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_174),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_174),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_309),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_181),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_314),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_181),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_329),
.Y(n_369)
);

NOR2xp67_ASAP7_75t_L g370 ( 
.A(n_173),
.B(n_0),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_205),
.B(n_2),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_191),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_179),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_182),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_191),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_188),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_199),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_304),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_190),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_263),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_296),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_286),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_199),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_286),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_238),
.B(n_3),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_195),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_196),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_204),
.B(n_4),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_204),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_207),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_207),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_209),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_209),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_210),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_193),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_193),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_203),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_193),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_210),
.B(n_4),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_226),
.B(n_5),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_226),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_217),
.B(n_7),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_234),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_234),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_237),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_237),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_212),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_239),
.B(n_8),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_304),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_239),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_236),
.B(n_9),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_236),
.B(n_9),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_323),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_323),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_213),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_216),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_323),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_259),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_259),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_219),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_260),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_260),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_217),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_217),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_304),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_225),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_266),
.B(n_17),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_217),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_266),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_232),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_409),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_378),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_346),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_349),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_380),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_351),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_362),
.Y(n_438)
);

OA21x2_ASAP7_75t_L g439 ( 
.A1(n_378),
.A2(n_313),
.B(n_273),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_425),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g441 ( 
.A(n_365),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_367),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_366),
.B(n_224),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_366),
.B(n_273),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_382),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_358),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_348),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_355),
.B(n_224),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_348),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_350),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_369),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_350),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_353),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_373),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_416),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_353),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_374),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_356),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_384),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_385),
.B(n_313),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_356),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_359),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_359),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_381),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_360),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_430),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_360),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_363),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_363),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_364),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_368),
.B(n_304),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_364),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_347),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_376),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_368),
.Y(n_476)
);

NAND3xp33_ASAP7_75t_L g477 ( 
.A(n_388),
.B(n_408),
.C(n_371),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_372),
.B(n_331),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_372),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_402),
.A2(n_285),
.B1(n_295),
.B2(n_305),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_375),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_375),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_379),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_377),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_R g485 ( 
.A(n_354),
.B(n_177),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_386),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_371),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_377),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_387),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_355),
.B(n_178),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_383),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_397),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_383),
.B(n_389),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_389),
.B(n_331),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_407),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_415),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_390),
.B(n_201),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_426),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_402),
.B(n_201),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_395),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_390),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_391),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_391),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_392),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_396),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_392),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_423),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_451),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_479),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_487),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_487),
.B(n_398),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_479),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_451),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_481),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_487),
.B(n_413),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_345),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_431),
.B(n_414),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_469),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_481),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_469),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_482),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_454),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_441),
.B(n_352),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_R g524 ( 
.A(n_435),
.B(n_357),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_431),
.B(n_417),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_482),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_437),
.Y(n_527)
);

INVx8_ASAP7_75t_L g528 ( 
.A(n_493),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_493),
.B(n_411),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_484),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_461),
.B(n_393),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_477),
.B(n_461),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_493),
.B(n_393),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_493),
.B(n_176),
.Y(n_534)
);

OR2x6_ASAP7_75t_L g535 ( 
.A(n_467),
.B(n_486),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_477),
.B(n_420),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_493),
.B(n_394),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_448),
.B(n_411),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_500),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_454),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_438),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_454),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_469),
.B(n_176),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_451),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_484),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_442),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_451),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_456),
.B(n_394),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_505),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_467),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_R g551 ( 
.A(n_455),
.B(n_424),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_488),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_501),
.B(n_401),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_468),
.B(n_176),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_462),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_488),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_502),
.Y(n_557)
);

OR2x6_ASAP7_75t_L g558 ( 
.A(n_486),
.B(n_412),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_501),
.B(n_401),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_446),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_456),
.A2(n_412),
.B1(n_370),
.B2(n_361),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_462),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_499),
.B(n_502),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_501),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_501),
.B(n_403),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_503),
.B(n_403),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_468),
.B(n_227),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_468),
.B(n_462),
.Y(n_568)
);

AND2x6_ASAP7_75t_L g569 ( 
.A(n_472),
.B(n_227),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_503),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_441),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_451),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_506),
.B(n_458),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_506),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_448),
.B(n_404),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_468),
.B(n_404),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_476),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_433),
.B(n_405),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_473),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_433),
.B(n_405),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_476),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_473),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_443),
.B(n_406),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_475),
.B(n_406),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_476),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_491),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_490),
.A2(n_399),
.B1(n_427),
.B2(n_400),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_451),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_443),
.B(n_410),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_451),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_491),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_473),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_490),
.A2(n_248),
.B1(n_243),
.B2(n_244),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_491),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_504),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_480),
.A2(n_429),
.B1(n_410),
.B2(n_422),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_434),
.B(n_418),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_434),
.B(n_418),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_453),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_453),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_448),
.B(n_419),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_504),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_447),
.B(n_227),
.Y(n_603)
);

INVx4_ASAP7_75t_L g604 ( 
.A(n_453),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_432),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_447),
.B(n_233),
.Y(n_606)
);

AND2x2_ASAP7_75t_SL g607 ( 
.A(n_492),
.B(n_233),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_490),
.B(n_419),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_436),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_504),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_453),
.Y(n_611)
);

NAND2x1p5_ASAP7_75t_L g612 ( 
.A(n_443),
.B(n_421),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_432),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_443),
.B(n_444),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_452),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_453),
.Y(n_616)
);

OR2x6_ASAP7_75t_L g617 ( 
.A(n_492),
.B(n_180),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_453),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_453),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_432),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_443),
.B(n_421),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_449),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_449),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_470),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_449),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_445),
.B(n_422),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_483),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_489),
.B(n_429),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_450),
.B(n_198),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_444),
.B(n_178),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_472),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_470),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_450),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_478),
.B(n_220),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_470),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_470),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_478),
.B(n_220),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_495),
.B(n_428),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_457),
.B(n_233),
.Y(n_639)
);

INVx4_ASAP7_75t_SL g640 ( 
.A(n_470),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_470),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_465),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_472),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_457),
.B(n_257),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_472),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_472),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_480),
.A2(n_310),
.B1(n_272),
.B2(n_283),
.Y(n_647)
);

AND2x6_ASAP7_75t_L g648 ( 
.A(n_459),
.B(n_257),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_497),
.B(n_272),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_496),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_445),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_459),
.B(n_317),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_470),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_471),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_471),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_471),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_463),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_471),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_460),
.Y(n_659)
);

AND2x6_ASAP7_75t_L g660 ( 
.A(n_463),
.B(n_257),
.Y(n_660)
);

BUFx12f_ASAP7_75t_SL g661 ( 
.A(n_535),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_532),
.B(n_498),
.C(n_460),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_523),
.B(n_474),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_584),
.B(n_497),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_628),
.B(n_464),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_577),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_522),
.Y(n_667)
);

NOR2x2_ASAP7_75t_L g668 ( 
.A(n_535),
.B(n_507),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_531),
.B(n_464),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_548),
.B(n_466),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_607),
.B(n_494),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_510),
.B(n_466),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_650),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_510),
.B(n_494),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_614),
.B(n_485),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_607),
.B(n_439),
.Y(n_676)
);

BUFx8_ASAP7_75t_L g677 ( 
.A(n_627),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_650),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_522),
.Y(n_679)
);

NAND2x1p5_ASAP7_75t_L g680 ( 
.A(n_564),
.B(n_518),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_614),
.B(n_485),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_608),
.B(n_439),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_536),
.A2(n_573),
.B1(n_529),
.B2(n_587),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_528),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_540),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_581),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_516),
.B(n_471),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_630),
.B(n_471),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_585),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_523),
.B(n_246),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_511),
.B(n_247),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_528),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_515),
.B(n_250),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_586),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_630),
.B(n_471),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_647),
.A2(n_439),
.B1(n_180),
.B2(n_304),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_563),
.A2(n_283),
.B(n_284),
.C(n_291),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_540),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_634),
.B(n_439),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_634),
.B(n_637),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_538),
.A2(n_439),
.B1(n_304),
.B2(n_339),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_568),
.A2(n_249),
.B(n_229),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_538),
.A2(n_339),
.B1(n_229),
.B2(n_249),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_637),
.B(n_284),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_608),
.B(n_251),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_591),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_542),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_571),
.Y(n_708)
);

AND2x2_ASAP7_75t_SL g709 ( 
.A(n_596),
.B(n_297),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_649),
.B(n_291),
.Y(n_710)
);

NOR2x1p5_ASAP7_75t_L g711 ( 
.A(n_527),
.B(n_252),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_528),
.A2(n_276),
.B1(n_344),
.B2(n_274),
.Y(n_712)
);

NOR3xp33_ASAP7_75t_L g713 ( 
.A(n_550),
.B(n_310),
.C(n_294),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_608),
.B(n_256),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_651),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_528),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_542),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_649),
.B(n_294),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_575),
.B(n_311),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_626),
.Y(n_720)
);

BUFx6f_ASAP7_75t_SL g721 ( 
.A(n_535),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_649),
.B(n_311),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_555),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_538),
.A2(n_339),
.B1(n_297),
.B2(n_322),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_626),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_575),
.B(n_315),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_518),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_575),
.B(n_315),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_601),
.B(n_325),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_601),
.B(n_325),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_648),
.B(n_660),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_555),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_517),
.B(n_525),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_529),
.A2(n_339),
.B1(n_322),
.B2(n_326),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_513),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_562),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_659),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_558),
.B(n_261),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_SL g739 ( 
.A1(n_657),
.A2(n_327),
.B(n_328),
.C(n_326),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_513),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_558),
.B(n_262),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_564),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_529),
.B(n_264),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_601),
.B(n_327),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_562),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_583),
.B(n_328),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_564),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_612),
.B(n_265),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_569),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_612),
.B(n_267),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_568),
.A2(n_641),
.B(n_636),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_627),
.B(n_268),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_636),
.A2(n_440),
.B(n_340),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_629),
.B(n_269),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_569),
.A2(n_214),
.B1(n_343),
.B2(n_228),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_569),
.A2(n_208),
.B1(n_222),
.B2(n_221),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_652),
.B(n_280),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_569),
.A2(n_339),
.B1(n_297),
.B2(n_326),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_583),
.B(n_281),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_579),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_594),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_595),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_569),
.A2(n_561),
.B1(n_621),
.B2(n_589),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_569),
.A2(n_339),
.B1(n_322),
.B2(n_340),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_589),
.B(n_288),
.Y(n_765)
);

NOR2x1p5_ASAP7_75t_L g766 ( 
.A(n_527),
.B(n_289),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_621),
.B(n_617),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_534),
.A2(n_194),
.B1(n_189),
.B2(n_197),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_533),
.B(n_537),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_558),
.B(n_290),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_L g771 ( 
.A(n_541),
.B(n_183),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_558),
.B(n_292),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_509),
.B(n_293),
.Y(n_773)
);

BUFx2_ASAP7_75t_SL g774 ( 
.A(n_648),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_579),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_535),
.Y(n_776)
);

NOR2x2_ASAP7_75t_L g777 ( 
.A(n_617),
.B(n_340),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_512),
.B(n_298),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_534),
.A2(n_330),
.B1(n_342),
.B2(n_341),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_602),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_560),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_610),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_541),
.B(n_299),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_514),
.B(n_519),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_631),
.B(n_301),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_521),
.B(n_526),
.Y(n_786)
);

INVx8_ASAP7_75t_L g787 ( 
.A(n_648),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_520),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_530),
.B(n_303),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_582),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_593),
.B(n_306),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_545),
.B(n_308),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_SL g793 ( 
.A1(n_552),
.A2(n_338),
.B(n_318),
.C(n_319),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_520),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_556),
.B(n_324),
.Y(n_795)
);

OR2x6_ASAP7_75t_L g796 ( 
.A(n_617),
.B(n_440),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_582),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_617),
.B(n_333),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_638),
.B(n_335),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_546),
.B(n_539),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_557),
.B(n_336),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_633),
.A2(n_255),
.B1(n_206),
.B2(n_192),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_592),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_570),
.B(n_337),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_633),
.A2(n_440),
.B1(n_334),
.B2(n_186),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_609),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_592),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_551),
.B(n_200),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_549),
.B(n_202),
.Y(n_809)
);

NAND2x1p5_ASAP7_75t_L g810 ( 
.A(n_599),
.B(n_600),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_574),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_605),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_643),
.B(n_211),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_645),
.B(n_223),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_646),
.B(n_440),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_553),
.B(n_230),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_566),
.B(n_231),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_605),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_613),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_613),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_576),
.A2(n_275),
.B(n_235),
.C(n_332),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_599),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_642),
.B(n_241),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_559),
.B(n_242),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_565),
.B(n_245),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_578),
.B(n_253),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_580),
.B(n_597),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_620),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_560),
.B(n_254),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_615),
.B(n_258),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_648),
.A2(n_440),
.B1(n_334),
.B2(n_186),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_598),
.B(n_270),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_811),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_684),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_664),
.B(n_733),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_671),
.B(n_648),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_684),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_684),
.Y(n_838)
);

INVx4_ASAP7_75t_L g839 ( 
.A(n_684),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_811),
.Y(n_840)
);

INVx4_ASAP7_75t_L g841 ( 
.A(n_684),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_673),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_819),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_673),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_671),
.B(n_648),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_715),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_666),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_665),
.B(n_700),
.Y(n_848)
);

NOR3xp33_ASAP7_75t_SL g849 ( 
.A(n_678),
.B(n_615),
.C(n_524),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_819),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_767),
.B(n_640),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_827),
.B(n_660),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_827),
.B(n_660),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_767),
.B(n_640),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_749),
.Y(n_855)
);

INVx5_ASAP7_75t_L g856 ( 
.A(n_749),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_666),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_683),
.B(n_660),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_677),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_691),
.B(n_660),
.Y(n_860)
);

INVx3_ASAP7_75t_SL g861 ( 
.A(n_678),
.Y(n_861)
);

INVx4_ASAP7_75t_L g862 ( 
.A(n_749),
.Y(n_862)
);

NOR3xp33_ASAP7_75t_SL g863 ( 
.A(n_783),
.B(n_567),
.C(n_554),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_675),
.B(n_599),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_670),
.B(n_660),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_681),
.B(n_600),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_735),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_686),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_677),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_677),
.Y(n_870)
);

NAND2x1p5_ASAP7_75t_L g871 ( 
.A(n_692),
.B(n_600),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_690),
.B(n_604),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_720),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_720),
.B(n_543),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_799),
.B(n_604),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_806),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_R g877 ( 
.A(n_708),
.B(n_513),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_667),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_767),
.A2(n_567),
.B1(n_554),
.B2(n_543),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_686),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_689),
.Y(n_881)
);

OR2x6_ASAP7_75t_L g882 ( 
.A(n_796),
.B(n_603),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_667),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_788),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_692),
.B(n_640),
.Y(n_885)
);

BUFx4f_ASAP7_75t_L g886 ( 
.A(n_781),
.Y(n_886)
);

NOR3xp33_ASAP7_75t_SL g887 ( 
.A(n_752),
.B(n_321),
.C(n_320),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_679),
.Y(n_888)
);

INVx5_ASAP7_75t_L g889 ( 
.A(n_787),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_725),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_689),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_694),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_694),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_679),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_788),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_725),
.B(n_603),
.Y(n_896)
);

CKINVDCx16_ASAP7_75t_R g897 ( 
.A(n_708),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_669),
.B(n_604),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_794),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_663),
.B(n_606),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_706),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_693),
.B(n_616),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_706),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_794),
.Y(n_904)
);

BUFx4f_ASAP7_75t_L g905 ( 
.A(n_781),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_761),
.Y(n_906)
);

NOR3xp33_ASAP7_75t_SL g907 ( 
.A(n_705),
.B(n_316),
.C(n_312),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_761),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_762),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_776),
.B(n_616),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_762),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_780),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_800),
.B(n_606),
.C(n_644),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_SL g914 ( 
.A(n_714),
.B(n_302),
.C(n_287),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_780),
.Y(n_915)
);

AND2x6_ASAP7_75t_L g916 ( 
.A(n_676),
.B(n_641),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_754),
.B(n_757),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_782),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_782),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_742),
.B(n_508),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_735),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_784),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_709),
.B(n_769),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_786),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_661),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_716),
.B(n_640),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_815),
.Y(n_927)
);

NOR3xp33_ASAP7_75t_SL g928 ( 
.A(n_829),
.B(n_282),
.C(n_278),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_815),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_709),
.B(n_616),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_742),
.B(n_508),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_742),
.B(n_508),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_735),
.Y(n_933)
);

OR2x6_ASAP7_75t_L g934 ( 
.A(n_796),
.B(n_639),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_716),
.B(n_618),
.Y(n_935)
);

BUFx4f_ASAP7_75t_L g936 ( 
.A(n_796),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_763),
.B(n_618),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_747),
.B(n_682),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_685),
.Y(n_939)
);

INVx2_ASAP7_75t_SL g940 ( 
.A(n_711),
.Y(n_940)
);

INVx5_ASAP7_75t_L g941 ( 
.A(n_787),
.Y(n_941)
);

INVxp67_ASAP7_75t_L g942 ( 
.A(n_737),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_735),
.Y(n_943)
);

INVx4_ASAP7_75t_L g944 ( 
.A(n_787),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_823),
.Y(n_945)
);

BUFx10_ASAP7_75t_L g946 ( 
.A(n_830),
.Y(n_946)
);

CKINVDCx11_ASAP7_75t_R g947 ( 
.A(n_796),
.Y(n_947)
);

NAND2x1p5_ASAP7_75t_L g948 ( 
.A(n_727),
.B(n_618),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_682),
.B(n_619),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_674),
.B(n_619),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_735),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_728),
.B(n_639),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_790),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_746),
.B(n_619),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_685),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_748),
.B(n_635),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_746),
.B(n_635),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_766),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_704),
.B(n_635),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_719),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_790),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_740),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_719),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_807),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_785),
.B(n_644),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_698),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_807),
.Y(n_967)
);

OR2x4_ASAP7_75t_L g968 ( 
.A(n_809),
.B(n_508),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_726),
.B(n_653),
.Y(n_969)
);

INVx5_ASAP7_75t_L g970 ( 
.A(n_787),
.Y(n_970)
);

NOR3xp33_ASAP7_75t_SL g971 ( 
.A(n_712),
.B(n_271),
.C(n_277),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_750),
.B(n_653),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_661),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_785),
.B(n_620),
.Y(n_974)
);

INVx8_ASAP7_75t_L g975 ( 
.A(n_721),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_688),
.B(n_622),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_726),
.B(n_622),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_759),
.B(n_655),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_740),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_812),
.Y(n_980)
);

NOR3xp33_ASAP7_75t_SL g981 ( 
.A(n_821),
.B(n_17),
.C(n_19),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_695),
.B(n_623),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_740),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_SL g984 ( 
.A(n_743),
.B(n_19),
.C(n_22),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_710),
.B(n_623),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_729),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_740),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_740),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_R g989 ( 
.A(n_721),
.B(n_513),
.Y(n_989)
);

NAND2x1p5_ASAP7_75t_L g990 ( 
.A(n_727),
.B(n_544),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_698),
.Y(n_991)
);

NAND2x1p5_ASAP7_75t_L g992 ( 
.A(n_676),
.B(n_544),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_680),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_707),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_680),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_810),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_680),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_812),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_747),
.B(n_508),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_721),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_810),
.Y(n_1001)
);

CKINVDCx8_ASAP7_75t_R g1002 ( 
.A(n_798),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_707),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_818),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_818),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_820),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_822),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_668),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_717),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_717),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_820),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_765),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_672),
.A2(n_658),
.B(n_655),
.Y(n_1013)
);

AND2x2_ASAP7_75t_SL g1014 ( 
.A(n_731),
.B(n_184),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_828),
.Y(n_1015)
);

NOR3xp33_ASAP7_75t_SL g1016 ( 
.A(n_817),
.B(n_22),
.C(n_24),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_810),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_L g1018 ( 
.A(n_668),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_718),
.B(n_625),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_747),
.B(n_654),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_828),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_662),
.A2(n_738),
.B1(n_741),
.B2(n_772),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_722),
.B(n_625),
.Y(n_1023)
);

OR2x6_ASAP7_75t_L g1024 ( 
.A(n_774),
.B(n_658),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_723),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_875),
.A2(n_835),
.B(n_848),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_1013),
.A2(n_751),
.B(n_753),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_872),
.A2(n_731),
.B(n_687),
.Y(n_1028)
);

NOR3xp33_ASAP7_75t_L g1029 ( 
.A(n_945),
.B(n_1012),
.C(n_917),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_833),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_922),
.B(n_770),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_851),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_924),
.B(n_730),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_851),
.B(n_822),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_860),
.A2(n_898),
.B(n_865),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_897),
.Y(n_1036)
);

AOI21xp33_ASAP7_75t_L g1037 ( 
.A1(n_900),
.A2(n_791),
.B(n_699),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_978),
.A2(n_702),
.B(n_822),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_917),
.A2(n_697),
.B(n_713),
.C(n_778),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_992),
.A2(n_732),
.B(n_797),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_1014),
.B(n_654),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_960),
.B(n_963),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_986),
.B(n_744),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_978),
.A2(n_824),
.B(n_816),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_923),
.A2(n_703),
.B1(n_696),
.B2(n_724),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_843),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1014),
.A2(n_832),
.B1(n_826),
.B2(n_825),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_873),
.B(n_890),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_840),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_938),
.A2(n_755),
.B(n_756),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_886),
.B(n_771),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_937),
.B(n_654),
.Y(n_1052)
);

AO31x2_ASAP7_75t_L g1053 ( 
.A1(n_972),
.A2(n_760),
.A3(n_745),
.B(n_732),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_847),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_873),
.B(n_890),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_992),
.A2(n_736),
.B(n_797),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_938),
.A2(n_813),
.B(n_814),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_846),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_1002),
.B(n_773),
.Y(n_1059)
);

NOR2xp67_ASAP7_75t_L g1060 ( 
.A(n_876),
.B(n_808),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_976),
.A2(n_745),
.B(n_736),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_977),
.B(n_789),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1022),
.B(n_792),
.Y(n_1063)
);

AOI211x1_ASAP7_75t_L g1064 ( 
.A1(n_857),
.A2(n_795),
.B(n_801),
.C(n_804),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_846),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_851),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_843),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_842),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_950),
.A2(n_723),
.B(n_803),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_982),
.A2(n_931),
.B(n_920),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_864),
.A2(n_803),
.B(n_760),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_937),
.A2(n_775),
.B(n_779),
.C(n_764),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_864),
.A2(n_775),
.B(n_654),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_954),
.A2(n_701),
.B(n_802),
.Y(n_1074)
);

INVx5_ASAP7_75t_L g1075 ( 
.A(n_916),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_996),
.B(n_654),
.Y(n_1076)
);

INVxp67_ASAP7_75t_SL g1077 ( 
.A(n_936),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_854),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_L g1079 ( 
.A(n_844),
.B(n_768),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_868),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_896),
.B(n_734),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_969),
.B(n_758),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_957),
.A2(n_866),
.B(n_959),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_969),
.B(n_774),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_866),
.A2(n_853),
.B(n_852),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_877),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_969),
.B(n_544),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_880),
.B(n_881),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_891),
.A2(n_831),
.B1(n_656),
.B2(n_588),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_942),
.B(n_777),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_892),
.A2(n_656),
.B1(n_544),
.B2(n_572),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_SL g1092 ( 
.A1(n_858),
.A2(n_805),
.B(n_739),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_920),
.A2(n_656),
.B(n_547),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_931),
.A2(n_793),
.B(n_656),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_893),
.B(n_901),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_932),
.A2(n_656),
.B(n_590),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_903),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_SL g1098 ( 
.A1(n_862),
.A2(n_572),
.B(n_632),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_SL g1099 ( 
.A1(n_965),
.A2(n_908),
.B(n_906),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_909),
.B(n_590),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_877),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_1016),
.A2(n_777),
.B(n_632),
.C(n_624),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_911),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_932),
.A2(n_632),
.B(n_624),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_912),
.B(n_632),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_999),
.A2(n_624),
.B(n_611),
.Y(n_1106)
);

NOR2xp67_ASAP7_75t_SL g1107 ( 
.A(n_859),
.B(n_624),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_999),
.A2(n_611),
.B(n_590),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1020),
.A2(n_611),
.B(n_590),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1020),
.A2(n_611),
.B(n_588),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_993),
.A2(n_588),
.B(n_572),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_993),
.A2(n_588),
.B(n_572),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_886),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_915),
.B(n_547),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_956),
.A2(n_547),
.B(n_334),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_918),
.B(n_547),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_905),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_956),
.A2(n_334),
.B(n_218),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_995),
.A2(n_440),
.B(n_334),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_850),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_919),
.B(n_26),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_995),
.A2(n_440),
.B(n_334),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_930),
.A2(n_27),
.B(n_29),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_856),
.A2(n_218),
.B(n_186),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_854),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_927),
.B(n_29),
.Y(n_1126)
);

O2A1O1Ixp5_ASAP7_75t_L g1127 ( 
.A1(n_902),
.A2(n_30),
.B(n_31),
.C(n_34),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_929),
.B(n_35),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_SL g1129 ( 
.A1(n_862),
.A2(n_1007),
.B(n_845),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_953),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_854),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_946),
.B(n_37),
.Y(n_1132)
);

O2A1O1Ixp5_ASAP7_75t_L g1133 ( 
.A1(n_902),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_856),
.A2(n_218),
.B(n_186),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_948),
.A2(n_218),
.B(n_186),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_948),
.A2(n_218),
.B(n_186),
.Y(n_1136)
);

OAI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_972),
.A2(n_949),
.B(n_974),
.Y(n_1137)
);

AO22x2_ASAP7_75t_L g1138 ( 
.A1(n_913),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_850),
.A2(n_991),
.A3(n_878),
.B(n_939),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_874),
.B(n_42),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_946),
.B(n_43),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_990),
.A2(n_218),
.B(n_184),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_990),
.A2(n_184),
.B(n_171),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_884),
.B(n_895),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_878),
.A2(n_184),
.B(n_170),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_961),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_884),
.B(n_46),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_867),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_905),
.B(n_47),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_856),
.A2(n_184),
.B(n_165),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_895),
.B(n_48),
.Y(n_1151)
);

INVx4_ASAP7_75t_L g1152 ( 
.A(n_889),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_910),
.B(n_49),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1016),
.A2(n_184),
.B(n_52),
.C(n_55),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_981),
.A2(n_50),
.B(n_55),
.C(n_56),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_910),
.B(n_56),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_883),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_836),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_1158)
);

NAND2xp33_ASAP7_75t_SL g1159 ( 
.A(n_944),
.B(n_61),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_949),
.A2(n_62),
.B(n_64),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_883),
.A2(n_84),
.B(n_145),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_856),
.A2(n_82),
.B(n_143),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_996),
.B(n_62),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_964),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_952),
.B(n_967),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_980),
.B(n_64),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_975),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1007),
.A2(n_85),
.B(n_133),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_998),
.B(n_66),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_996),
.B(n_68),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1004),
.B(n_69),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_981),
.A2(n_69),
.B(n_70),
.C(n_77),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_949),
.A2(n_70),
.B(n_130),
.Y(n_1173)
);

INVxp67_ASAP7_75t_L g1174 ( 
.A(n_925),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_935),
.A2(n_132),
.B(n_154),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1005),
.A2(n_1011),
.B(n_1006),
.Y(n_1176)
);

NOR2xp67_ASAP7_75t_SL g1177 ( 
.A(n_859),
.B(n_869),
.Y(n_1177)
);

AO31x2_ASAP7_75t_L g1178 ( 
.A1(n_888),
.A2(n_894),
.A3(n_966),
.B(n_991),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_935),
.A2(n_855),
.B(n_1023),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_935),
.A2(n_855),
.B(n_985),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1015),
.A2(n_1021),
.B(n_879),
.Y(n_1181)
);

AO22x2_ASAP7_75t_L g1182 ( 
.A1(n_1025),
.A2(n_1003),
.B1(n_1009),
.B2(n_994),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_899),
.B(n_904),
.Y(n_1183)
);

AO21x2_ASAP7_75t_L g1184 ( 
.A1(n_1019),
.A2(n_863),
.B(n_966),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_996),
.B(n_867),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1024),
.A2(n_979),
.B(n_921),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_899),
.B(n_904),
.Y(n_1187)
);

AOI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1024),
.A2(n_1003),
.B(n_939),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1029),
.A2(n_1018),
.B1(n_1008),
.B2(n_1031),
.Y(n_1189)
);

AOI22x1_ASAP7_75t_L g1190 ( 
.A1(n_1026),
.A2(n_871),
.B1(n_921),
.B2(n_933),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1027),
.A2(n_1061),
.B(n_1119),
.Y(n_1191)
);

OR2x6_ASAP7_75t_L g1192 ( 
.A(n_1101),
.B(n_975),
.Y(n_1192)
);

NOR2x1_ASAP7_75t_SL g1193 ( 
.A(n_1075),
.B(n_1024),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_SL g1194 ( 
.A1(n_1099),
.A2(n_841),
.B(n_839),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_SL g1195 ( 
.A1(n_1149),
.A2(n_1018),
.B1(n_975),
.B2(n_869),
.Y(n_1195)
);

INVxp67_ASAP7_75t_SL g1196 ( 
.A(n_1048),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1027),
.A2(n_1010),
.B(n_894),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_SL g1198 ( 
.A1(n_1063),
.A2(n_834),
.B(n_838),
.C(n_940),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1075),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1039),
.A2(n_1047),
.B(n_1173),
.C(n_1123),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1030),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1139),
.Y(n_1202)
);

NOR2x1_ASAP7_75t_L g1203 ( 
.A(n_1144),
.B(n_870),
.Y(n_1203)
);

CKINVDCx11_ASAP7_75t_R g1204 ( 
.A(n_1036),
.Y(n_1204)
);

BUFx12f_ASAP7_75t_L g1205 ( 
.A(n_1068),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_SL g1206 ( 
.A1(n_1149),
.A2(n_870),
.B1(n_989),
.B2(n_936),
.Y(n_1206)
);

INVx6_ASAP7_75t_L g1207 ( 
.A(n_1066),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1028),
.A2(n_943),
.B(n_921),
.Y(n_1208)
);

AO21x2_ASAP7_75t_L g1209 ( 
.A1(n_1035),
.A2(n_863),
.B(n_1010),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1139),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1167),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_1036),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1061),
.A2(n_994),
.B(n_1009),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1075),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1119),
.A2(n_888),
.B(n_955),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_SL g1216 ( 
.A1(n_1129),
.A2(n_841),
.B(n_839),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1032),
.B(n_934),
.Y(n_1217)
);

OAI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1090),
.A2(n_861),
.B1(n_968),
.B2(n_882),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1122),
.A2(n_955),
.B(n_871),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1058),
.A2(n_1062),
.B1(n_1138),
.B2(n_1160),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1059),
.B(n_861),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1139),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1049),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1032),
.B(n_1017),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1059),
.B(n_973),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_1071),
.A2(n_968),
.A3(n_944),
.B(n_916),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1181),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_1072),
.A2(n_916),
.A3(n_934),
.B(n_882),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1083),
.A2(n_928),
.B(n_914),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1153),
.A2(n_971),
.B1(n_849),
.B2(n_984),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1139),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1054),
.Y(n_1232)
);

NAND2xp33_ASAP7_75t_SL g1233 ( 
.A(n_1088),
.B(n_989),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1080),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1075),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1138),
.A2(n_947),
.B1(n_916),
.B2(n_934),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1178),
.Y(n_1237)
);

AOI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1052),
.A2(n_1115),
.B(n_1118),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1097),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1065),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1167),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1066),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1178),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1066),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1103),
.Y(n_1245)
);

NAND3xp33_ASAP7_75t_L g1246 ( 
.A(n_1154),
.B(n_984),
.C(n_971),
.Y(n_1246)
);

AOI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1052),
.A2(n_882),
.B(n_885),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1072),
.A2(n_916),
.A3(n_997),
.B(n_1001),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1122),
.A2(n_834),
.B(n_838),
.Y(n_1249)
);

OA21x2_ASAP7_75t_L g1250 ( 
.A1(n_1145),
.A2(n_928),
.B(n_914),
.Y(n_1250)
);

O2A1O1Ixp5_ASAP7_75t_L g1251 ( 
.A1(n_1044),
.A2(n_926),
.B(n_885),
.C(n_907),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1033),
.B(n_849),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1130),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1178),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1156),
.A2(n_907),
.B(n_887),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1055),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_1068),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1146),
.Y(n_1258)
);

AO22x1_ASAP7_75t_L g1259 ( 
.A1(n_1132),
.A2(n_1000),
.B1(n_997),
.B2(n_958),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1034),
.Y(n_1260)
);

INVxp67_ASAP7_75t_L g1261 ( 
.A(n_1132),
.Y(n_1261)
);

AOI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1188),
.A2(n_926),
.B(n_885),
.Y(n_1262)
);

CKINVDCx6p67_ASAP7_75t_R g1263 ( 
.A(n_1051),
.Y(n_1263)
);

NAND2x1p5_ASAP7_75t_L g1264 ( 
.A(n_1148),
.B(n_941),
.Y(n_1264)
);

NAND2xp33_ASAP7_75t_SL g1265 ( 
.A(n_1095),
.B(n_887),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1178),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1078),
.B(n_1017),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1046),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1042),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1079),
.A2(n_947),
.B1(n_1000),
.B2(n_1001),
.Y(n_1270)
);

AO21x2_ASAP7_75t_L g1271 ( 
.A1(n_1092),
.A2(n_926),
.B(n_983),
.Y(n_1271)
);

BUFx10_ASAP7_75t_L g1272 ( 
.A(n_1034),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1145),
.A2(n_951),
.B(n_867),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1135),
.A2(n_951),
.B(n_867),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1165),
.B(n_988),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1066),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1064),
.A2(n_889),
.B1(n_970),
.B2(n_941),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1152),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1138),
.A2(n_988),
.B1(n_983),
.B2(n_962),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1117),
.B(n_962),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1043),
.B(n_1077),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1069),
.A2(n_943),
.A3(n_979),
.B(n_921),
.Y(n_1282)
);

AOI22x1_ASAP7_75t_L g1283 ( 
.A1(n_1057),
.A2(n_943),
.B1(n_979),
.B2(n_933),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1078),
.B(n_943),
.Y(n_1284)
);

NAND2x1p5_ASAP7_75t_L g1285 ( 
.A(n_1148),
.B(n_970),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1125),
.B(n_951),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1174),
.Y(n_1287)
);

AO21x2_ASAP7_75t_L g1288 ( 
.A1(n_1085),
.A2(n_951),
.B(n_979),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1113),
.B(n_1125),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1135),
.A2(n_933),
.B(n_987),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1136),
.A2(n_933),
.B(n_987),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1034),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1137),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1086),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1136),
.A2(n_987),
.B(n_889),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1154),
.A2(n_837),
.B(n_987),
.C(n_941),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1131),
.B(n_837),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1148),
.Y(n_1298)
);

AOI221xp5_ASAP7_75t_L g1299 ( 
.A1(n_1155),
.A2(n_837),
.B1(n_889),
.B2(n_941),
.C(n_970),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1131),
.B(n_837),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1141),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1046),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1067),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1074),
.A2(n_970),
.B1(n_1045),
.B2(n_1081),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1147),
.B(n_1151),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1164),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1038),
.A2(n_1041),
.B(n_1073),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1155),
.A2(n_1158),
.B1(n_1140),
.B2(n_1102),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1096),
.A2(n_1104),
.B(n_1106),
.Y(n_1309)
);

BUFx12f_ASAP7_75t_L g1310 ( 
.A(n_1148),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1060),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1096),
.A2(n_1104),
.B(n_1106),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1121),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1070),
.A2(n_1142),
.B(n_1093),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1067),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1120),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1110),
.A2(n_1142),
.B(n_1040),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1120),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1157),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1126),
.Y(n_1320)
);

NOR2x1_ASAP7_75t_SL g1321 ( 
.A(n_1185),
.B(n_1184),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1040),
.A2(n_1056),
.B(n_1112),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1152),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1045),
.A2(n_1037),
.B1(n_1050),
.B2(n_1159),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1053),
.B(n_1176),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1102),
.A2(n_1128),
.B1(n_1171),
.B2(n_1169),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1166),
.A2(n_1172),
.B1(n_1116),
.B2(n_1114),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1177),
.B(n_1157),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1182),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1183),
.B(n_1187),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1159),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1056),
.A2(n_1112),
.B(n_1143),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1172),
.B(n_1184),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_1152),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1179),
.A2(n_1180),
.B(n_1091),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1087),
.Y(n_1336)
);

BUFx10_ASAP7_75t_L g1337 ( 
.A(n_1107),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1143),
.A2(n_1094),
.B(n_1161),
.Y(n_1338)
);

AO21x2_ASAP7_75t_L g1339 ( 
.A1(n_1041),
.A2(n_1076),
.B(n_1185),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1084),
.Y(n_1340)
);

INVx3_ASAP7_75t_SL g1341 ( 
.A(n_1163),
.Y(n_1341)
);

INVx4_ASAP7_75t_L g1342 ( 
.A(n_1182),
.Y(n_1342)
);

INVx6_ASAP7_75t_L g1343 ( 
.A(n_1182),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1163),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1186),
.B(n_1076),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1082),
.A2(n_1170),
.B1(n_1105),
.B2(n_1100),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1170),
.A2(n_1089),
.B1(n_1175),
.B2(n_1094),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1053),
.Y(n_1348)
);

OA21x2_ASAP7_75t_L g1349 ( 
.A1(n_1127),
.A2(n_1133),
.B(n_1111),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1053),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1053),
.B(n_1108),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_1098),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1109),
.A2(n_1150),
.B(n_1134),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1124),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1168),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_SL g1356 ( 
.A1(n_1162),
.A2(n_733),
.B1(n_607),
.B2(n_369),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1061),
.A2(n_1027),
.B(n_1145),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1211),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1356),
.A2(n_1220),
.B1(n_1331),
.B2(n_1324),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1201),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1256),
.B(n_1225),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1331),
.A2(n_1343),
.B1(n_1246),
.B2(n_1344),
.Y(n_1362)
);

OAI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1261),
.A2(n_1344),
.B1(n_1227),
.B2(n_1308),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1260),
.B(n_1292),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1310),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1288),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1240),
.B(n_1196),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1236),
.A2(n_1227),
.B1(n_1301),
.B2(n_1265),
.Y(n_1368)
);

OAI222xp33_ASAP7_75t_L g1369 ( 
.A1(n_1206),
.A2(n_1301),
.B1(n_1342),
.B2(n_1230),
.C1(n_1304),
.C2(n_1195),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1302),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1211),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1217),
.B(n_1260),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1281),
.B(n_1305),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1191),
.A2(n_1273),
.B(n_1353),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1265),
.A2(n_1293),
.B1(n_1313),
.B2(n_1255),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1205),
.Y(n_1376)
);

INVx4_ASAP7_75t_L g1377 ( 
.A(n_1310),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1292),
.B(n_1221),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1293),
.A2(n_1320),
.B1(n_1341),
.B2(n_1229),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_1294),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1272),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1200),
.A2(n_1252),
.B1(n_1326),
.B2(n_1341),
.Y(n_1382)
);

CKINVDCx16_ASAP7_75t_R g1383 ( 
.A(n_1212),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1223),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1269),
.B(n_1287),
.Y(n_1385)
);

INVx6_ASAP7_75t_L g1386 ( 
.A(n_1272),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1303),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1343),
.A2(n_1270),
.B1(n_1263),
.B2(n_1192),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1232),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1189),
.A2(n_1343),
.B1(n_1346),
.B2(n_1299),
.Y(n_1390)
);

INVx4_ASAP7_75t_L g1391 ( 
.A(n_1205),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1234),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1217),
.B(n_1284),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1272),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_R g1395 ( 
.A(n_1233),
.B(n_1257),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1343),
.A2(n_1342),
.B1(n_1333),
.B2(n_1352),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1244),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1303),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1212),
.A2(n_1330),
.B1(n_1294),
.B2(n_1296),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1327),
.A2(n_1352),
.B1(n_1333),
.B2(n_1263),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1335),
.A2(n_1355),
.B(n_1190),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_1244),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1239),
.B(n_1245),
.Y(n_1403)
);

INVx3_ASAP7_75t_SL g1404 ( 
.A(n_1257),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1288),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1279),
.A2(n_1347),
.B1(n_1218),
.B2(n_1192),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1253),
.B(n_1258),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_1204),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1288),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1306),
.B(n_1241),
.Y(n_1410)
);

INVx4_ASAP7_75t_L g1411 ( 
.A(n_1323),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1191),
.A2(n_1273),
.B(n_1353),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1355),
.A2(n_1190),
.B(n_1208),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1316),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1311),
.A2(n_1233),
.B1(n_1325),
.B2(n_1348),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1325),
.A2(n_1348),
.B1(n_1342),
.B2(n_1250),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1241),
.B(n_1284),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1207),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1192),
.A2(n_1280),
.B1(n_1275),
.B2(n_1250),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1315),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1318),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1315),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1259),
.B(n_1336),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1207),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1244),
.Y(n_1425)
);

OAI221xp5_ASAP7_75t_L g1426 ( 
.A1(n_1251),
.A2(n_1289),
.B1(n_1250),
.B2(n_1203),
.C(n_1328),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1207),
.Y(n_1427)
);

AO21x1_ASAP7_75t_L g1428 ( 
.A1(n_1345),
.A2(n_1247),
.B(n_1351),
.Y(n_1428)
);

INVx5_ASAP7_75t_L g1429 ( 
.A(n_1192),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1268),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1250),
.A2(n_1350),
.B1(n_1336),
.B2(n_1222),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1259),
.B(n_1242),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1207),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1323),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1298),
.Y(n_1435)
);

AOI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1198),
.A2(n_1351),
.B1(n_1329),
.B2(n_1209),
.C(n_1340),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1319),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1286),
.B(n_1224),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1268),
.B(n_1242),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1244),
.B(n_1276),
.Y(n_1440)
);

OR2x6_ASAP7_75t_L g1441 ( 
.A(n_1247),
.B(n_1235),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1286),
.B(n_1297),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1323),
.Y(n_1443)
);

AOI332xp33_ASAP7_75t_L g1444 ( 
.A1(n_1297),
.A2(n_1345),
.A3(n_1222),
.B1(n_1267),
.B2(n_1224),
.B3(n_1278),
.C1(n_1300),
.C2(n_1319),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1244),
.Y(n_1445)
);

OR2x6_ASAP7_75t_L g1446 ( 
.A(n_1199),
.B(n_1214),
.Y(n_1446)
);

NAND3xp33_ASAP7_75t_L g1447 ( 
.A(n_1283),
.B(n_1340),
.C(n_1276),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1202),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1340),
.A2(n_1267),
.B1(n_1224),
.B2(n_1209),
.Y(n_1449)
);

AND2x4_ASAP7_75t_L g1450 ( 
.A(n_1267),
.B(n_1276),
.Y(n_1450)
);

AOI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1340),
.A2(n_1345),
.B1(n_1276),
.B2(n_1235),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1276),
.B(n_1340),
.Y(n_1452)
);

NAND2x1_ASAP7_75t_L g1453 ( 
.A(n_1194),
.B(n_1216),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1277),
.A2(n_1194),
.B(n_1216),
.C(n_1278),
.Y(n_1454)
);

OAI21xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1334),
.A2(n_1278),
.B(n_1295),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1202),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1210),
.Y(n_1457)
);

OAI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1199),
.A2(n_1214),
.B1(n_1235),
.B2(n_1334),
.Y(n_1458)
);

CKINVDCx6p67_ASAP7_75t_R g1459 ( 
.A(n_1337),
.Y(n_1459)
);

NAND2xp33_ASAP7_75t_SL g1460 ( 
.A(n_1323),
.B(n_1199),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1298),
.B(n_1228),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1317),
.A2(n_1332),
.B(n_1290),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1210),
.Y(n_1463)
);

A2O1A1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1214),
.A2(n_1197),
.B(n_1295),
.C(n_1290),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1209),
.A2(n_1266),
.B1(n_1231),
.B2(n_1243),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1231),
.A2(n_1266),
.B1(n_1243),
.B2(n_1254),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1237),
.Y(n_1467)
);

INVx4_ASAP7_75t_L g1468 ( 
.A(n_1323),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1264),
.Y(n_1469)
);

AO32x2_ASAP7_75t_L g1470 ( 
.A1(n_1248),
.A2(n_1228),
.A3(n_1321),
.B1(n_1254),
.B2(n_1237),
.Y(n_1470)
);

AOI21xp33_ASAP7_75t_L g1471 ( 
.A1(n_1271),
.A2(n_1307),
.B(n_1349),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1271),
.A2(n_1339),
.B1(n_1307),
.B2(n_1283),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1271),
.A2(n_1339),
.B1(n_1307),
.B2(n_1337),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1213),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1193),
.B(n_1226),
.Y(n_1475)
);

BUFx4f_ASAP7_75t_SL g1476 ( 
.A(n_1337),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1197),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1228),
.B(n_1248),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1228),
.B(n_1248),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1228),
.B(n_1339),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1264),
.A2(n_1285),
.B1(n_1349),
.B2(n_1238),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1282),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1354),
.Y(n_1483)
);

AOI221xp5_ASAP7_75t_L g1484 ( 
.A1(n_1354),
.A2(n_1248),
.B1(n_1264),
.B2(n_1285),
.C(n_1238),
.Y(n_1484)
);

NAND2xp33_ASAP7_75t_R g1485 ( 
.A(n_1349),
.B(n_1338),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1213),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1349),
.A2(n_1285),
.B1(n_1219),
.B2(n_1338),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1193),
.B(n_1226),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1215),
.A2(n_1219),
.B1(n_1357),
.B2(n_1338),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1321),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1226),
.B(n_1248),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1215),
.A2(n_1357),
.B1(n_1338),
.B2(n_1249),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1226),
.B(n_1282),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1262),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1274),
.A2(n_1291),
.B1(n_1226),
.B2(n_1332),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1282),
.B(n_1274),
.Y(n_1496)
);

NAND2xp33_ASAP7_75t_R g1497 ( 
.A(n_1357),
.B(n_1314),
.Y(n_1497)
);

CKINVDCx11_ASAP7_75t_R g1498 ( 
.A(n_1282),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1249),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1291),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1322),
.B(n_1317),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1314),
.A2(n_1357),
.B(n_1322),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1309),
.Y(n_1503)
);

CKINVDCx20_ASAP7_75t_R g1504 ( 
.A(n_1314),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1309),
.A2(n_1312),
.B(n_1314),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1312),
.Y(n_1506)
);

NAND2xp33_ASAP7_75t_R g1507 ( 
.A(n_1227),
.B(n_989),
.Y(n_1507)
);

INVx3_ASAP7_75t_L g1508 ( 
.A(n_1310),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1310),
.Y(n_1509)
);

INVx4_ASAP7_75t_L g1510 ( 
.A(n_1310),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1201),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1201),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1430),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1359),
.A2(n_1363),
.B1(n_1400),
.B2(n_1390),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1373),
.B(n_1361),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1359),
.A2(n_1363),
.B1(n_1368),
.B2(n_1396),
.Y(n_1516)
);

OAI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1382),
.A2(n_1399),
.B1(n_1406),
.B2(n_1383),
.Y(n_1517)
);

BUFx2_ASAP7_75t_L g1518 ( 
.A(n_1455),
.Y(n_1518)
);

AOI222xp33_ASAP7_75t_L g1519 ( 
.A1(n_1369),
.A2(n_1368),
.B1(n_1375),
.B2(n_1379),
.C1(n_1388),
.C2(n_1478),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1442),
.B(n_1393),
.Y(n_1520)
);

AOI211xp5_ASAP7_75t_L g1521 ( 
.A1(n_1388),
.A2(n_1419),
.B(n_1426),
.C(n_1367),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1401),
.A2(n_1502),
.B(n_1471),
.Y(n_1522)
);

AOI221xp5_ASAP7_75t_L g1523 ( 
.A1(n_1375),
.A2(n_1379),
.B1(n_1360),
.B2(n_1392),
.C(n_1512),
.Y(n_1523)
);

OAI211xp5_ASAP7_75t_L g1524 ( 
.A1(n_1395),
.A2(n_1362),
.B(n_1444),
.C(n_1385),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1476),
.A2(n_1459),
.B1(n_1380),
.B2(n_1504),
.Y(n_1525)
);

AOI21xp33_ASAP7_75t_L g1526 ( 
.A1(n_1423),
.A2(n_1507),
.B(n_1483),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1413),
.A2(n_1412),
.B(n_1374),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1376),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1476),
.A2(n_1504),
.B1(n_1415),
.B2(n_1404),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1404),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1414),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1408),
.Y(n_1532)
);

OAI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1415),
.A2(n_1473),
.B1(n_1431),
.B2(n_1389),
.C(n_1384),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1489),
.A2(n_1492),
.B(n_1462),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1358),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_SL g1536 ( 
.A1(n_1479),
.A2(n_1395),
.B1(n_1493),
.B2(n_1429),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1378),
.B(n_1403),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1435),
.A2(n_1365),
.B1(n_1510),
.B2(n_1377),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1377),
.A2(n_1510),
.B1(n_1509),
.B2(n_1508),
.Y(n_1539)
);

INVx2_ASAP7_75t_SL g1540 ( 
.A(n_1429),
.Y(n_1540)
);

A2O1A1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1436),
.A2(n_1416),
.B(n_1410),
.C(n_1473),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1393),
.B(n_1511),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1429),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1498),
.A2(n_1428),
.B1(n_1491),
.B2(n_1393),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1397),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1372),
.B(n_1416),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1461),
.B(n_1480),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1498),
.A2(n_1421),
.B1(n_1372),
.B2(n_1432),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1489),
.A2(n_1492),
.B(n_1472),
.Y(n_1549)
);

OAI221xp5_ASAP7_75t_L g1550 ( 
.A1(n_1431),
.A2(n_1472),
.B1(n_1407),
.B2(n_1449),
.C(n_1507),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1417),
.B(n_1364),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1372),
.A2(n_1438),
.B1(n_1475),
.B2(n_1488),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1438),
.A2(n_1475),
.B1(n_1488),
.B2(n_1449),
.Y(n_1553)
);

OAI221xp5_ASAP7_75t_L g1554 ( 
.A1(n_1391),
.A2(n_1484),
.B1(n_1485),
.B2(n_1495),
.C(n_1427),
.Y(n_1554)
);

OAI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1391),
.A2(n_1485),
.B1(n_1487),
.B2(n_1424),
.C(n_1451),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1438),
.A2(n_1475),
.B1(n_1429),
.B2(n_1420),
.Y(n_1556)
);

OAI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1358),
.A2(n_1371),
.B1(n_1386),
.B2(n_1381),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1387),
.A2(n_1420),
.B1(n_1422),
.B2(n_1437),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_SL g1559 ( 
.A1(n_1490),
.A2(n_1482),
.B1(n_1371),
.B2(n_1386),
.Y(n_1559)
);

BUFx8_ASAP7_75t_SL g1560 ( 
.A(n_1433),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1387),
.A2(n_1422),
.B1(n_1437),
.B2(n_1398),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1398),
.A2(n_1457),
.B1(n_1467),
.B2(n_1456),
.Y(n_1562)
);

AO31x2_ASAP7_75t_L g1563 ( 
.A1(n_1464),
.A2(n_1463),
.A3(n_1477),
.B(n_1474),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1448),
.A2(n_1450),
.B1(n_1465),
.B2(n_1366),
.Y(n_1564)
);

OAI21xp33_ASAP7_75t_L g1565 ( 
.A1(n_1503),
.A2(n_1506),
.B(n_1496),
.Y(n_1565)
);

OAI222xp33_ASAP7_75t_L g1566 ( 
.A1(n_1439),
.A2(n_1441),
.B1(n_1465),
.B2(n_1463),
.C1(n_1466),
.C2(n_1452),
.Y(n_1566)
);

NAND2x1_ASAP7_75t_L g1567 ( 
.A(n_1446),
.B(n_1425),
.Y(n_1567)
);

OAI211xp5_ASAP7_75t_L g1568 ( 
.A1(n_1454),
.A2(n_1453),
.B(n_1499),
.C(n_1434),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1418),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1482),
.B(n_1500),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1440),
.Y(n_1571)
);

OAI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1381),
.A2(n_1447),
.B1(n_1418),
.B2(n_1441),
.Y(n_1572)
);

BUFx12f_ASAP7_75t_L g1573 ( 
.A(n_1397),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1450),
.A2(n_1366),
.B1(n_1409),
.B2(n_1405),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1397),
.Y(n_1575)
);

OAI221xp5_ASAP7_75t_L g1576 ( 
.A1(n_1394),
.A2(n_1497),
.B1(n_1460),
.B2(n_1409),
.C(n_1405),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1470),
.B(n_1397),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1460),
.A2(n_1481),
.B(n_1458),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1470),
.B(n_1445),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1441),
.A2(n_1466),
.B1(n_1494),
.B2(n_1381),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1402),
.B(n_1445),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1458),
.A2(n_1481),
.B(n_1464),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_SL g1583 ( 
.A1(n_1381),
.A2(n_1494),
.B1(n_1469),
.B2(n_1394),
.Y(n_1583)
);

CKINVDCx11_ASAP7_75t_R g1584 ( 
.A(n_1446),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1411),
.A2(n_1468),
.B1(n_1443),
.B2(n_1434),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1494),
.A2(n_1402),
.B1(n_1425),
.B2(n_1411),
.Y(n_1586)
);

OA21x2_ASAP7_75t_L g1587 ( 
.A1(n_1486),
.A2(n_1501),
.B(n_1497),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1470),
.B(n_1501),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1470),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1443),
.B(n_1468),
.Y(n_1590)
);

OAI221xp5_ASAP7_75t_L g1591 ( 
.A1(n_1505),
.A2(n_733),
.B1(n_1022),
.B2(n_799),
.C(n_945),
.Y(n_1591)
);

OAI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1505),
.A2(n_733),
.B1(n_1022),
.B2(n_799),
.C(n_945),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1367),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1359),
.A2(n_733),
.B1(n_1018),
.B2(n_1356),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1442),
.B(n_1393),
.Y(n_1595)
);

AOI222xp33_ASAP7_75t_L g1596 ( 
.A1(n_1359),
.A2(n_607),
.B1(n_733),
.B2(n_709),
.C1(n_1369),
.C2(n_690),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1359),
.A2(n_733),
.B1(n_1018),
.B2(n_1356),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1373),
.B(n_1361),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1430),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1373),
.B(n_1361),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1375),
.A2(n_1331),
.B1(n_683),
.B2(n_1356),
.Y(n_1601)
);

OAI211xp5_ASAP7_75t_L g1602 ( 
.A1(n_1375),
.A2(n_799),
.B(n_691),
.C(n_1149),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1367),
.Y(n_1603)
);

AND2x4_ASAP7_75t_SL g1604 ( 
.A(n_1450),
.B(n_1438),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1367),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_1383),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1413),
.A2(n_1401),
.B(n_1374),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1359),
.A2(n_733),
.B1(n_1018),
.B2(n_1356),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1359),
.A2(n_733),
.B1(n_1018),
.B2(n_1356),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1359),
.A2(n_733),
.B1(n_1018),
.B2(n_1356),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1442),
.B(n_1393),
.Y(n_1611)
);

AOI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1363),
.A2(n_733),
.B1(n_799),
.B2(n_690),
.C(n_536),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1430),
.Y(n_1613)
);

OAI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1375),
.A2(n_733),
.B1(n_1022),
.B2(n_799),
.C(n_945),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1359),
.A2(n_733),
.B1(n_1018),
.B2(n_1356),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1359),
.A2(n_733),
.B1(n_1018),
.B2(n_1356),
.Y(n_1616)
);

O2A1O1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1382),
.A2(n_733),
.B(n_835),
.C(n_799),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1359),
.A2(n_733),
.B1(n_1018),
.B2(n_1356),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1375),
.A2(n_1331),
.B1(n_683),
.B2(n_1356),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1359),
.A2(n_733),
.B1(n_1018),
.B2(n_1356),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_SL g1621 ( 
.A1(n_1400),
.A2(n_733),
.B1(n_1331),
.B2(n_607),
.Y(n_1621)
);

NAND3xp33_ASAP7_75t_L g1622 ( 
.A(n_1375),
.B(n_733),
.C(n_1382),
.Y(n_1622)
);

AO221x2_ASAP7_75t_L g1623 ( 
.A1(n_1363),
.A2(n_1382),
.B1(n_1400),
.B2(n_1246),
.C(n_1369),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1375),
.A2(n_1331),
.B1(n_683),
.B2(n_1356),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1370),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1430),
.Y(n_1626)
);

AOI222xp33_ASAP7_75t_L g1627 ( 
.A1(n_1359),
.A2(n_607),
.B1(n_733),
.B2(n_709),
.C1(n_1369),
.C2(n_690),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1358),
.Y(n_1628)
);

INVx3_ASAP7_75t_L g1629 ( 
.A(n_1397),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1375),
.A2(n_1331),
.B1(n_683),
.B2(n_1356),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1430),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1430),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1588),
.B(n_1518),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1528),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1587),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1513),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1513),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1588),
.B(n_1518),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1535),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1577),
.B(n_1579),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1579),
.B(n_1577),
.Y(n_1641)
);

OR2x6_ASAP7_75t_SL g1642 ( 
.A(n_1529),
.B(n_1622),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1587),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1599),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1582),
.B(n_1552),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1599),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1587),
.B(n_1549),
.Y(n_1647)
);

AOI221xp5_ASAP7_75t_L g1648 ( 
.A1(n_1612),
.A2(n_1617),
.B1(n_1614),
.B2(n_1619),
.C(n_1630),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1587),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1593),
.B(n_1603),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1549),
.B(n_1534),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1605),
.B(n_1613),
.Y(n_1652)
);

NOR2x1_ASAP7_75t_L g1653 ( 
.A(n_1554),
.B(n_1535),
.Y(n_1653)
);

AOI21xp33_ASAP7_75t_L g1654 ( 
.A1(n_1596),
.A2(n_1627),
.B(n_1602),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1534),
.B(n_1589),
.Y(n_1655)
);

INVx3_ASAP7_75t_L g1656 ( 
.A(n_1534),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1626),
.B(n_1631),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1623),
.A2(n_1610),
.B1(n_1594),
.B2(n_1608),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1623),
.A2(n_1597),
.B1(n_1609),
.B2(n_1615),
.Y(n_1659)
);

AND2x2_ASAP7_75t_SL g1660 ( 
.A(n_1514),
.B(n_1516),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1589),
.B(n_1547),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1547),
.B(n_1570),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1570),
.B(n_1537),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1534),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1628),
.Y(n_1665)
);

OR2x6_ASAP7_75t_L g1666 ( 
.A(n_1578),
.B(n_1546),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1576),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1522),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1571),
.B(n_1632),
.Y(n_1669)
);

NAND2xp33_ASAP7_75t_SL g1670 ( 
.A(n_1606),
.B(n_1525),
.Y(n_1670)
);

AND2x4_ASAP7_75t_SL g1671 ( 
.A(n_1542),
.B(n_1520),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1531),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1522),
.B(n_1563),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1623),
.A2(n_1618),
.B1(n_1616),
.B2(n_1620),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1531),
.Y(n_1675)
);

AO21x2_ASAP7_75t_L g1676 ( 
.A1(n_1541),
.A2(n_1566),
.B(n_1607),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1522),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_1575),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1563),
.B(n_1520),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1515),
.B(n_1598),
.Y(n_1680)
);

AOI211xp5_ASAP7_75t_L g1681 ( 
.A1(n_1517),
.A2(n_1601),
.B(n_1624),
.C(n_1592),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1551),
.B(n_1600),
.Y(n_1682)
);

AOI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1591),
.A2(n_1621),
.B1(n_1524),
.B2(n_1521),
.C(n_1523),
.Y(n_1683)
);

OAI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1654),
.A2(n_1623),
.B1(n_1550),
.B2(n_1533),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_SL g1685 ( 
.A1(n_1660),
.A2(n_1519),
.B1(n_1555),
.B2(n_1611),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1633),
.B(n_1611),
.Y(n_1686)
);

OA21x2_ASAP7_75t_L g1687 ( 
.A1(n_1649),
.A2(n_1607),
.B(n_1527),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1648),
.A2(n_1606),
.B1(n_1530),
.B2(n_1536),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1654),
.A2(n_1683),
.B1(n_1660),
.B2(n_1648),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1660),
.A2(n_1548),
.B1(n_1584),
.B2(n_1544),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1681),
.A2(n_1586),
.B1(n_1575),
.B2(n_1559),
.Y(n_1691)
);

AOI33xp33_ASAP7_75t_L g1692 ( 
.A1(n_1681),
.A2(n_1595),
.A3(n_1583),
.B1(n_1574),
.B2(n_1564),
.B3(n_1553),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1636),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1636),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1683),
.A2(n_1526),
.B1(n_1580),
.B2(n_1556),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1637),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1667),
.A2(n_1565),
.B1(n_1538),
.B2(n_1572),
.C(n_1539),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1637),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1679),
.B(n_1640),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_SL g1700 ( 
.A1(n_1660),
.A2(n_1645),
.B1(n_1649),
.B2(n_1676),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1638),
.B(n_1595),
.Y(n_1701)
);

NOR2x1_ASAP7_75t_L g1702 ( 
.A(n_1639),
.B(n_1568),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1633),
.B(n_1625),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1642),
.A2(n_1532),
.B1(n_1567),
.B2(n_1569),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1644),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1665),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1662),
.Y(n_1707)
);

OAI31xp33_ASAP7_75t_L g1708 ( 
.A1(n_1658),
.A2(n_1557),
.A3(n_1604),
.B(n_1569),
.Y(n_1708)
);

OAI33xp33_ASAP7_75t_L g1709 ( 
.A1(n_1667),
.A2(n_1650),
.A3(n_1652),
.B1(n_1680),
.B2(n_1682),
.B3(n_1661),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1662),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1644),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1662),
.B(n_1581),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1646),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1658),
.A2(n_1584),
.B1(n_1562),
.B2(n_1561),
.Y(n_1714)
);

AO21x2_ASAP7_75t_L g1715 ( 
.A1(n_1676),
.A2(n_1590),
.B(n_1585),
.Y(n_1715)
);

OAI221xp5_ASAP7_75t_L g1716 ( 
.A1(n_1659),
.A2(n_1558),
.B1(n_1543),
.B2(n_1540),
.C(n_1629),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1679),
.B(n_1640),
.Y(n_1717)
);

A2O1A1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1659),
.A2(n_1674),
.B(n_1645),
.C(n_1653),
.Y(n_1718)
);

AOI31xp33_ASAP7_75t_SL g1719 ( 
.A1(n_1633),
.A2(n_1560),
.A3(n_1532),
.B(n_1528),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1680),
.B(n_1629),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1638),
.B(n_1545),
.Y(n_1721)
);

HB1xp67_ASAP7_75t_L g1722 ( 
.A(n_1661),
.Y(n_1722)
);

NOR4xp25_ASAP7_75t_SL g1723 ( 
.A(n_1670),
.B(n_1560),
.C(n_1573),
.D(n_1545),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1661),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1634),
.B(n_1573),
.Y(n_1725)
);

INVxp67_ASAP7_75t_L g1726 ( 
.A(n_1665),
.Y(n_1726)
);

INVx4_ASAP7_75t_L g1727 ( 
.A(n_1715),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1693),
.Y(n_1728)
);

INVxp67_ASAP7_75t_SL g1729 ( 
.A(n_1687),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1693),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1699),
.B(n_1640),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1699),
.B(n_1640),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1707),
.B(n_1655),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1699),
.B(n_1640),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1699),
.B(n_1641),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1717),
.B(n_1641),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1710),
.B(n_1650),
.Y(n_1737)
);

NAND3xp33_ASAP7_75t_L g1738 ( 
.A(n_1689),
.B(n_1674),
.C(n_1673),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1694),
.Y(n_1739)
);

NOR3xp33_ASAP7_75t_L g1740 ( 
.A(n_1684),
.B(n_1668),
.C(n_1677),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1717),
.B(n_1655),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1694),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1722),
.B(n_1655),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1717),
.B(n_1635),
.Y(n_1744)
);

NOR3xp33_ASAP7_75t_L g1745 ( 
.A(n_1718),
.B(n_1668),
.C(n_1677),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1696),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1717),
.B(n_1635),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1696),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1701),
.B(n_1679),
.Y(n_1749)
);

OA21x2_ASAP7_75t_L g1750 ( 
.A1(n_1697),
.A2(n_1649),
.B(n_1673),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1724),
.B(n_1652),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1698),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1701),
.B(n_1651),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1698),
.B(n_1682),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1703),
.B(n_1663),
.Y(n_1755)
);

OR2x2_ASAP7_75t_SL g1756 ( 
.A(n_1686),
.B(n_1682),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1721),
.B(n_1647),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1705),
.B(n_1672),
.Y(n_1758)
);

OAI33xp33_ASAP7_75t_L g1759 ( 
.A1(n_1688),
.A2(n_1669),
.A3(n_1657),
.B1(n_1663),
.B2(n_1675),
.B3(n_1672),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1721),
.B(n_1647),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1711),
.B(n_1675),
.Y(n_1761)
);

AND2x4_ASAP7_75t_SL g1762 ( 
.A(n_1690),
.B(n_1666),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1686),
.B(n_1669),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_SL g1764 ( 
.A(n_1738),
.B(n_1708),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1728),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1728),
.Y(n_1766)
);

INVxp67_ASAP7_75t_L g1767 ( 
.A(n_1740),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1749),
.B(n_1706),
.Y(n_1768)
);

INVxp67_ASAP7_75t_SL g1769 ( 
.A(n_1740),
.Y(n_1769)
);

AND2x2_ASAP7_75t_SL g1770 ( 
.A(n_1750),
.B(n_1645),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1759),
.B(n_1725),
.Y(n_1771)
);

NOR2xp67_ASAP7_75t_SL g1772 ( 
.A(n_1750),
.B(n_1716),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1730),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1730),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1739),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1754),
.B(n_1711),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1749),
.B(n_1731),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1756),
.B(n_1712),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1739),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1750),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1742),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1750),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1742),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1750),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1746),
.Y(n_1785)
);

NAND2x1_ASAP7_75t_L g1786 ( 
.A(n_1731),
.B(n_1702),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1749),
.B(n_1726),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1756),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1746),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1754),
.B(n_1713),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1748),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1737),
.B(n_1720),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1751),
.B(n_1713),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1737),
.Y(n_1794)
);

NOR2x1_ASAP7_75t_L g1795 ( 
.A(n_1727),
.B(n_1719),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1731),
.B(n_1671),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1731),
.B(n_1671),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1763),
.B(n_1669),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1748),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1752),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1745),
.B(n_1702),
.Y(n_1801)
);

NAND2x1_ASAP7_75t_L g1802 ( 
.A(n_1731),
.B(n_1666),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1770),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1798),
.B(n_1763),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1777),
.B(n_1744),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1775),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1767),
.B(n_1745),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1798),
.B(n_1763),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1777),
.B(n_1732),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1795),
.B(n_1732),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1767),
.B(n_1738),
.Y(n_1811)
);

NOR3xp33_ASAP7_75t_L g1812 ( 
.A(n_1769),
.B(n_1727),
.C(n_1759),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1795),
.B(n_1732),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1794),
.B(n_1751),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1775),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1791),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_SL g1817 ( 
.A(n_1770),
.B(n_1708),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1770),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1771),
.B(n_1709),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1780),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1786),
.B(n_1734),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1764),
.A2(n_1685),
.B1(n_1700),
.B2(n_1645),
.Y(n_1822)
);

NOR2x1_ASAP7_75t_L g1823 ( 
.A(n_1801),
.B(n_1727),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1793),
.B(n_1733),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1769),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1778),
.B(n_1753),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1791),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1765),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1793),
.B(n_1733),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1778),
.B(n_1753),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1765),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1780),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1766),
.Y(n_1833)
);

INVx4_ASAP7_75t_L g1834 ( 
.A(n_1780),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1792),
.B(n_1743),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1786),
.B(n_1734),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1766),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1782),
.Y(n_1838)
);

OAI21x1_ASAP7_75t_SL g1839 ( 
.A1(n_1788),
.A2(n_1704),
.B(n_1727),
.Y(n_1839)
);

OAI211xp5_ASAP7_75t_SL g1840 ( 
.A1(n_1782),
.A2(n_1729),
.B(n_1761),
.C(n_1758),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1773),
.Y(n_1841)
);

NOR4xp25_ASAP7_75t_SL g1842 ( 
.A(n_1772),
.B(n_1670),
.C(n_1729),
.D(n_1678),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1773),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1782),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1774),
.Y(n_1845)
);

OAI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1819),
.A2(n_1764),
.B1(n_1772),
.B2(n_1784),
.C(n_1788),
.Y(n_1846)
);

NAND2xp33_ASAP7_75t_L g1847 ( 
.A(n_1825),
.B(n_1788),
.Y(n_1847)
);

OAI221xp5_ASAP7_75t_SL g1848 ( 
.A1(n_1807),
.A2(n_1784),
.B1(n_1692),
.B2(n_1690),
.C(n_1666),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1811),
.B(n_1792),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1837),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1812),
.B(n_1768),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1834),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1845),
.Y(n_1853)
);

OAI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1817),
.A2(n_1784),
.B1(n_1727),
.B2(n_1802),
.C(n_1695),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1815),
.Y(n_1855)
);

XOR2xp5_ASAP7_75t_L g1856 ( 
.A(n_1822),
.B(n_1691),
.Y(n_1856)
);

INVx2_ASAP7_75t_SL g1857 ( 
.A(n_1814),
.Y(n_1857)
);

OAI21xp33_ASAP7_75t_SL g1858 ( 
.A1(n_1810),
.A2(n_1735),
.B(n_1736),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1834),
.Y(n_1859)
);

OAI21xp5_ASAP7_75t_SL g1860 ( 
.A1(n_1823),
.A2(n_1653),
.B(n_1762),
.Y(n_1860)
);

OAI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1822),
.A2(n_1642),
.B1(n_1666),
.B2(n_1802),
.Y(n_1861)
);

OAI21xp33_ASAP7_75t_SL g1862 ( 
.A1(n_1810),
.A2(n_1736),
.B(n_1735),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1814),
.B(n_1768),
.Y(n_1863)
);

INVxp67_ASAP7_75t_SL g1864 ( 
.A(n_1820),
.Y(n_1864)
);

INVxp67_ASAP7_75t_L g1865 ( 
.A(n_1806),
.Y(n_1865)
);

INVx1_ASAP7_75t_SL g1866 ( 
.A(n_1803),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1828),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1804),
.B(n_1776),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1809),
.B(n_1796),
.Y(n_1869)
);

OAI211xp5_ASAP7_75t_L g1870 ( 
.A1(n_1842),
.A2(n_1723),
.B(n_1678),
.C(n_1677),
.Y(n_1870)
);

NAND2xp33_ASAP7_75t_SL g1871 ( 
.A(n_1842),
.B(n_1796),
.Y(n_1871)
);

AOI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1803),
.A2(n_1676),
.B1(n_1647),
.B2(n_1645),
.Y(n_1872)
);

O2A1O1Ixp33_ASAP7_75t_R g1873 ( 
.A1(n_1804),
.A2(n_1776),
.B(n_1790),
.C(n_1755),
.Y(n_1873)
);

OAI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1823),
.A2(n_1642),
.B1(n_1818),
.B2(n_1803),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1808),
.B(n_1790),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1828),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1806),
.B(n_1787),
.Y(n_1877)
);

AOI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1818),
.A2(n_1676),
.B1(n_1762),
.B2(n_1666),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1805),
.Y(n_1879)
);

NOR2x1_ASAP7_75t_L g1880 ( 
.A(n_1834),
.B(n_1774),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1816),
.B(n_1787),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1867),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1876),
.Y(n_1883)
);

AOI211xp5_ASAP7_75t_L g1884 ( 
.A1(n_1874),
.A2(n_1840),
.B(n_1818),
.C(n_1813),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1856),
.A2(n_1839),
.B(n_1832),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1850),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1879),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1853),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1855),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_L g1890 ( 
.A(n_1849),
.B(n_1808),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1879),
.Y(n_1891)
);

INVx1_ASAP7_75t_SL g1892 ( 
.A(n_1847),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1846),
.A2(n_1826),
.B1(n_1830),
.B2(n_1813),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1849),
.B(n_1834),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1880),
.Y(n_1895)
);

INVxp33_ASAP7_75t_L g1896 ( 
.A(n_1852),
.Y(n_1896)
);

AOI211xp5_ASAP7_75t_L g1897 ( 
.A1(n_1873),
.A2(n_1827),
.B(n_1816),
.C(n_1832),
.Y(n_1897)
);

AOI332xp33_ASAP7_75t_L g1898 ( 
.A1(n_1851),
.A2(n_1827),
.A3(n_1843),
.B1(n_1841),
.B2(n_1831),
.B3(n_1833),
.C1(n_1832),
.C2(n_1820),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1857),
.B(n_1835),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1863),
.B(n_1835),
.Y(n_1900)
);

A2O1A1Ixp33_ASAP7_75t_L g1901 ( 
.A1(n_1848),
.A2(n_1844),
.B(n_1820),
.C(n_1838),
.Y(n_1901)
);

NAND3xp33_ASAP7_75t_L g1902 ( 
.A(n_1865),
.B(n_1844),
.C(n_1838),
.Y(n_1902)
);

AOI221xp5_ASAP7_75t_L g1903 ( 
.A1(n_1854),
.A2(n_1839),
.B1(n_1844),
.B2(n_1838),
.C(n_1843),
.Y(n_1903)
);

INVx1_ASAP7_75t_SL g1904 ( 
.A(n_1866),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1864),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1868),
.B(n_1824),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1861),
.A2(n_1871),
.B(n_1860),
.Y(n_1907)
);

INVx1_ASAP7_75t_SL g1908 ( 
.A(n_1892),
.Y(n_1908)
);

NAND2xp33_ASAP7_75t_R g1909 ( 
.A(n_1907),
.B(n_1852),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1905),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1905),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_1887),
.Y(n_1912)
);

XNOR2xp5_ASAP7_75t_L g1913 ( 
.A(n_1904),
.B(n_1861),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1882),
.Y(n_1914)
);

INVxp67_ASAP7_75t_L g1915 ( 
.A(n_1887),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1882),
.Y(n_1916)
);

XOR2x2_ASAP7_75t_L g1917 ( 
.A(n_1885),
.B(n_1872),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1902),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1883),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1890),
.B(n_1865),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1900),
.B(n_1875),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1906),
.B(n_1869),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1889),
.Y(n_1923)
);

BUFx2_ASAP7_75t_L g1924 ( 
.A(n_1891),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1891),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1886),
.Y(n_1926)
);

XOR2x2_ASAP7_75t_L g1927 ( 
.A(n_1903),
.B(n_1878),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1922),
.B(n_1899),
.Y(n_1928)
);

OAI21xp33_ASAP7_75t_L g1929 ( 
.A1(n_1908),
.A2(n_1893),
.B(n_1894),
.Y(n_1929)
);

AOI221x1_ASAP7_75t_L g1930 ( 
.A1(n_1918),
.A2(n_1888),
.B1(n_1895),
.B2(n_1901),
.C(n_1871),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1917),
.A2(n_1901),
.B1(n_1884),
.B2(n_1864),
.Y(n_1931)
);

NAND4xp25_ASAP7_75t_L g1932 ( 
.A(n_1909),
.B(n_1897),
.C(n_1895),
.D(n_1859),
.Y(n_1932)
);

NOR2x1_ASAP7_75t_L g1933 ( 
.A(n_1912),
.B(n_1859),
.Y(n_1933)
);

NAND3xp33_ASAP7_75t_SL g1934 ( 
.A(n_1918),
.B(n_1898),
.C(n_1896),
.Y(n_1934)
);

AOI22xp33_ASAP7_75t_L g1935 ( 
.A1(n_1927),
.A2(n_1896),
.B1(n_1666),
.B2(n_1635),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1913),
.A2(n_1881),
.B(n_1877),
.Y(n_1936)
);

NOR4xp75_ASAP7_75t_L g1937 ( 
.A(n_1920),
.B(n_1821),
.C(n_1836),
.D(n_1809),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1912),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1924),
.Y(n_1939)
);

AOI322xp5_ASAP7_75t_L g1940 ( 
.A1(n_1934),
.A2(n_1910),
.A3(n_1911),
.B1(n_1917),
.B2(n_1923),
.C1(n_1926),
.C2(n_1916),
.Y(n_1940)
);

AOI211xp5_ASAP7_75t_L g1941 ( 
.A1(n_1932),
.A2(n_1913),
.B(n_1915),
.C(n_1924),
.Y(n_1941)
);

AOI311xp33_ASAP7_75t_L g1942 ( 
.A1(n_1938),
.A2(n_1919),
.A3(n_1914),
.B(n_1858),
.C(n_1862),
.Y(n_1942)
);

AOI221x1_ASAP7_75t_L g1943 ( 
.A1(n_1939),
.A2(n_1925),
.B1(n_1922),
.B2(n_1927),
.C(n_1831),
.Y(n_1943)
);

OAI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1930),
.A2(n_1931),
.B(n_1936),
.Y(n_1944)
);

AOI211xp5_ASAP7_75t_L g1945 ( 
.A1(n_1929),
.A2(n_1925),
.B(n_1921),
.C(n_1870),
.Y(n_1945)
);

OAI21xp33_ASAP7_75t_L g1946 ( 
.A1(n_1928),
.A2(n_1921),
.B(n_1841),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_L g1947 ( 
.A(n_1933),
.B(n_1833),
.Y(n_1947)
);

AOI221xp5_ASAP7_75t_L g1948 ( 
.A1(n_1935),
.A2(n_1635),
.B1(n_1643),
.B2(n_1664),
.C(n_1656),
.Y(n_1948)
);

AOI211xp5_ASAP7_75t_SL g1949 ( 
.A1(n_1937),
.A2(n_1821),
.B(n_1836),
.C(n_1805),
.Y(n_1949)
);

AOI21xp33_ASAP7_75t_SL g1950 ( 
.A1(n_1928),
.A2(n_1805),
.B(n_1824),
.Y(n_1950)
);

INVx1_ASAP7_75t_SL g1951 ( 
.A(n_1944),
.Y(n_1951)
);

INVx5_ASAP7_75t_L g1952 ( 
.A(n_1943),
.Y(n_1952)
);

AOI22xp33_ASAP7_75t_SL g1953 ( 
.A1(n_1947),
.A2(n_1762),
.B1(n_1635),
.B2(n_1664),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1946),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1941),
.Y(n_1955)
);

INVx1_ASAP7_75t_SL g1956 ( 
.A(n_1945),
.Y(n_1956)
);

AOI222xp33_ASAP7_75t_L g1957 ( 
.A1(n_1940),
.A2(n_1643),
.B1(n_1714),
.B2(n_1673),
.C1(n_1656),
.C2(n_1664),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1951),
.B(n_1805),
.Y(n_1958)
);

NAND4xp25_ASAP7_75t_SL g1959 ( 
.A(n_1956),
.B(n_1950),
.C(n_1942),
.D(n_1949),
.Y(n_1959)
);

A2O1A1Ixp33_ASAP7_75t_L g1960 ( 
.A1(n_1952),
.A2(n_1948),
.B(n_1829),
.C(n_1668),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1952),
.A2(n_1829),
.B(n_1800),
.Y(n_1961)
);

NOR4xp75_ASAP7_75t_SL g1962 ( 
.A(n_1954),
.B(n_1743),
.C(n_1758),
.D(n_1761),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1955),
.Y(n_1963)
);

OAI221xp5_ASAP7_75t_L g1964 ( 
.A1(n_1961),
.A2(n_1957),
.B1(n_1953),
.B2(n_1800),
.C(n_1779),
.Y(n_1964)
);

NAND3xp33_ASAP7_75t_L g1965 ( 
.A(n_1963),
.B(n_1799),
.C(n_1779),
.Y(n_1965)
);

NOR4xp25_ASAP7_75t_L g1966 ( 
.A(n_1959),
.B(n_1799),
.C(n_1783),
.D(n_1789),
.Y(n_1966)
);

AO221x1_ASAP7_75t_L g1967 ( 
.A1(n_1962),
.A2(n_1783),
.B1(n_1789),
.B2(n_1785),
.C(n_1781),
.Y(n_1967)
);

NAND3xp33_ASAP7_75t_L g1968 ( 
.A(n_1958),
.B(n_1785),
.C(n_1781),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1965),
.Y(n_1969)
);

CKINVDCx12_ASAP7_75t_R g1970 ( 
.A(n_1966),
.Y(n_1970)
);

CKINVDCx20_ASAP7_75t_R g1971 ( 
.A(n_1968),
.Y(n_1971)
);

AOI22xp5_ASAP7_75t_SL g1972 ( 
.A1(n_1971),
.A2(n_1967),
.B1(n_1960),
.B2(n_1964),
.Y(n_1972)
);

OAI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1972),
.A2(n_1969),
.B1(n_1970),
.B2(n_1735),
.Y(n_1973)
);

BUFx2_ASAP7_75t_L g1974 ( 
.A(n_1973),
.Y(n_1974)
);

CKINVDCx20_ASAP7_75t_R g1975 ( 
.A(n_1973),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1974),
.B(n_1969),
.Y(n_1976)
);

INVx1_ASAP7_75t_SL g1977 ( 
.A(n_1975),
.Y(n_1977)
);

AOI222xp33_ASAP7_75t_L g1978 ( 
.A1(n_1977),
.A2(n_1741),
.B1(n_1643),
.B2(n_1753),
.C1(n_1744),
.C2(n_1747),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1976),
.Y(n_1979)
);

AOI322xp5_ASAP7_75t_L g1980 ( 
.A1(n_1979),
.A2(n_1741),
.A3(n_1744),
.B1(n_1747),
.B2(n_1736),
.C1(n_1757),
.C2(n_1760),
.Y(n_1980)
);

OAI221xp5_ASAP7_75t_R g1981 ( 
.A1(n_1980),
.A2(n_1978),
.B1(n_1797),
.B2(n_1747),
.C(n_1744),
.Y(n_1981)
);

AOI211xp5_ASAP7_75t_L g1982 ( 
.A1(n_1981),
.A2(n_1744),
.B(n_1747),
.C(n_1741),
.Y(n_1982)
);


endmodule