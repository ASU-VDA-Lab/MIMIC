module fake_jpeg_25291_n_62 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_62);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_62;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_44;
wire n_36;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx12_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_26),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_42),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_14),
.B1(n_24),
.B2(n_23),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_40),
.B1(n_35),
.B2(n_13),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_12),
.B1(n_22),
.B2(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_46),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_35),
.B1(n_30),
.B2(n_28),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_5),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_49)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_52),
.Y(n_54)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_51),
.B(n_48),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_55),
.A2(n_47),
.B1(n_53),
.B2(n_45),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_54),
.B(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

NOR3xp33_ASAP7_75t_SL g59 ( 
.A(n_58),
.B(n_53),
.C(n_9),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_6),
.Y(n_60)
);

AOI31xp33_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_15),
.A3(n_16),
.B(n_17),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_27),
.Y(n_62)
);


endmodule