module fake_jpeg_598_n_201 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_201);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_17),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_16),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_12),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_18),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_49),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_66),
.C(n_55),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_63),
.B1(n_53),
.B2(n_65),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_51),
.B1(n_68),
.B2(n_54),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_88),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_74),
.A2(n_63),
.B1(n_65),
.B2(n_70),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_92),
.B1(n_68),
.B2(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_51),
.B1(n_68),
.B2(n_67),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_67),
.B1(n_71),
.B2(n_69),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_102),
.B1(n_80),
.B2(n_57),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_104),
.Y(n_110)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_54),
.B1(n_58),
.B2(n_56),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_81),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_108),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_58),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_72),
.B1(n_64),
.B2(n_62),
.Y(n_109)
);

AO22x1_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_99),
.B1(n_96),
.B2(n_94),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_108),
.A2(n_90),
.B1(n_83),
.B2(n_52),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_128),
.B1(n_94),
.B2(n_6),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_109),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_117),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_46),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_9),
.C(n_10),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_123),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_1),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_129),
.Y(n_138)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_95),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_134),
.B1(n_139),
.B2(n_13),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_120),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_133),
.B(n_149),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_4),
.B(n_7),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_150),
.B(n_45),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_8),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_137),
.C(n_143),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_24),
.B1(n_44),
.B2(n_43),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_148),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_21),
.C(n_42),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_110),
.A2(n_31),
.B(n_41),
.C(n_40),
.D(n_33),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_119),
.B1(n_129),
.B2(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_153),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_146),
.A2(n_129),
.B1(n_12),
.B2(n_13),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_155),
.B(n_156),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_28),
.A3(n_27),
.B1(n_22),
.B2(n_29),
.C1(n_16),
.C2(n_17),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_11),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_158),
.B(n_160),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_147),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_131),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_163),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_136),
.B(n_14),
.Y(n_165)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_140),
.B(n_14),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_148),
.C(n_138),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_175),
.C(n_151),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_134),
.B(n_150),
.C(n_145),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_151),
.B(n_153),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_143),
.C(n_18),
.Y(n_175)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_167),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_186),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_173),
.B(n_178),
.Y(n_187)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_183),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_177),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_185),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_161),
.C(n_154),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_170),
.A2(n_161),
.B1(n_162),
.B2(n_155),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_185),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_180),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_192),
.B(n_193),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_R g194 ( 
.A(n_190),
.B(n_184),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_191),
.B(n_189),
.Y(n_196)
);

AO221x1_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_194),
.B1(n_172),
.B2(n_187),
.C(n_175),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_188),
.C(n_174),
.Y(n_198)
);

A2O1A1O1Ixp25_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_178),
.B(n_19),
.C(n_20),
.D(n_15),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_15),
.B(n_19),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_20),
.Y(n_201)
);


endmodule