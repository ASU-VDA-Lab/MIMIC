module fake_jpeg_26372_n_290 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx11_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_23),
.A2(n_0),
.B(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_29),
.B1(n_22),
.B2(n_34),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_48),
.A2(n_60),
.B1(n_68),
.B2(n_70),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_22),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_22),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_29),
.B1(n_31),
.B2(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_59),
.Y(n_80)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_29),
.B1(n_18),
.B2(n_32),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_57),
.A2(n_71),
.B1(n_0),
.B2(n_1),
.Y(n_109)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_18),
.B1(n_21),
.B2(n_35),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_31),
.B1(n_27),
.B2(n_21),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_67),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_35),
.B1(n_24),
.B2(n_32),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_24),
.B1(n_32),
.B2(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_45),
.B1(n_18),
.B2(n_24),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_38),
.B1(n_20),
.B2(n_26),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_25),
.B1(n_33),
.B2(n_28),
.Y(n_71)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_43),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_28),
.B1(n_33),
.B2(n_25),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_20),
.B(n_30),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_74),
.A2(n_84),
.B(n_94),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_82),
.Y(n_124)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_37),
.C(n_26),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_88),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_73),
.B(n_37),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_83),
.B(n_93),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_33),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_86),
.B(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_36),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_70),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_66),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_33),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_50),
.A2(n_28),
.B1(n_25),
.B2(n_11),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_96),
.A2(n_110),
.B1(n_111),
.B2(n_72),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_61),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_100),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_36),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_65),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_28),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_53),
.A2(n_36),
.B(n_9),
.C(n_11),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_103),
.B(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_25),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_104),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_57),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_8),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_72),
.B(n_8),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_108),
.A2(n_17),
.B1(n_9),
.B2(n_12),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_72),
.B1(n_69),
.B2(n_62),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_71),
.B(n_0),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_1),
.B(n_2),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_119),
.A2(n_133),
.B1(n_139),
.B2(n_92),
.Y(n_160)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_130),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_SL g168 ( 
.A(n_123),
.B(n_137),
.C(n_12),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_13),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_117),
.B(n_124),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_99),
.A2(n_56),
.B1(n_69),
.B2(n_62),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_56),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_132),
.B1(n_108),
.B2(n_83),
.Y(n_145)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_87),
.B1(n_77),
.B2(n_82),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_90),
.B1(n_109),
.B2(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_140),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_94),
.A2(n_84),
.B1(n_87),
.B2(n_76),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_78),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_79),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_143),
.A2(n_161),
.B(n_168),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_152),
.B1(n_128),
.B2(n_116),
.Y(n_172)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_135),
.A2(n_111),
.B(n_93),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_112),
.B(n_16),
.Y(n_181)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_166),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_125),
.B(n_86),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_150),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_121),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_80),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_153),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_110),
.B1(n_105),
.B2(n_103),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_102),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_80),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_107),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_130),
.B(n_92),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_157),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_92),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_158),
.B(n_164),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_98),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_163),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_162),
.B1(n_129),
.B2(n_156),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_2),
.B(n_3),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_133),
.A2(n_91),
.B1(n_89),
.B2(n_98),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_91),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_89),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_165),
.B(n_170),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_98),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_116),
.A2(n_89),
.B1(n_78),
.B2(n_13),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_85),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_172),
.A2(n_175),
.B1(n_179),
.B2(n_166),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_173),
.A2(n_182),
.B1(n_191),
.B2(n_148),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_152),
.A2(n_119),
.B1(n_126),
.B2(n_138),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_154),
.A2(n_120),
.B1(n_112),
.B2(n_134),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_181),
.A2(n_197),
.B(n_158),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_140),
.B1(n_122),
.B2(n_134),
.Y(n_182)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_113),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_142),
.B(n_113),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_144),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_141),
.B1(n_114),
.B2(n_85),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_146),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_193),
.B(n_195),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_149),
.B(n_85),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_196),
.B(n_144),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_170),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_176),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_206),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_185),
.B(n_155),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_207),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_175),
.B1(n_192),
.B2(n_186),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_216),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_151),
.B(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_147),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_198),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_214),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_153),
.C(n_150),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_174),
.C(n_180),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_188),
.A2(n_171),
.B(n_145),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_218),
.B(n_195),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_157),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_172),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_213),
.A2(n_217),
.B1(n_220),
.B2(n_196),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_178),
.B(n_161),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_114),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_215),
.Y(n_235)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_222),
.C(n_229),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_187),
.C(n_193),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_233),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_226),
.B(n_202),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_184),
.B(n_198),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_178),
.C(n_177),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_174),
.Y(n_233)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_234),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_203),
.A2(n_173),
.B1(n_182),
.B2(n_177),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_197),
.B1(n_216),
.B2(n_220),
.Y(n_247)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_184),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_218),
.C(n_209),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_248),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_227),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_246),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_233),
.B(n_217),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_247),
.A2(n_249),
.B1(n_204),
.B2(n_208),
.Y(n_257)
);

NAND2x1_ASAP7_75t_SL g249 ( 
.A(n_224),
.B(n_186),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_211),
.C(n_197),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_250),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_235),
.Y(n_253)
);

NOR3xp33_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_243),
.C(n_240),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_252),
.A2(n_234),
.B1(n_225),
.B2(n_226),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_255),
.B(n_260),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_261),
.B1(n_223),
.B2(n_258),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_232),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_247),
.A2(n_236),
.B1(n_229),
.B2(n_211),
.Y(n_261)
);

NOR2x1_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_231),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_239),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_264),
.A2(n_244),
.A3(n_253),
.B1(n_248),
.B2(n_261),
.C1(n_262),
.C2(n_245),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_272),
.Y(n_273)
);

AOI21x1_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_249),
.B(n_252),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_269),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_268),
.A2(n_270),
.B1(n_191),
.B2(n_164),
.Y(n_277)
);

OAI221xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_251),
.B1(n_239),
.B2(n_176),
.C(n_221),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_271),
.A2(n_241),
.B1(n_250),
.B2(n_258),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_241),
.C(n_242),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_277),
.Y(n_280)
);

NOR2x1_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_257),
.Y(n_276)
);

AOI311xp33_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_238),
.A3(n_230),
.B(n_254),
.C(n_201),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_272),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_278),
.A2(n_275),
.B(n_276),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_L g283 ( 
.A1(n_279),
.A2(n_281),
.A3(n_274),
.B1(n_278),
.B2(n_230),
.C1(n_201),
.C2(n_148),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_169),
.C(n_7),
.Y(n_285)
);

AOI322xp5_ASAP7_75t_L g287 ( 
.A1(n_283),
.A2(n_284),
.A3(n_285),
.B1(n_169),
.B2(n_13),
.C1(n_6),
.C2(n_14),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_274),
.A3(n_201),
.B1(n_169),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_283),
.A2(n_169),
.B(n_7),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_287),
.B(n_14),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_14),
.Y(n_289)
);

NOR3xp33_ASAP7_75t_L g290 ( 
.A(n_289),
.B(n_15),
.C(n_3),
.Y(n_290)
);


endmodule