module fake_netlist_5_879_n_1724 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1724);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1724;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx2_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_41),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_122),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_10),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_6),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_0),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_116),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_92),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_97),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_81),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_82),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_73),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_62),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_84),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_68),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_83),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_123),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_6),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_31),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_39),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_127),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_76),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_135),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_55),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_99),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_0),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_104),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_74),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_50),
.Y(n_187)
);

CKINVDCx6p67_ASAP7_75t_R g188 ( 
.A(n_152),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_142),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_67),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_77),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_42),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_42),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_19),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_52),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_38),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_138),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_91),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_37),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_90),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_32),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_29),
.Y(n_202)
);

INVxp67_ASAP7_75t_SL g203 ( 
.A(n_121),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_33),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_126),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_26),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_45),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_19),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_79),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_71),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_48),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_53),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_56),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_57),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_7),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_149),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_21),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_141),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_16),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_1),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_31),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_93),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_28),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_59),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_61),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_41),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_151),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_49),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_9),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_9),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_154),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_69),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_100),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g234 ( 
.A(n_18),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_33),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_133),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_89),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_113),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_34),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_16),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_70),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_107),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_43),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_95),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_13),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_98),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_26),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_29),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_17),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_21),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_18),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_128),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_80),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_43),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_36),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_88),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_63),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_143),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_1),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_27),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_101),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_118),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_72),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_111),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_94),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_34),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_32),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_5),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_139),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_87),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_145),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_54),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_11),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_22),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_125),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_58),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_45),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_108),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_86),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_112),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_114),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_39),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_131),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_144),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_65),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_64),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_3),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_60),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_75),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_22),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_115),
.Y(n_291)
);

BUFx2_ASAP7_75t_SL g292 ( 
.A(n_13),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_36),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_66),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_85),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_37),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_7),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_10),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_132),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_119),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_40),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_51),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_96),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_15),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_28),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_20),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_46),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_30),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_109),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_226),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_234),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_257),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_234),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_234),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_156),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_202),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_234),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_234),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_176),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_254),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_165),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_179),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_281),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_234),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_234),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_234),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_180),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_181),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g329 ( 
.A(n_178),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_268),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_221),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_268),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

BUFx10_ASAP7_75t_L g334 ( 
.A(n_269),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_268),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_268),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_257),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_186),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_230),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_158),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_230),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_198),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_158),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_184),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_257),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_248),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_182),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_210),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g349 ( 
.A(n_160),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_248),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_183),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_266),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_160),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_266),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_184),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_259),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_194),
.Y(n_357)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_188),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_259),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_185),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_217),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_229),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_189),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_239),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_190),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_243),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_245),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_195),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_209),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_249),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_211),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_166),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_274),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_282),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_298),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_212),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_155),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_155),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_286),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_273),
.Y(n_380)
);

INVxp33_ASAP7_75t_L g381 ( 
.A(n_167),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_172),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_222),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_191),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_311),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_330),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_315),
.B(n_269),
.Y(n_388)
);

INVxp33_ASAP7_75t_SL g389 ( 
.A(n_319),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_311),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_313),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

NOR2x1_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_191),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_332),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_314),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_332),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_314),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_333),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_333),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_335),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_331),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_335),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_336),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_315),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_315),
.B(n_289),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_372),
.B(n_382),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_317),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_317),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_318),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_344),
.B(n_286),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_318),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_324),
.B(n_289),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_324),
.B(n_157),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_325),
.B(n_157),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_350),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_325),
.B(n_159),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_350),
.Y(n_418)
);

INVx6_ASAP7_75t_L g419 ( 
.A(n_334),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_326),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_326),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_377),
.B(n_261),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_357),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_378),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_357),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_378),
.B(n_261),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_R g427 ( 
.A(n_358),
.B(n_365),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_362),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_384),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_362),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_384),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_375),
.B(n_294),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_322),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_361),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_355),
.B(n_286),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_355),
.B(n_188),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_361),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_321),
.B(n_192),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_364),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_356),
.B(n_159),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_364),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_339),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_366),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_356),
.B(n_163),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_366),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_380),
.Y(n_447)
);

NOR2x1_ASAP7_75t_L g448 ( 
.A(n_312),
.B(n_294),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_327),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_367),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_339),
.A2(n_187),
.B(n_175),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_359),
.B(n_163),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_341),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_340),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_367),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_439),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_421),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_408),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_404),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_445),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_390),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_421),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_389),
.B(n_345),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_390),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_436),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_436),
.B(n_359),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_390),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_391),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_391),
.Y(n_469)
);

OAI22xp33_ASAP7_75t_L g470 ( 
.A1(n_407),
.A2(n_345),
.B1(n_379),
.B2(n_381),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_391),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_414),
.A2(n_310),
.B1(n_323),
.B2(n_320),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_392),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_404),
.B(n_328),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_392),
.Y(n_475)
);

OR2x6_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_292),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_392),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_408),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_434),
.B(n_379),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_395),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_404),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_401),
.Y(n_482)
);

NOR2x1p5_ASAP7_75t_L g483 ( 
.A(n_449),
.B(n_312),
.Y(n_483)
);

BUFx10_ASAP7_75t_L g484 ( 
.A(n_419),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_395),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_395),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_397),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_407),
.B(n_347),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_L g489 ( 
.A(n_414),
.B(n_351),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_397),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_SL g492 ( 
.A(n_447),
.B(n_383),
.Y(n_492)
);

NAND3xp33_ASAP7_75t_L g493 ( 
.A(n_415),
.B(n_373),
.C(n_370),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_410),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_408),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_415),
.A2(n_310),
.B1(n_349),
.B2(n_353),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_411),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_417),
.B(n_360),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_410),
.Y(n_499)
);

XOR2x2_ASAP7_75t_L g500 ( 
.A(n_439),
.B(n_343),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_410),
.Y(n_501)
);

OAI22x1_ASAP7_75t_L g502 ( 
.A1(n_454),
.A2(n_174),
.B1(n_162),
.B2(n_161),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_408),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_412),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_412),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_427),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_412),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_420),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_401),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_408),
.Y(n_510)
);

AO21x2_ASAP7_75t_L g511 ( 
.A1(n_451),
.A2(n_205),
.B(n_197),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_411),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_417),
.B(n_363),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_420),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_447),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_454),
.Y(n_517)
);

OR2x6_ASAP7_75t_L g518 ( 
.A(n_448),
.B(n_213),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_419),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_443),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_437),
.Y(n_521)
);

OA22x2_ASAP7_75t_L g522 ( 
.A1(n_441),
.A2(n_374),
.B1(n_373),
.B2(n_370),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_388),
.B(n_376),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_437),
.B(n_316),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_443),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_443),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_443),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_388),
.B(n_334),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_419),
.B(n_368),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_419),
.B(n_369),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_385),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_388),
.B(n_334),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_443),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_443),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_405),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_385),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_408),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_385),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_387),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_441),
.B(n_316),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_387),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_409),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_452),
.B(n_214),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_394),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_394),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_385),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_452),
.B(n_371),
.Y(n_547)
);

INVx8_ASAP7_75t_L g548 ( 
.A(n_405),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_396),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_405),
.B(n_334),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_405),
.B(n_203),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_409),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_409),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_396),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_398),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_398),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_SL g557 ( 
.A(n_413),
.B(n_235),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_400),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_432),
.B(n_337),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_400),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_403),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_403),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_429),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_409),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_409),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_409),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_419),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_432),
.B(n_337),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_386),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_432),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_432),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_435),
.B(n_164),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_SL g573 ( 
.A1(n_435),
.A2(n_260),
.B1(n_267),
.B2(n_308),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_386),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_413),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_438),
.B(n_164),
.Y(n_576)
);

INVxp33_ASAP7_75t_L g577 ( 
.A(n_438),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_440),
.B(n_168),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_422),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_433),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_433),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_440),
.B(n_168),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_442),
.B(n_169),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_433),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_433),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_386),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_442),
.B(n_329),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_429),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_444),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_433),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_429),
.Y(n_591)
);

BUFx4f_ASAP7_75t_L g592 ( 
.A(n_433),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_444),
.B(n_169),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_446),
.B(n_338),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g595 ( 
.A(n_386),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_386),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_386),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_431),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_446),
.B(n_170),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_431),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_422),
.A2(n_263),
.B1(n_200),
.B2(n_374),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_431),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_422),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_422),
.A2(n_200),
.B1(n_263),
.B2(n_302),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_424),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_488),
.B(n_426),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_571),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_570),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_497),
.A2(n_342),
.B1(n_348),
.B2(n_228),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_535),
.B(n_426),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_535),
.B(n_575),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_575),
.B(n_426),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_546),
.Y(n_613)
);

OAI22xp33_ASAP7_75t_L g614 ( 
.A1(n_497),
.A2(n_232),
.B1(n_216),
.B2(n_307),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_539),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_459),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_512),
.B(n_170),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_551),
.B(n_498),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_539),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_541),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_603),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_551),
.B(n_426),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_587),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_543),
.A2(n_451),
.B1(n_263),
.B2(n_200),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_506),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_551),
.B(n_424),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_R g627 ( 
.A(n_506),
.B(n_171),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_541),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_551),
.B(n_424),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_512),
.B(n_171),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_603),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_513),
.B(n_424),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_521),
.B(n_200),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_589),
.B(n_450),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_548),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_543),
.A2(n_451),
.B1(n_200),
.B2(n_263),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_521),
.B(n_460),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_544),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_517),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_544),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_460),
.B(n_263),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_465),
.B(n_424),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_482),
.B(n_455),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_579),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_465),
.B(n_589),
.Y(n_645)
);

NOR2x1_ASAP7_75t_L g646 ( 
.A(n_529),
.B(n_530),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_579),
.B(n_424),
.Y(n_647)
);

NOR2xp67_ASAP7_75t_L g648 ( 
.A(n_493),
.B(n_450),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_554),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_519),
.B(n_173),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_554),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_577),
.B(n_173),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_548),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_545),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_548),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_457),
.B(n_399),
.Y(n_656)
);

O2A1O1Ixp5_ASAP7_75t_L g657 ( 
.A1(n_457),
.A2(n_224),
.B(n_227),
.C(n_218),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_545),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_555),
.Y(n_659)
);

NOR3xp33_ASAP7_75t_L g660 ( 
.A(n_470),
.B(n_455),
.C(n_240),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_549),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_549),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_459),
.B(n_481),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_519),
.B(n_303),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_523),
.B(n_303),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_466),
.B(n_273),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_555),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_462),
.B(n_399),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_528),
.B(n_225),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_548),
.B(n_399),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_560),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_548),
.B(n_466),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_517),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_556),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_556),
.B(n_399),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_558),
.B(n_399),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_558),
.B(n_402),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_543),
.A2(n_241),
.B1(n_252),
.B2(n_246),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_561),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_561),
.B(n_531),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_531),
.B(n_536),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_540),
.B(n_177),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_546),
.B(n_276),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_536),
.B(n_402),
.Y(n_684)
);

INVxp67_ASAP7_75t_SL g685 ( 
.A(n_546),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_547),
.B(n_193),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_560),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_538),
.B(n_402),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_524),
.B(n_196),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_543),
.A2(n_300),
.B1(n_283),
.B2(n_393),
.Y(n_690)
);

NAND3xp33_ASAP7_75t_L g691 ( 
.A(n_472),
.B(n_255),
.C(n_251),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_562),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_538),
.B(n_402),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_459),
.B(n_423),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_532),
.B(n_231),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_543),
.B(n_402),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_550),
.B(n_481),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_482),
.B(n_273),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_481),
.B(n_567),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_496),
.B(n_233),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_594),
.B(n_474),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_559),
.B(n_423),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_458),
.Y(n_703)
);

A2O1A1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_493),
.A2(n_393),
.B(n_453),
.C(n_428),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_567),
.B(n_402),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_516),
.B(n_236),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_553),
.B(n_406),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_562),
.B(n_406),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_574),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_563),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_509),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_563),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_489),
.B(n_406),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_516),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_511),
.A2(n_162),
.B1(n_306),
.B2(n_305),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_564),
.B(n_406),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_564),
.B(n_406),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_565),
.B(n_406),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_568),
.B(n_425),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_588),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_565),
.B(n_566),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_566),
.B(n_453),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_588),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_458),
.B(n_478),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_591),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_573),
.B(n_297),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_458),
.B(n_453),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_476),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_572),
.B(n_199),
.Y(n_729)
);

AO221x1_ASAP7_75t_L g730 ( 
.A1(n_502),
.A2(n_537),
.B1(n_503),
.B2(n_510),
.C(n_495),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_576),
.B(n_201),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_478),
.B(n_416),
.Y(n_732)
);

NOR2xp67_ASAP7_75t_L g733 ( 
.A(n_463),
.B(n_416),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_478),
.B(n_418),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_578),
.B(n_204),
.Y(n_735)
);

OAI22xp33_ASAP7_75t_SL g736 ( 
.A1(n_476),
.A2(n_301),
.B1(n_174),
.B2(n_304),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_591),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_557),
.B(n_237),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_484),
.B(n_479),
.Y(n_739)
);

INVxp67_ASAP7_75t_SL g740 ( 
.A(n_495),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_495),
.B(n_503),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_598),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_483),
.B(n_297),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_484),
.B(n_238),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_492),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_503),
.B(n_510),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_484),
.B(n_242),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_598),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_510),
.B(n_418),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_456),
.B(n_301),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_476),
.Y(n_751)
);

OAI22xp33_ASAP7_75t_L g752 ( 
.A1(n_476),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_537),
.B(n_425),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_483),
.B(n_297),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_537),
.B(n_428),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_582),
.B(n_206),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_600),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_542),
.B(n_552),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_600),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_583),
.B(n_207),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_602),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_542),
.B(n_430),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_542),
.B(n_430),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_L g764 ( 
.A(n_502),
.B(n_244),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_520),
.B(n_253),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_593),
.B(n_208),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_599),
.B(n_215),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_552),
.B(n_256),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_602),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_552),
.B(n_258),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_476),
.B(n_219),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_518),
.A2(n_280),
.B1(n_262),
.B2(n_264),
.Y(n_772)
);

AND2x2_ASAP7_75t_SL g773 ( 
.A(n_604),
.B(n_341),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_518),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_618),
.B(n_464),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_634),
.B(n_601),
.Y(n_776)
);

BUFx4f_ASAP7_75t_SL g777 ( 
.A(n_711),
.Y(n_777)
);

INVx5_ASAP7_75t_L g778 ( 
.A(n_653),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_615),
.Y(n_779)
);

INVx5_ASAP7_75t_L g780 ( 
.A(n_653),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_608),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_623),
.B(n_518),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_607),
.B(n_518),
.Y(n_783)
);

INVx5_ASAP7_75t_L g784 ( 
.A(n_653),
.Y(n_784)
);

INVx8_ASAP7_75t_L g785 ( 
.A(n_663),
.Y(n_785)
);

INVxp67_ASAP7_75t_SL g786 ( 
.A(n_613),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_646),
.B(n_592),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_730),
.A2(n_518),
.B1(n_511),
.B2(n_467),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_643),
.Y(n_789)
);

AND3x1_ASAP7_75t_L g790 ( 
.A(n_726),
.B(n_500),
.C(n_354),
.Y(n_790)
);

AOI21xp33_ASAP7_75t_L g791 ( 
.A1(n_690),
.A2(n_715),
.B(n_686),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_701),
.B(n_595),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_715),
.A2(n_511),
.B1(n_490),
.B2(n_464),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_606),
.B(n_467),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_663),
.B(n_616),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_642),
.B(n_649),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_613),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_625),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_619),
.Y(n_799)
);

AO22x1_ASAP7_75t_L g800 ( 
.A1(n_686),
.A2(n_290),
.B1(n_223),
.B2(n_247),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_651),
.B(n_473),
.Y(n_801)
);

BUFx12f_ASAP7_75t_L g802 ( 
.A(n_714),
.Y(n_802)
);

OAI21xp5_ASAP7_75t_L g803 ( 
.A1(n_624),
.A2(n_508),
.B(n_473),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_621),
.Y(n_804)
);

BUFx8_ASAP7_75t_L g805 ( 
.A(n_698),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_659),
.B(n_475),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_667),
.B(n_475),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_666),
.B(n_522),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_639),
.B(n_522),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_673),
.B(n_522),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_750),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_631),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_620),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_616),
.B(n_520),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_645),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_652),
.B(n_500),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_628),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_613),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_652),
.B(n_611),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_637),
.B(n_728),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_704),
.A2(n_505),
.B(n_490),
.C(n_491),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_R g822 ( 
.A(n_751),
.B(n_265),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_628),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_674),
.B(n_485),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_613),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_709),
.Y(n_826)
);

BUFx4f_ASAP7_75t_L g827 ( 
.A(n_743),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_638),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_612),
.B(n_592),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_638),
.Y(n_830)
);

INVx5_ASAP7_75t_L g831 ( 
.A(n_653),
.Y(n_831)
);

NAND3xp33_ASAP7_75t_SL g832 ( 
.A(n_660),
.B(n_293),
.C(n_250),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_672),
.A2(n_644),
.B1(n_697),
.B2(n_774),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_697),
.A2(n_648),
.B1(n_771),
.B2(n_637),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_SL g835 ( 
.A1(n_729),
.A2(n_605),
.B(n_525),
.C(n_533),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_771),
.B(n_270),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_640),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_640),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_624),
.A2(n_220),
.B1(n_277),
.B2(n_287),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_694),
.B(n_702),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_702),
.B(n_271),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_682),
.B(n_346),
.Y(n_842)
);

AND2x4_ASAP7_75t_L g843 ( 
.A(n_694),
.B(n_525),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_682),
.B(n_346),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_679),
.B(n_485),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_654),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_754),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_719),
.B(n_526),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_609),
.Y(n_849)
);

BUFx4f_ASAP7_75t_L g850 ( 
.A(n_719),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_680),
.B(n_491),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_654),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_689),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_733),
.B(n_272),
.Y(n_854)
);

NOR2xp67_ASAP7_75t_L g855 ( 
.A(n_745),
.B(n_526),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_729),
.B(n_275),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_709),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_709),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_706),
.B(n_296),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_617),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_658),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_658),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_630),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_661),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_709),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_661),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_662),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_662),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_671),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_671),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_692),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_690),
.A2(n_508),
.B1(n_499),
.B2(n_501),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_632),
.B(n_687),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_681),
.B(n_499),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_731),
.B(n_278),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_622),
.B(n_501),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_700),
.B(n_689),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_636),
.A2(n_515),
.B1(n_504),
.B2(n_505),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_731),
.B(n_279),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_735),
.B(n_284),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_710),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_735),
.B(n_352),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_720),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_725),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_696),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_685),
.B(n_504),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_756),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_737),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_756),
.B(n_285),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_737),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_773),
.B(n_748),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_748),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_627),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_773),
.B(n_515),
.Y(n_894)
);

INVx4_ASAP7_75t_L g895 ( 
.A(n_635),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_678),
.Y(n_896)
);

BUFx5_ASAP7_75t_L g897 ( 
.A(n_712),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_760),
.B(n_288),
.Y(n_898)
);

O2A1O1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_641),
.A2(n_487),
.B(n_461),
.C(n_486),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_627),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_760),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_695),
.A2(n_585),
.B1(n_580),
.B2(n_581),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_764),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_766),
.Y(n_904)
);

OR2x6_ASAP7_75t_L g905 ( 
.A(n_739),
.B(n_352),
.Y(n_905)
);

NOR3xp33_ASAP7_75t_SL g906 ( 
.A(n_752),
.B(n_291),
.C(n_295),
.Y(n_906)
);

OAI21xp33_ASAP7_75t_SL g907 ( 
.A1(n_636),
.A2(n_581),
.B(n_584),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_767),
.B(n_299),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_759),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_759),
.B(n_769),
.Y(n_910)
);

INVx5_ASAP7_75t_L g911 ( 
.A(n_635),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_769),
.B(n_514),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_699),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_753),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_610),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_772),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_767),
.Y(n_917)
);

O2A1O1Ixp5_ASAP7_75t_L g918 ( 
.A1(n_641),
.A2(n_633),
.B(n_683),
.C(n_657),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_691),
.B(n_354),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_SL g920 ( 
.A(n_655),
.B(n_309),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_723),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_755),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_762),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_763),
.Y(n_924)
);

OR2x6_ASAP7_75t_L g925 ( 
.A(n_738),
.B(n_605),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_626),
.B(n_629),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_742),
.B(n_514),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_757),
.B(n_461),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_665),
.B(n_527),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_761),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_721),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_732),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_734),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_749),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_683),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_722),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_633),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_695),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_703),
.B(n_468),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_SL g940 ( 
.A1(n_736),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_740),
.B(n_468),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_650),
.B(n_584),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_656),
.B(n_469),
.Y(n_943)
);

NOR2xp67_ASAP7_75t_L g944 ( 
.A(n_664),
.B(n_533),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_765),
.A2(n_590),
.B1(n_585),
.B2(n_527),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_768),
.Y(n_946)
);

AND2x6_ASAP7_75t_L g947 ( 
.A(n_724),
.B(n_534),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_669),
.B(n_471),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_668),
.B(n_507),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_765),
.B(n_471),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_675),
.B(n_477),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_676),
.B(n_477),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_677),
.B(n_480),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_614),
.B(n_596),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_926),
.A2(n_670),
.B(n_713),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_777),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_887),
.B(n_770),
.Y(n_957)
);

INVx5_ASAP7_75t_L g958 ( 
.A(n_826),
.Y(n_958)
);

BUFx12f_ASAP7_75t_L g959 ( 
.A(n_802),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_819),
.B(n_747),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_791),
.A2(n_747),
.B(n_647),
.C(n_758),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_888),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_789),
.B(n_708),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_781),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_SL g965 ( 
.A(n_798),
.B(n_741),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_853),
.B(n_727),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_888),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_917),
.B(n_744),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_796),
.B(n_746),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_796),
.B(n_684),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_805),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_SL g972 ( 
.A(n_791),
.B(n_688),
.Y(n_972)
);

NOR2x1_ASAP7_75t_L g973 ( 
.A(n_901),
.B(n_693),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_877),
.A2(n_718),
.B(n_717),
.C(n_716),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_850),
.A2(n_705),
.B1(n_707),
.B2(n_480),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_826),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_825),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_926),
.A2(n_597),
.B(n_574),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_804),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_896),
.A2(n_839),
.B(n_875),
.C(n_856),
.Y(n_980)
);

BUFx2_ASAP7_75t_L g981 ( 
.A(n_811),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_808),
.B(n_936),
.Y(n_982)
);

NAND2xp33_ASAP7_75t_SL g983 ( 
.A(n_906),
.B(n_597),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_842),
.B(n_486),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_775),
.A2(n_597),
.B(n_574),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_844),
.B(n_494),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_816),
.B(n_487),
.Y(n_987)
);

CKINVDCx20_ASAP7_75t_R g988 ( 
.A(n_805),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_882),
.B(n_494),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_809),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_826),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_850),
.A2(n_793),
.B1(n_776),
.B2(n_891),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_891),
.A2(n_596),
.B1(n_569),
.B2(n_574),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_919),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_914),
.B(n_597),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_922),
.B(n_586),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_899),
.A2(n_586),
.B(n_47),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_923),
.B(n_586),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_783),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_839),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_879),
.A2(n_8),
.B(n_11),
.C(n_12),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_840),
.B(n_586),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_812),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_782),
.B(n_8),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_932),
.B(n_586),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_881),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_778),
.A2(n_586),
.B(n_105),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_858),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_894),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_894),
.A2(n_14),
.B1(n_17),
.B2(n_20),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_R g1011 ( 
.A(n_832),
.B(n_117),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_794),
.B(n_110),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_849),
.B(n_23),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_SL g1014 ( 
.A(n_832),
.B(n_23),
.C(n_24),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_840),
.B(n_120),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_827),
.B(n_124),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_827),
.B(n_106),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_778),
.A2(n_130),
.B(n_150),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_785),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_783),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_SL g1021 ( 
.A(n_893),
.B(n_78),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_795),
.B(n_153),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_880),
.A2(n_24),
.B(n_25),
.C(n_27),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_825),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_825),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_795),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_778),
.A2(n_136),
.B(n_146),
.Y(n_1027)
);

OAI21xp33_ASAP7_75t_SL g1028 ( 
.A1(n_803),
.A2(n_25),
.B(n_30),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_778),
.A2(n_784),
.B(n_780),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_820),
.B(n_137),
.Y(n_1030)
);

INVx8_ASAP7_75t_L g1031 ( 
.A(n_785),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_813),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_889),
.A2(n_35),
.B(n_38),
.C(n_40),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_815),
.B(n_35),
.Y(n_1034)
);

OAI21xp33_ASAP7_75t_L g1035 ( 
.A1(n_859),
.A2(n_44),
.B(n_140),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_SL g1036 ( 
.A1(n_790),
.A2(n_940),
.B1(n_916),
.B2(n_847),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_810),
.B(n_44),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_834),
.A2(n_148),
.B1(n_878),
.B2(n_794),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_858),
.Y(n_1039)
);

AOI21xp33_ASAP7_75t_L g1040 ( 
.A1(n_898),
.A2(n_908),
.B(n_938),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_779),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_858),
.Y(n_1042)
);

BUFx4f_ASAP7_75t_L g1043 ( 
.A(n_900),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_931),
.B(n_934),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_863),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_885),
.A2(n_935),
.B1(n_915),
.B2(n_931),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_830),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_860),
.B(n_915),
.Y(n_1048)
);

AOI21x1_ASAP7_75t_L g1049 ( 
.A1(n_829),
.A2(n_787),
.B(n_873),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_931),
.B(n_792),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_841),
.B(n_915),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_924),
.B(n_933),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_937),
.B(n_873),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_851),
.A2(n_937),
.B1(n_940),
.B2(n_803),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_865),
.Y(n_1055)
);

NAND2xp33_ASAP7_75t_SL g1056 ( 
.A(n_903),
.B(n_895),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_851),
.B(n_874),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_843),
.B(n_885),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_836),
.A2(n_854),
.B(n_954),
.C(n_806),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_885),
.B(n_911),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_837),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_874),
.B(n_876),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_797),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_905),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_780),
.A2(n_784),
.B(n_831),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_799),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_780),
.A2(n_784),
.B(n_831),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_911),
.B(n_833),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_876),
.B(n_801),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_905),
.Y(n_1070)
);

NAND2x1p5_ASAP7_75t_L g1071 ( 
.A(n_911),
.B(n_895),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_801),
.B(n_806),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_911),
.B(n_780),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_929),
.A2(n_942),
.B1(n_946),
.B2(n_848),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_822),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_872),
.A2(n_845),
.B1(n_807),
.B2(n_824),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_807),
.A2(n_845),
.B1(n_824),
.B2(n_788),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_784),
.B(n_831),
.Y(n_1078)
);

INVx4_ASAP7_75t_L g1079 ( 
.A(n_865),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_905),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_800),
.B(n_848),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_913),
.B(n_930),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_831),
.A2(n_886),
.B(n_939),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_865),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_929),
.A2(n_843),
.B1(n_913),
.B2(n_948),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_913),
.B(n_920),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_886),
.A2(n_941),
.B(n_939),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_855),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_930),
.B(n_866),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_921),
.A2(n_814),
.B1(n_950),
.B2(n_944),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_814),
.B(n_797),
.Y(n_1091)
);

AOI21xp33_ASAP7_75t_L g1092 ( 
.A1(n_980),
.A2(n_925),
.B(n_907),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_SL g1093 ( 
.A(n_956),
.B(n_920),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_964),
.Y(n_1094)
);

NAND3xp33_ASAP7_75t_SL g1095 ( 
.A(n_1013),
.B(n_918),
.C(n_902),
.Y(n_1095)
);

AOI211x1_ASAP7_75t_L g1096 ( 
.A1(n_1054),
.A2(n_982),
.B(n_1010),
.C(n_1009),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_1059),
.A2(n_821),
.B(n_945),
.C(n_846),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1057),
.B(n_953),
.Y(n_1098)
);

NAND2x1p5_ASAP7_75t_L g1099 ( 
.A(n_1019),
.B(n_857),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_955),
.A2(n_912),
.B(n_910),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_994),
.B(n_866),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_981),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1036),
.A2(n_864),
.B1(n_868),
.B2(n_871),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_979),
.Y(n_1104)
);

NOR2x1_ASAP7_75t_SL g1105 ( 
.A(n_1073),
.B(n_925),
.Y(n_1105)
);

NOR4xp25_ASAP7_75t_L g1106 ( 
.A(n_1000),
.B(n_861),
.C(n_838),
.D(n_862),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1057),
.A2(n_953),
.B(n_952),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1087),
.A2(n_951),
.B(n_949),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_985),
.A2(n_912),
.B(n_910),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_976),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_1091),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1003),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_987),
.B(n_870),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_R g1114 ( 
.A(n_1075),
.B(n_818),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_1045),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1049),
.A2(n_943),
.B(n_927),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1062),
.B(n_1053),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_990),
.B(n_869),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1062),
.B(n_943),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_999),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1069),
.B(n_786),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1032),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1038),
.A2(n_928),
.B(n_927),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1072),
.A2(n_835),
.B(n_857),
.Y(n_1124)
);

OR2x6_ASAP7_75t_L g1125 ( 
.A(n_1031),
.B(n_925),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1072),
.A2(n_928),
.B(n_866),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1069),
.B(n_817),
.Y(n_1127)
);

AOI31xp67_ASAP7_75t_L g1128 ( 
.A1(n_1068),
.A2(n_1012),
.A3(n_1086),
.B(n_957),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1034),
.B(n_823),
.Y(n_1129)
);

CKINVDCx6p67_ASAP7_75t_R g1130 ( 
.A(n_959),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_966),
.B(n_828),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_970),
.A2(n_890),
.B(n_909),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_970),
.A2(n_883),
.B(n_884),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_982),
.B(n_852),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1047),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1083),
.A2(n_892),
.B(n_867),
.Y(n_1136)
);

INVxp67_ASAP7_75t_SL g1137 ( 
.A(n_1044),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1038),
.A2(n_961),
.B(n_1077),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_993),
.A2(n_947),
.B(n_897),
.Y(n_1139)
);

AOI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1076),
.A2(n_947),
.B(n_897),
.Y(n_1140)
);

O2A1O1Ixp5_ASAP7_75t_SL g1141 ( 
.A1(n_1009),
.A2(n_897),
.B(n_947),
.C(n_1010),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1076),
.A2(n_897),
.B(n_947),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_993),
.A2(n_897),
.B(n_1029),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1061),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1065),
.A2(n_1067),
.B(n_975),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1006),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_975),
.A2(n_995),
.B(n_1012),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_1043),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1074),
.A2(n_1046),
.B1(n_1085),
.B2(n_1050),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_R g1150 ( 
.A(n_1056),
.B(n_1031),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1054),
.A2(n_960),
.B1(n_1077),
.B2(n_1090),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_1052),
.B(n_1020),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_1064),
.Y(n_1153)
);

BUFx8_ASAP7_75t_L g1154 ( 
.A(n_1070),
.Y(n_1154)
);

INVx5_ASAP7_75t_L g1155 ( 
.A(n_976),
.Y(n_1155)
);

AND2x6_ASAP7_75t_L g1156 ( 
.A(n_1058),
.B(n_1081),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_963),
.B(n_968),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1041),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_969),
.A2(n_984),
.B(n_986),
.Y(n_1159)
);

NOR2xp67_ASAP7_75t_L g1160 ( 
.A(n_958),
.B(n_1051),
.Y(n_1160)
);

O2A1O1Ixp5_ASAP7_75t_SL g1161 ( 
.A1(n_1040),
.A2(n_992),
.B(n_1030),
.C(n_1088),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_992),
.A2(n_974),
.B(n_972),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1026),
.B(n_1019),
.Y(n_1163)
);

AO32x2_ASAP7_75t_L g1164 ( 
.A1(n_1028),
.A2(n_1042),
.A3(n_1079),
.B1(n_1004),
.B2(n_1035),
.Y(n_1164)
);

NOR3xp33_ASAP7_75t_L g1165 ( 
.A(n_1040),
.B(n_1015),
.C(n_1001),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_969),
.A2(n_989),
.B(n_1060),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1048),
.B(n_1080),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_995),
.A2(n_1089),
.B(n_1082),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_971),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_996),
.A2(n_998),
.B(n_1005),
.Y(n_1170)
);

AOI21xp33_ASAP7_75t_L g1171 ( 
.A1(n_1023),
.A2(n_1033),
.B(n_973),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1037),
.A2(n_1014),
.B(n_983),
.C(n_965),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1078),
.A2(n_1005),
.B(n_998),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1043),
.A2(n_1022),
.B(n_1017),
.C(n_1016),
.Y(n_1174)
);

INVx5_ASAP7_75t_L g1175 ( 
.A(n_976),
.Y(n_1175)
);

NOR2xp67_ASAP7_75t_L g1176 ( 
.A(n_958),
.B(n_1063),
.Y(n_1176)
);

AOI221x1_ASAP7_75t_L g1177 ( 
.A1(n_996),
.A2(n_1007),
.B1(n_1018),
.B2(n_1027),
.C(n_1063),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1066),
.A2(n_1021),
.B(n_962),
.C(n_967),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1071),
.A2(n_1002),
.B(n_977),
.Y(n_1179)
);

NOR2xp67_ASAP7_75t_L g1180 ( 
.A(n_958),
.B(n_977),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1024),
.B(n_1025),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_991),
.A2(n_1008),
.B(n_1039),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_991),
.A2(n_1008),
.B(n_1039),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_991),
.B(n_1008),
.Y(n_1184)
);

INVxp67_ASAP7_75t_L g1185 ( 
.A(n_1039),
.Y(n_1185)
);

AOI211x1_ASAP7_75t_L g1186 ( 
.A1(n_1011),
.A2(n_1084),
.B(n_1055),
.C(n_988),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1055),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1055),
.A2(n_791),
.B(n_877),
.Y(n_1188)
);

OAI21xp33_ASAP7_75t_L g1189 ( 
.A1(n_1084),
.A2(n_816),
.B(n_791),
.Y(n_1189)
);

AOI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1084),
.A2(n_1068),
.B(n_1049),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_987),
.B(n_623),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1057),
.B(n_819),
.Y(n_1192)
);

INVx5_ASAP7_75t_L g1193 ( 
.A(n_976),
.Y(n_1193)
);

AOI21xp33_ASAP7_75t_L g1194 ( 
.A1(n_980),
.A2(n_877),
.B(n_816),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_994),
.B(n_887),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1057),
.B(n_819),
.Y(n_1196)
);

CKINVDCx6p67_ASAP7_75t_R g1197 ( 
.A(n_959),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_976),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1057),
.B(n_819),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1026),
.B(n_1019),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_964),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_997),
.A2(n_978),
.B(n_955),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_987),
.B(n_623),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_997),
.A2(n_978),
.B(n_955),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_997),
.A2(n_978),
.B(n_955),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_980),
.A2(n_877),
.B(n_791),
.C(n_887),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_987),
.B(n_623),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_964),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_964),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1026),
.B(n_1019),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_976),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1057),
.B(n_819),
.Y(n_1212)
);

O2A1O1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1013),
.A2(n_887),
.B(n_917),
.C(n_904),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1038),
.A2(n_791),
.B(n_877),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_981),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1057),
.A2(n_653),
.B(n_955),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1038),
.A2(n_791),
.B(n_877),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1057),
.A2(n_653),
.B(n_955),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1038),
.A2(n_791),
.B(n_877),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_956),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_976),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_994),
.B(n_887),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_964),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1157),
.B(n_1152),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1115),
.Y(n_1225)
);

AOI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1140),
.A2(n_1142),
.B(n_1124),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1192),
.B(n_1196),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1191),
.B(n_1203),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1205),
.A2(n_1100),
.B(n_1145),
.Y(n_1229)
);

AND2x6_ASAP7_75t_L g1230 ( 
.A(n_1103),
.B(n_1098),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1207),
.B(n_1129),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1104),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1163),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1117),
.A2(n_1219),
.B1(n_1217),
.B2(n_1214),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1094),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1143),
.A2(n_1170),
.B(n_1116),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1169),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1111),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1102),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1112),
.Y(n_1240)
);

AO21x2_ASAP7_75t_L g1241 ( 
.A1(n_1138),
.A2(n_1162),
.B(n_1092),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1136),
.A2(n_1139),
.B(n_1216),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1194),
.A2(n_1189),
.B1(n_1093),
.B2(n_1165),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_L g1244 ( 
.A(n_1206),
.B(n_1213),
.C(n_1161),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1189),
.B(n_1199),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1163),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1108),
.A2(n_1218),
.B(n_1107),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1212),
.B(n_1153),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1113),
.B(n_1137),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1118),
.B(n_1195),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1200),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1222),
.A2(n_1103),
.B1(n_1119),
.B2(n_1121),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1159),
.A2(n_1123),
.B(n_1126),
.Y(n_1253)
);

OAI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1151),
.A2(n_1149),
.B1(n_1131),
.B2(n_1127),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1168),
.A2(n_1095),
.B(n_1128),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1215),
.B(n_1120),
.Y(n_1256)
);

OA21x2_ASAP7_75t_L g1257 ( 
.A1(n_1147),
.A2(n_1097),
.B(n_1173),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1188),
.A2(n_1172),
.B(n_1166),
.C(n_1171),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1132),
.A2(n_1133),
.B(n_1177),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1174),
.A2(n_1178),
.B(n_1122),
.C(n_1135),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1167),
.A2(n_1186),
.B1(n_1160),
.B2(n_1101),
.Y(n_1261)
);

INVx4_ASAP7_75t_L g1262 ( 
.A(n_1155),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1179),
.A2(n_1141),
.B(n_1144),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1201),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1156),
.A2(n_1223),
.B1(n_1208),
.B2(n_1209),
.Y(n_1265)
);

AND2x4_ASAP7_75t_L g1266 ( 
.A(n_1125),
.B(n_1156),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1156),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1155),
.Y(n_1268)
);

INVx1_ASAP7_75t_SL g1269 ( 
.A(n_1114),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1146),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1130),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1134),
.Y(n_1272)
);

AO21x1_ASAP7_75t_L g1273 ( 
.A1(n_1181),
.A2(n_1182),
.B(n_1183),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1158),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_1220),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1156),
.A2(n_1154),
.B1(n_1125),
.B2(n_1096),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1125),
.A2(n_1160),
.B(n_1106),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1099),
.A2(n_1176),
.B(n_1187),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1148),
.B(n_1185),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1164),
.Y(n_1280)
);

BUFx10_ASAP7_75t_L g1281 ( 
.A(n_1210),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1176),
.A2(n_1180),
.B(n_1164),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1154),
.B(n_1184),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1110),
.B(n_1221),
.Y(n_1284)
);

BUFx4f_ASAP7_75t_L g1285 ( 
.A(n_1197),
.Y(n_1285)
);

OR2x6_ASAP7_75t_L g1286 ( 
.A(n_1186),
.B(n_1096),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1180),
.A2(n_1164),
.B(n_1150),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1110),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1110),
.A2(n_1198),
.B1(n_1211),
.B2(n_1221),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1175),
.A2(n_1193),
.B(n_1211),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1104),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1115),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1138),
.A2(n_1162),
.B(n_1202),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1157),
.B(n_1152),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1115),
.Y(n_1295)
);

AO21x2_ASAP7_75t_L g1296 ( 
.A1(n_1214),
.A2(n_1219),
.B(n_1217),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1191),
.B(n_1203),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1117),
.A2(n_887),
.B1(n_917),
.B2(n_904),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1191),
.B(n_1203),
.Y(n_1299)
);

BUFx2_ASAP7_75t_SL g1300 ( 
.A(n_1155),
.Y(n_1300)
);

OR2x6_ASAP7_75t_L g1301 ( 
.A(n_1186),
.B(n_1125),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1190),
.Y(n_1302)
);

AND2x6_ASAP7_75t_L g1303 ( 
.A(n_1103),
.B(n_1081),
.Y(n_1303)
);

AOI22x1_ASAP7_75t_L g1304 ( 
.A1(n_1214),
.A2(n_1219),
.B1(n_1217),
.B2(n_904),
.Y(n_1304)
);

BUFx10_ASAP7_75t_L g1305 ( 
.A(n_1195),
.Y(n_1305)
);

NOR2x1_ASAP7_75t_SL g1306 ( 
.A(n_1125),
.B(n_1068),
.Y(n_1306)
);

INVx3_ASAP7_75t_SL g1307 ( 
.A(n_1220),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1104),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1104),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1151),
.A2(n_1142),
.A3(n_1097),
.B(n_1206),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1191),
.B(n_1203),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1104),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1157),
.B(n_1152),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1109),
.A2(n_1204),
.B(n_1202),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1115),
.Y(n_1315)
);

BUFx2_ASAP7_75t_SL g1316 ( 
.A(n_1155),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_SL g1317 ( 
.A1(n_1105),
.A2(n_1103),
.B(n_1214),
.Y(n_1317)
);

A2O1A1Ixp33_ASAP7_75t_L g1318 ( 
.A1(n_1214),
.A2(n_1219),
.B(n_1217),
.C(n_791),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1202),
.A2(n_1205),
.B(n_1204),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_SL g1320 ( 
.A1(n_1206),
.A2(n_791),
.B(n_1217),
.C(n_1214),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1202),
.A2(n_1205),
.B(n_1204),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1202),
.A2(n_1205),
.B(n_1204),
.Y(n_1322)
);

INVx4_ASAP7_75t_L g1323 ( 
.A(n_1155),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1194),
.A2(n_1217),
.B(n_1219),
.C(n_1214),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1202),
.A2(n_1205),
.B(n_1204),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1194),
.B(n_1189),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1192),
.B(n_1196),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1191),
.B(n_1203),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1104),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1202),
.A2(n_1205),
.B(n_1204),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1157),
.B(n_1152),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1194),
.A2(n_791),
.B1(n_1219),
.B2(n_1217),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1214),
.A2(n_1219),
.B(n_1217),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1194),
.B(n_1214),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1104),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1214),
.A2(n_1219),
.B(n_1217),
.C(n_791),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_1191),
.Y(n_1337)
);

AOI221xp5_ASAP7_75t_L g1338 ( 
.A1(n_1324),
.A2(n_1320),
.B1(n_1333),
.B2(n_1234),
.C(n_1334),
.Y(n_1338)
);

INVx2_ASAP7_75t_SL g1339 ( 
.A(n_1225),
.Y(n_1339)
);

BUFx8_ASAP7_75t_L g1340 ( 
.A(n_1275),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1231),
.B(n_1228),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1332),
.A2(n_1243),
.B1(n_1276),
.B2(n_1336),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1297),
.B(n_1299),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1332),
.A2(n_1276),
.B1(n_1318),
.B2(n_1336),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1252),
.B(n_1337),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_SL g1346 ( 
.A1(n_1318),
.A2(n_1260),
.B(n_1258),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1235),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1227),
.B(n_1327),
.Y(n_1348)
);

AOI31xp33_ASAP7_75t_L g1349 ( 
.A1(n_1261),
.A2(n_1265),
.A3(n_1326),
.B(n_1334),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1250),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1311),
.B(n_1328),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1265),
.A2(n_1304),
.B1(n_1244),
.B2(n_1286),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1266),
.B(n_1301),
.Y(n_1353)
);

A2O1A1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1326),
.A2(n_1253),
.B(n_1258),
.C(n_1245),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1260),
.A2(n_1266),
.B(n_1298),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1225),
.Y(n_1356)
);

OAI211xp5_ASAP7_75t_L g1357 ( 
.A1(n_1320),
.A2(n_1255),
.B(n_1249),
.C(n_1245),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1224),
.B(n_1294),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1313),
.B(n_1331),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1272),
.B(n_1248),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1266),
.B(n_1301),
.Y(n_1361)
);

A2O1A1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1277),
.A2(n_1247),
.B(n_1287),
.C(n_1282),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1254),
.B(n_1230),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1267),
.A2(n_1296),
.B(n_1230),
.C(n_1259),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1237),
.Y(n_1365)
);

AOI221xp5_ASAP7_75t_L g1366 ( 
.A1(n_1254),
.A2(n_1317),
.B1(n_1296),
.B2(n_1241),
.C(n_1256),
.Y(n_1366)
);

O2A1O1Ixp5_ASAP7_75t_L g1367 ( 
.A1(n_1273),
.A2(n_1226),
.B(n_1267),
.C(n_1280),
.Y(n_1367)
);

OAI21xp33_ASAP7_75t_L g1368 ( 
.A1(n_1286),
.A2(n_1256),
.B(n_1239),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_SL g1369 ( 
.A1(n_1306),
.A2(n_1262),
.B(n_1323),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1263),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1263),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1269),
.A2(n_1279),
.B1(n_1315),
.B2(n_1292),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1230),
.B(n_1329),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1263),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1230),
.B(n_1329),
.Y(n_1375)
);

NOR2xp67_ASAP7_75t_L g1376 ( 
.A(n_1232),
.B(n_1291),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1308),
.B(n_1309),
.Y(n_1377)
);

NOR2xp67_ASAP7_75t_L g1378 ( 
.A(n_1312),
.B(n_1335),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1295),
.A2(n_1251),
.B1(n_1246),
.B2(n_1233),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1283),
.A2(n_1264),
.B1(n_1240),
.B2(n_1285),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1230),
.B(n_1270),
.Y(n_1381)
);

OAI22x1_ASAP7_75t_L g1382 ( 
.A1(n_1274),
.A2(n_1280),
.B1(n_1289),
.B2(n_1307),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1257),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1283),
.A2(n_1285),
.B1(n_1238),
.B2(n_1307),
.Y(n_1384)
);

AOI221xp5_ASAP7_75t_L g1385 ( 
.A1(n_1238),
.A2(n_1237),
.B1(n_1271),
.B2(n_1284),
.C(n_1288),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1303),
.B(n_1305),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1305),
.B(n_1281),
.Y(n_1387)
);

INVx1_ASAP7_75t_SL g1388 ( 
.A(n_1275),
.Y(n_1388)
);

INVxp33_ASAP7_75t_L g1389 ( 
.A(n_1284),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1271),
.A2(n_1316),
.B1(n_1300),
.B2(n_1323),
.Y(n_1390)
);

O2A1O1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1293),
.A2(n_1303),
.B(n_1310),
.C(n_1281),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1281),
.B(n_1303),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1242),
.A2(n_1229),
.B(n_1236),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1268),
.A2(n_1303),
.B1(n_1278),
.B2(n_1290),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1268),
.B(n_1314),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1319),
.B(n_1321),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1322),
.B(n_1325),
.Y(n_1397)
);

OA21x2_ASAP7_75t_L g1398 ( 
.A1(n_1322),
.A2(n_1325),
.B(n_1330),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1330),
.A2(n_1186),
.B1(n_887),
.B2(n_917),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1302),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1332),
.A2(n_1186),
.B1(n_887),
.B2(n_917),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1227),
.B(n_1327),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1227),
.B(n_1327),
.Y(n_1403)
);

CKINVDCx14_ASAP7_75t_R g1404 ( 
.A(n_1237),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1237),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1224),
.B(n_1331),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1255),
.A2(n_1259),
.B(n_1247),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1333),
.A2(n_1217),
.B(n_1219),
.C(n_1214),
.Y(n_1408)
);

A2O1A1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1333),
.A2(n_1217),
.B(n_1219),
.C(n_1214),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1224),
.B(n_1331),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1231),
.B(n_1228),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1227),
.B(n_1327),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1332),
.A2(n_1186),
.B1(n_887),
.B2(n_917),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1255),
.A2(n_1259),
.B(n_1247),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1224),
.B(n_1331),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1227),
.B(n_1327),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1266),
.B(n_1301),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1231),
.B(n_1228),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1231),
.B(n_1228),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1371),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1347),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1383),
.B(n_1370),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1383),
.B(n_1370),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1374),
.B(n_1407),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1395),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1396),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1387),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1397),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1356),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1400),
.Y(n_1430)
);

CKINVDCx16_ASAP7_75t_R g1431 ( 
.A(n_1404),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1353),
.B(n_1361),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1362),
.A2(n_1367),
.B(n_1364),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1398),
.Y(n_1434)
);

INVxp67_ASAP7_75t_L g1435 ( 
.A(n_1345),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1400),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1381),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1373),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1375),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1345),
.B(n_1354),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1354),
.B(n_1338),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_1376),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1414),
.B(n_1364),
.Y(n_1443)
);

INVxp67_ASAP7_75t_SL g1444 ( 
.A(n_1391),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1377),
.Y(n_1445)
);

OR2x6_ASAP7_75t_L g1446 ( 
.A(n_1346),
.B(n_1361),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1362),
.A2(n_1408),
.B(n_1409),
.Y(n_1447)
);

OR2x6_ASAP7_75t_L g1448 ( 
.A(n_1417),
.B(n_1355),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1378),
.Y(n_1449)
);

BUFx4f_ASAP7_75t_SL g1450 ( 
.A(n_1340),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1417),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1393),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1349),
.B(n_1401),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1408),
.A2(n_1409),
.B(n_1413),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1363),
.B(n_1359),
.Y(n_1455)
);

AOI222xp33_ASAP7_75t_L g1456 ( 
.A1(n_1342),
.A2(n_1344),
.B1(n_1352),
.B2(n_1366),
.C1(n_1416),
.C2(n_1403),
.Y(n_1456)
);

OR2x6_ASAP7_75t_L g1457 ( 
.A(n_1392),
.B(n_1394),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1435),
.B(n_1360),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1422),
.B(n_1423),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1422),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1446),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1441),
.A2(n_1402),
.B(n_1412),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1420),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1426),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1434),
.Y(n_1465)
);

INVx4_ASAP7_75t_L g1466 ( 
.A(n_1446),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1426),
.B(n_1428),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1434),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1435),
.B(n_1357),
.Y(n_1469)
);

AOI222xp33_ASAP7_75t_L g1470 ( 
.A1(n_1441),
.A2(n_1368),
.B1(n_1348),
.B2(n_1358),
.C1(n_1350),
.C2(n_1351),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1422),
.B(n_1410),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1453),
.A2(n_1343),
.B1(n_1411),
.B2(n_1341),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1456),
.B(n_1386),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1446),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1423),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1437),
.B(n_1415),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1423),
.B(n_1406),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1428),
.B(n_1419),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1452),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1443),
.B(n_1418),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1443),
.B(n_1382),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1453),
.A2(n_1380),
.B1(n_1399),
.B2(n_1385),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1424),
.B(n_1389),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1437),
.B(n_1389),
.Y(n_1484)
);

AOI221xp5_ASAP7_75t_L g1485 ( 
.A1(n_1462),
.A2(n_1454),
.B1(n_1473),
.B2(n_1440),
.C(n_1469),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1463),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1465),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1471),
.Y(n_1488)
);

OAI31xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1473),
.A2(n_1444),
.A3(n_1456),
.B(n_1390),
.Y(n_1489)
);

AOI33xp33_ASAP7_75t_L g1490 ( 
.A1(n_1472),
.A2(n_1438),
.A3(n_1439),
.B1(n_1445),
.B2(n_1449),
.B3(n_1421),
.Y(n_1490)
);

AOI211xp5_ASAP7_75t_L g1491 ( 
.A1(n_1462),
.A2(n_1440),
.B(n_1469),
.C(n_1444),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1483),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1484),
.B(n_1476),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1482),
.A2(n_1446),
.B1(n_1448),
.B2(n_1431),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1463),
.Y(n_1495)
);

OAI31xp33_ASAP7_75t_L g1496 ( 
.A1(n_1482),
.A2(n_1384),
.A3(n_1472),
.B(n_1372),
.Y(n_1496)
);

OAI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1466),
.A2(n_1446),
.B1(n_1448),
.B2(n_1447),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1468),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1463),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1480),
.B(n_1451),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1471),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_SL g1502 ( 
.A1(n_1481),
.A2(n_1447),
.B1(n_1446),
.B2(n_1448),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1480),
.B(n_1425),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_SL g1504 ( 
.A1(n_1481),
.A2(n_1447),
.B1(n_1446),
.B2(n_1448),
.Y(n_1504)
);

AOI221xp5_ASAP7_75t_L g1505 ( 
.A1(n_1484),
.A2(n_1439),
.B1(n_1438),
.B2(n_1442),
.C(n_1449),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1468),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1461),
.B(n_1432),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1459),
.B(n_1430),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1458),
.A2(n_1448),
.B1(n_1431),
.B2(n_1447),
.Y(n_1509)
);

AOI21xp33_ASAP7_75t_L g1510 ( 
.A1(n_1470),
.A2(n_1447),
.B(n_1442),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1466),
.Y(n_1511)
);

OAI221xp5_ASAP7_75t_L g1512 ( 
.A1(n_1470),
.A2(n_1476),
.B1(n_1455),
.B2(n_1448),
.C(n_1461),
.Y(n_1512)
);

NAND3xp33_ASAP7_75t_L g1513 ( 
.A(n_1458),
.B(n_1433),
.C(n_1455),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1459),
.B(n_1430),
.Y(n_1514)
);

NAND2xp33_ASAP7_75t_R g1515 ( 
.A(n_1481),
.B(n_1405),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1459),
.B(n_1436),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1461),
.A2(n_1448),
.B1(n_1457),
.B2(n_1427),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1480),
.B(n_1425),
.Y(n_1518)
);

OAI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1461),
.A2(n_1455),
.B1(n_1457),
.B2(n_1388),
.C(n_1339),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1511),
.B(n_1466),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1492),
.B(n_1467),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1501),
.B(n_1460),
.Y(n_1522)
);

NOR3xp33_ASAP7_75t_SL g1523 ( 
.A(n_1515),
.B(n_1405),
.C(n_1365),
.Y(n_1523)
);

INVx4_ASAP7_75t_SL g1524 ( 
.A(n_1507),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1486),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1498),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1492),
.B(n_1467),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1492),
.B(n_1467),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1486),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1495),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1495),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1499),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_SL g1533 ( 
.A(n_1491),
.B(n_1432),
.Y(n_1533)
);

INVx3_ASAP7_75t_L g1534 ( 
.A(n_1506),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1508),
.Y(n_1535)
);

BUFx8_ASAP7_75t_L g1536 ( 
.A(n_1507),
.Y(n_1536)
);

INVx1_ASAP7_75t_SL g1537 ( 
.A(n_1508),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1487),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1503),
.B(n_1464),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1488),
.B(n_1475),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1503),
.B(n_1464),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1493),
.B(n_1475),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1513),
.B(n_1479),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1513),
.B(n_1479),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1511),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1511),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1499),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1529),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1529),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1530),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1542),
.B(n_1491),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1535),
.B(n_1516),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1530),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1531),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1531),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1524),
.B(n_1511),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1542),
.B(n_1485),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1533),
.B(n_1505),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1524),
.B(n_1518),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1524),
.B(n_1518),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1525),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1540),
.B(n_1471),
.Y(n_1562)
);

NOR3xp33_ASAP7_75t_SL g1563 ( 
.A(n_1533),
.B(n_1512),
.C(n_1519),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_1536),
.Y(n_1564)
);

NOR3xp33_ASAP7_75t_L g1565 ( 
.A(n_1543),
.B(n_1494),
.C(n_1509),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1525),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1524),
.B(n_1507),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1536),
.Y(n_1568)
);

NOR3xp33_ASAP7_75t_L g1569 ( 
.A(n_1543),
.B(n_1510),
.C(n_1497),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1535),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1537),
.B(n_1516),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1537),
.B(n_1490),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1540),
.B(n_1514),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1538),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1543),
.B(n_1514),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1544),
.B(n_1489),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_SL g1577 ( 
.A(n_1523),
.B(n_1489),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1524),
.B(n_1507),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1538),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1544),
.B(n_1478),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1544),
.B(n_1477),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1538),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1532),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1532),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1522),
.B(n_1477),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1524),
.B(n_1500),
.Y(n_1586)
);

INVxp67_ASAP7_75t_L g1587 ( 
.A(n_1545),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1538),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1547),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1521),
.B(n_1500),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1561),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1568),
.B(n_1545),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1557),
.B(n_1539),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1566),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1576),
.A2(n_1502),
.B1(n_1504),
.B2(n_1523),
.Y(n_1595)
);

NOR3xp33_ASAP7_75t_L g1596 ( 
.A(n_1577),
.B(n_1545),
.C(n_1546),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1570),
.B(n_1477),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1583),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1577),
.A2(n_1520),
.B1(n_1536),
.B2(n_1466),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1584),
.Y(n_1600)
);

BUFx3_ASAP7_75t_L g1601 ( 
.A(n_1568),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1568),
.B(n_1545),
.Y(n_1602)
);

OAI21xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1558),
.A2(n_1496),
.B(n_1517),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1565),
.A2(n_1520),
.B1(n_1536),
.B2(n_1466),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1564),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1572),
.B(n_1522),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1556),
.B(n_1546),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1564),
.Y(n_1608)
);

AOI211x1_ASAP7_75t_SL g1609 ( 
.A1(n_1551),
.A2(n_1580),
.B(n_1563),
.C(n_1588),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1589),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1587),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1574),
.Y(n_1612)
);

OAI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1585),
.A2(n_1581),
.B1(n_1562),
.B2(n_1466),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1573),
.B(n_1404),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1556),
.B(n_1546),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1569),
.B(n_1539),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1548),
.Y(n_1617)
);

A2O1A1Ixp33_ASAP7_75t_L g1618 ( 
.A1(n_1581),
.A2(n_1496),
.B(n_1474),
.C(n_1546),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1574),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1549),
.A2(n_1433),
.B1(n_1450),
.B2(n_1474),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1590),
.B(n_1539),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1550),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1573),
.B(n_1450),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1585),
.B(n_1522),
.Y(n_1624)
);

NAND3xp33_ASAP7_75t_L g1625 ( 
.A(n_1553),
.B(n_1536),
.C(n_1433),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1590),
.B(n_1541),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1611),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1605),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1601),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1591),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1601),
.Y(n_1631)
);

NAND3x1_ASAP7_75t_L g1632 ( 
.A(n_1596),
.B(n_1567),
.C(n_1578),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1624),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1595),
.A2(n_1559),
.B1(n_1560),
.B2(n_1520),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1608),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1594),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1607),
.B(n_1556),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1598),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1624),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1606),
.B(n_1575),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1600),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1607),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1597),
.B(n_1575),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1614),
.B(n_1340),
.Y(n_1644)
);

BUFx3_ASAP7_75t_L g1645 ( 
.A(n_1592),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1612),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1592),
.B(n_1559),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1610),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1609),
.B(n_1552),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1617),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1603),
.B(n_1552),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1629),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_SL g1653 ( 
.A1(n_1649),
.A2(n_1625),
.B1(n_1614),
.B2(n_1599),
.Y(n_1653)
);

OAI21xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1634),
.A2(n_1616),
.B(n_1604),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1639),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1639),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1627),
.B(n_1593),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1632),
.A2(n_1618),
.B1(n_1620),
.B2(n_1623),
.Y(n_1658)
);

OAI21x1_ASAP7_75t_SL g1659 ( 
.A1(n_1651),
.A2(n_1622),
.B(n_1619),
.Y(n_1659)
);

AOI21xp33_ASAP7_75t_L g1660 ( 
.A1(n_1632),
.A2(n_1623),
.B(n_1618),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1639),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1633),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1633),
.Y(n_1663)
);

NAND2x1p5_ASAP7_75t_L g1664 ( 
.A(n_1629),
.B(n_1602),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1631),
.Y(n_1665)
);

NOR2x1_ASAP7_75t_L g1666 ( 
.A(n_1631),
.B(n_1602),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1647),
.B(n_1615),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1628),
.B(n_1615),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1645),
.B(n_1637),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1635),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1658),
.B(n_1640),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1652),
.B(n_1642),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1669),
.B(n_1666),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1655),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1656),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1660),
.A2(n_1644),
.B(n_1650),
.Y(n_1676)
);

HB1xp67_ASAP7_75t_L g1677 ( 
.A(n_1664),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1661),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1665),
.B(n_1645),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1662),
.Y(n_1680)
);

AOI31xp33_ASAP7_75t_L g1681 ( 
.A1(n_1670),
.A2(n_1640),
.A3(n_1650),
.B(n_1638),
.Y(n_1681)
);

HAxp5_ASAP7_75t_SL g1682 ( 
.A(n_1680),
.B(n_1663),
.CON(n_1682),
.SN(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1673),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1671),
.A2(n_1653),
.B1(n_1654),
.B2(n_1667),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_1681),
.B(n_1654),
.C(n_1669),
.Y(n_1685)
);

AOI21xp33_ASAP7_75t_L g1686 ( 
.A1(n_1677),
.A2(n_1659),
.B(n_1657),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1673),
.B(n_1637),
.Y(n_1687)
);

OAI21xp5_ASAP7_75t_SL g1688 ( 
.A1(n_1676),
.A2(n_1672),
.B(n_1668),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1676),
.A2(n_1653),
.B1(n_1636),
.B2(n_1648),
.C(n_1641),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1679),
.A2(n_1637),
.B(n_1645),
.Y(n_1690)
);

OAI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1674),
.A2(n_1647),
.B(n_1637),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1683),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1684),
.A2(n_1678),
.B1(n_1675),
.B2(n_1648),
.Y(n_1693)
);

OAI211xp5_ASAP7_75t_L g1694 ( 
.A1(n_1685),
.A2(n_1641),
.B(n_1638),
.C(n_1636),
.Y(n_1694)
);

O2A1O1Ixp5_ASAP7_75t_SL g1695 ( 
.A1(n_1687),
.A2(n_1630),
.B(n_1554),
.C(n_1555),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1691),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1696),
.A2(n_1689),
.B1(n_1686),
.B2(n_1688),
.C(n_1690),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1692),
.B(n_1630),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1694),
.Y(n_1699)
);

NOR2x1_ASAP7_75t_L g1700 ( 
.A(n_1695),
.B(n_1682),
.Y(n_1700)
);

NOR2x1_ASAP7_75t_L g1701 ( 
.A(n_1693),
.B(n_1646),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1692),
.B(n_1643),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1702),
.Y(n_1703)
);

NAND3xp33_ASAP7_75t_L g1704 ( 
.A(n_1700),
.B(n_1646),
.C(n_1643),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_R g1705 ( 
.A(n_1699),
.B(n_1340),
.Y(n_1705)
);

NOR2x1_ASAP7_75t_L g1706 ( 
.A(n_1701),
.B(n_1612),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1697),
.B(n_1621),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1706),
.Y(n_1708)
);

OAI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1704),
.A2(n_1698),
.B(n_1613),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1703),
.B(n_1626),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1709),
.B(n_1707),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1711),
.A2(n_1705),
.B1(n_1708),
.B2(n_1710),
.C(n_1619),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1712),
.A2(n_1579),
.B1(n_1588),
.B2(n_1582),
.Y(n_1713)
);

CKINVDCx20_ASAP7_75t_R g1714 ( 
.A(n_1712),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1714),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1713),
.A2(n_1579),
.B(n_1582),
.Y(n_1716)
);

XNOR2xp5_ASAP7_75t_L g1717 ( 
.A(n_1715),
.B(n_1620),
.Y(n_1717)
);

OAI22x1_ASAP7_75t_L g1718 ( 
.A1(n_1716),
.A2(n_1578),
.B1(n_1567),
.B2(n_1560),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1717),
.Y(n_1719)
);

AOI221x1_ASAP7_75t_L g1720 ( 
.A1(n_1719),
.A2(n_1718),
.B1(n_1534),
.B2(n_1586),
.C(n_1526),
.Y(n_1720)
);

AOI21xp33_ASAP7_75t_L g1721 ( 
.A1(n_1720),
.A2(n_1356),
.B(n_1571),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1586),
.B1(n_1571),
.B2(n_1520),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1722),
.A2(n_1520),
.B1(n_1527),
.B2(n_1528),
.Y(n_1723)
);

AOI211xp5_ASAP7_75t_L g1724 ( 
.A1(n_1723),
.A2(n_1369),
.B(n_1379),
.C(n_1429),
.Y(n_1724)
);


endmodule