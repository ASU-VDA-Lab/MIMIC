module fake_jpeg_10295_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_23),
.B(n_15),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx6p67_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx2_ASAP7_75t_SL g86 ( 
.A(n_44),
.Y(n_86)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_50),
.Y(n_81)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_23),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_55),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_22),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_36),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_38),
.B(n_36),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_62),
.A2(n_40),
.B(n_25),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_54),
.B1(n_29),
.B2(n_26),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_41),
.B1(n_29),
.B2(n_19),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_66),
.A2(n_41),
.B1(n_34),
.B2(n_55),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_59),
.B(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_68),
.B(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_36),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_74),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_36),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_41),
.B1(n_22),
.B2(n_29),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_82),
.B1(n_34),
.B2(n_26),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_36),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_80),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_41),
.B1(n_22),
.B2(n_29),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_17),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_84),
.Y(n_89)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_39),
.Y(n_108)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_90),
.B(n_92),
.Y(n_137)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_105),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_40),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_97),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_40),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_104),
.B1(n_113),
.B2(n_58),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_66),
.A2(n_41),
.B1(n_34),
.B2(n_39),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_40),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_80),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_107),
.A2(n_112),
.B1(n_115),
.B2(n_19),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_105),
.Y(n_134)
);

OAI22x1_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_27),
.B1(n_39),
.B2(n_34),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_111),
.A2(n_85),
.B1(n_72),
.B2(n_70),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_69),
.B1(n_88),
.B2(n_26),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_39),
.B1(n_58),
.B2(n_19),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_72),
.A2(n_24),
.B1(n_19),
.B2(n_39),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_119),
.B1(n_138),
.B2(n_106),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_63),
.B1(n_86),
.B2(n_51),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_120),
.B(n_122),
.Y(n_163)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_125),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_101),
.Y(n_125)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_127),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_84),
.Y(n_129)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_130),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_140),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_92),
.B1(n_99),
.B2(n_96),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_135),
.B1(n_136),
.B2(n_142),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_108),
.B(n_105),
.Y(n_150)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_95),
.A2(n_69),
.B1(n_70),
.B2(n_51),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_87),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_110),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_89),
.B(n_56),
.Y(n_143)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_51),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_97),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_91),
.C(n_108),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_157),
.C(n_165),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_95),
.B1(n_96),
.B2(n_89),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_160),
.B1(n_136),
.B2(n_16),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_150),
.B(n_177),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_151),
.A2(n_153),
.B1(n_161),
.B2(n_173),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_139),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_97),
.Y(n_156)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_91),
.C(n_94),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_117),
.A2(n_60),
.B1(n_103),
.B2(n_24),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_24),
.B1(n_27),
.B2(n_25),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_118),
.A2(n_60),
.B1(n_25),
.B2(n_28),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_162),
.A2(n_166),
.B1(n_152),
.B2(n_163),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_77),
.C(n_75),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_28),
.B1(n_20),
.B2(n_18),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_42),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_116),
.C(n_37),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_0),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_174),
.B(n_175),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_119),
.A2(n_18),
.B1(n_20),
.B2(n_28),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_132),
.B(n_137),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_119),
.A2(n_131),
.B(n_18),
.Y(n_175)
);

O2A1O1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_37),
.B(n_35),
.C(n_42),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_176),
.A2(n_48),
.B1(n_43),
.B2(n_35),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_126),
.A2(n_20),
.B(n_17),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_206),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_121),
.Y(n_180)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_127),
.Y(n_183)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_159),
.B(n_73),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_184),
.B(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_149),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_189),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_127),
.Y(n_186)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_162),
.B1(n_177),
.B2(n_146),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_164),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_196),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_168),
.B(n_67),
.Y(n_191)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_171),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_195),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_0),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_202),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_32),
.Y(n_196)
);

OA22x2_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_154),
.B1(n_48),
.B2(n_43),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_200),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_147),
.B(n_150),
.C(n_156),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_75),
.C(n_124),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_204),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_0),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_151),
.A2(n_48),
.B1(n_43),
.B2(n_33),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_160),
.B1(n_146),
.B2(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_13),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_207),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_208),
.A2(n_229),
.B1(n_30),
.B2(n_32),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_187),
.B1(n_198),
.B2(n_197),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g214 ( 
.A(n_196),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_201),
.Y(n_235)
);

XOR2x2_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_172),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_217),
.A2(n_193),
.B1(n_198),
.B2(n_194),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_155),
.Y(n_219)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_219),
.Y(n_233)
);

AND2x6_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_172),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_222),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_174),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_202),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_225),
.B(n_202),
.Y(n_236)
);

A2O1A1O1Ixp25_ASAP7_75t_L g226 ( 
.A1(n_182),
.A2(n_175),
.B(n_166),
.C(n_32),
.D(n_16),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_30),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_234),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_226),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_237),
.B(n_252),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_193),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_240),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_230),
.B(n_199),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_218),
.B1(n_219),
.B2(n_209),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_248),
.B1(n_249),
.B2(n_229),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_181),
.C(n_190),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_253),
.C(n_247),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_203),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_245),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_194),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_181),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_220),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_205),
.B1(n_75),
.B2(n_33),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_222),
.A2(n_33),
.B1(n_30),
.B2(n_16),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_33),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_212),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_251),
.B(n_245),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_37),
.C(n_35),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_249),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_260),
.C(n_268),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_238),
.A2(n_213),
.B1(n_215),
.B2(n_210),
.Y(n_258)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_224),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_9),
.C(n_14),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_231),
.C(n_220),
.Y(n_260)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_262),
.A2(n_248),
.B1(n_246),
.B2(n_252),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_1),
.Y(n_283)
);

XOR2x2_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_220),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_233),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_267),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_227),
.C(n_229),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_229),
.C(n_212),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_37),
.C(n_35),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_271),
.B(n_278),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_270),
.A2(n_233),
.B1(n_239),
.B2(n_237),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_276),
.B1(n_280),
.B2(n_265),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_274),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_10),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_11),
.B(n_15),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_279),
.A2(n_263),
.B(n_254),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_257),
.A2(n_30),
.B1(n_9),
.B2(n_14),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_284),
.C(n_264),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_7),
.Y(n_295)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_285),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_292),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_288),
.A2(n_296),
.B1(n_277),
.B2(n_293),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_256),
.B(n_269),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_284),
.C(n_7),
.Y(n_303)
);

INVx13_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_291),
.Y(n_301)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_265),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_295),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_298),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_283),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_275),
.C(n_281),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_303),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_6),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_305),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_302),
.A2(n_287),
.B1(n_290),
.B2(n_292),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_307),
.C(n_2),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_300),
.A2(n_295),
.B1(n_6),
.B2(n_5),
.Y(n_307)
);

OA21x2_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_11),
.B(n_12),
.Y(n_309)
);

OAI21xp33_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_2),
.B(n_3),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_304),
.A3(n_299),
.B1(n_301),
.B2(n_298),
.C1(n_12),
.C2(n_37),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_312),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_313),
.A3(n_314),
.B1(n_309),
.B2(n_308),
.C1(n_310),
.C2(n_37),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_308),
.C(n_3),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_3),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_4),
.B(n_302),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_4),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_4),
.Y(n_321)
);


endmodule