module fake_netlist_1_6952_n_1688 (n_117, n_44, n_361, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_360, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_362, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_365, n_179, n_315, n_363, n_86, n_143, n_295, n_263, n_166, n_186, n_364, n_75, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_359, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_343, n_127, n_291, n_170, n_356, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_355, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1688);
input n_117;
input n_44;
input n_361;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_360;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_362;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_365;
input n_179;
input n_315;
input n_363;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_364;
input n_75;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_359;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_343;
input n_127;
input n_291;
input n_170;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_355;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1688;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_1671;
wire n_646;
wire n_1334;
wire n_1627;
wire n_829;
wire n_1603;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1618;
wire n_1477;
wire n_1363;
wire n_1594;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_1646;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_1667;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_1663;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1672;
wire n_1342;
wire n_373;
wire n_1619;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1598;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_1631;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_367;
wire n_1661;
wire n_999;
wire n_769;
wire n_624;
wire n_1597;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1683;
wire n_1349;
wire n_1573;
wire n_1580;
wire n_1605;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_1656;
wire n_571;
wire n_1595;
wire n_1604;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_1654;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_1620;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_1623;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_1613;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1582;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_1662;
wire n_790;
wire n_761;
wire n_1660;
wire n_1287;
wire n_472;
wire n_1100;
wire n_1648;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1682;
wire n_1213;
wire n_1452;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_1639;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1615;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1590;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1628;
wire n_1533;
wire n_1611;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_1563;
wire n_1642;
wire n_824;
wire n_793;
wire n_753;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1600;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_395;
wire n_992;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1681;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1602;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1361;
wire n_1333;
wire n_1557;
wire n_911;
wire n_980;
wire n_1675;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_1606;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1625;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_1629;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1670;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_1581;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_1643;
wire n_1687;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1608;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1050;
wire n_1593;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_1647;
wire n_1621;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1668;
wire n_1153;
wire n_1657;
wire n_1655;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_1665;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_1638;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1645;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_1633;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1626;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_515;
wire n_1577;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1641;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_1583;
wire n_606;
wire n_1585;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_1586;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_1599;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1679;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_1634;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_400;
wire n_1455;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1653;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1640;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1658;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1659;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_1635;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_1576;
wire n_1609;
wire n_832;
wire n_996;
wire n_1578;
wire n_420;
wire n_1684;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1610;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_1678;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1674;
wire n_1351;
wire n_1318;
wire n_956;
wire n_1622;
wire n_1614;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_495;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1612;
wire n_1636;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1587;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1592;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_1624;
wire n_618;
wire n_1596;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1616;
wire n_1378;
wire n_1570;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_1676;
wire n_678;
wire n_1200;
wire n_384;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_401;
wire n_481;
wire n_443;
wire n_694;
wire n_1601;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_1666;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1680;
wire n_1644;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_1669;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1673;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_1589;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_1630;
wire n_784;
wire n_1491;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1637;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1617;
wire n_1632;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_1664;
wire n_682;
wire n_1607;
wire n_906;
wire n_1650;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1591;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_1685;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1677;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1649;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_1686;
wire n_600;
wire n_1531;
wire n_371;
wire n_1548;
wire n_1651;
wire n_1584;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_1588;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_1652;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
BUFx3_ASAP7_75t_L g366 ( .A(n_4), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_175), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_365), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_264), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_291), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_18), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_350), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_100), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_333), .Y(n_374) );
BUFx10_ASAP7_75t_L g375 ( .A(n_41), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_323), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_283), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_354), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_174), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_327), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_329), .Y(n_381) );
BUFx10_ASAP7_75t_L g382 ( .A(n_204), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_258), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_159), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_90), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_356), .Y(n_386) );
CKINVDCx14_ASAP7_75t_R g387 ( .A(n_57), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_312), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_142), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_181), .Y(n_390) );
CKINVDCx16_ASAP7_75t_R g391 ( .A(n_352), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_134), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_194), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_362), .Y(n_394) );
CKINVDCx14_ASAP7_75t_R g395 ( .A(n_34), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_60), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_64), .Y(n_397) );
INVx2_ASAP7_75t_SL g398 ( .A(n_82), .Y(n_398) );
CKINVDCx14_ASAP7_75t_R g399 ( .A(n_295), .Y(n_399) );
BUFx10_ASAP7_75t_L g400 ( .A(n_122), .Y(n_400) );
INVxp67_ASAP7_75t_L g401 ( .A(n_332), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_185), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_146), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_219), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_125), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_190), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_124), .Y(n_407) );
NOR2xp67_ASAP7_75t_L g408 ( .A(n_273), .B(n_80), .Y(n_408) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_191), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_265), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_316), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_315), .B(n_200), .Y(n_412) );
INVxp67_ASAP7_75t_L g413 ( .A(n_276), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_222), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_260), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_1), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_342), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_297), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_77), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_285), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_244), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_53), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_156), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_187), .Y(n_424) );
CKINVDCx16_ASAP7_75t_R g425 ( .A(n_355), .Y(n_425) );
CKINVDCx16_ASAP7_75t_R g426 ( .A(n_2), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_267), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_296), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_0), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_103), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_317), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_287), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_22), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_25), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_307), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_218), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_117), .Y(n_437) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_289), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_16), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_195), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_61), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_292), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_13), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_299), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_220), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_193), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_199), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_58), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_46), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_84), .Y(n_450) );
BUFx3_ASAP7_75t_L g451 ( .A(n_213), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_34), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_61), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_86), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_30), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_172), .Y(n_456) );
NOR2xp67_ASAP7_75t_L g457 ( .A(n_167), .B(n_16), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_178), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_311), .Y(n_459) );
INVxp33_ASAP7_75t_SL g460 ( .A(n_117), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_132), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_364), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_3), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_83), .Y(n_464) );
CKINVDCx16_ASAP7_75t_R g465 ( .A(n_33), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_229), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_50), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_293), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_339), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_171), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_251), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_255), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_221), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_225), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_64), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_147), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_82), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g478 ( .A(n_78), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_304), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_275), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_164), .Y(n_481) );
NOR2xp67_ASAP7_75t_L g482 ( .A(n_77), .B(n_310), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_202), .Y(n_483) );
INVxp33_ASAP7_75t_SL g484 ( .A(n_3), .Y(n_484) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_240), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_52), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_320), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_182), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_111), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_284), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_272), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_155), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_212), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_141), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_119), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_80), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_49), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_138), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_210), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_47), .Y(n_500) );
BUFx3_ASAP7_75t_L g501 ( .A(n_8), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_149), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_241), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_223), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_336), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_319), .Y(n_506) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_290), .Y(n_507) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_24), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_318), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_55), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_226), .Y(n_511) );
INVxp67_ASAP7_75t_L g512 ( .A(n_169), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_262), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_57), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_176), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_279), .Y(n_516) );
CKINVDCx14_ASAP7_75t_R g517 ( .A(n_158), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_39), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_130), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_201), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_118), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_186), .Y(n_522) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_207), .Y(n_523) );
NOR2xp67_ASAP7_75t_L g524 ( .A(n_298), .B(n_346), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_165), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_180), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_254), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_321), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_341), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_231), .Y(n_530) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_237), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_66), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_59), .Y(n_533) );
BUFx10_ASAP7_75t_L g534 ( .A(n_134), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_314), .Y(n_535) );
CKINVDCx16_ASAP7_75t_R g536 ( .A(n_75), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_236), .Y(n_537) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_211), .Y(n_538) );
BUFx3_ASAP7_75t_L g539 ( .A(n_66), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_261), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_330), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_88), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_39), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_196), .Y(n_544) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_286), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_179), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_115), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_348), .Y(n_548) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_161), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_249), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_8), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_131), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_177), .Y(n_553) );
BUFx3_ASAP7_75t_L g554 ( .A(n_92), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_123), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_256), .Y(n_556) );
CKINVDCx16_ASAP7_75t_R g557 ( .A(n_114), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_300), .Y(n_558) );
BUFx2_ASAP7_75t_L g559 ( .A(n_305), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_170), .Y(n_560) );
OAI22xp5_ASAP7_75t_SL g561 ( .A1(n_407), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_561) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_438), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_434), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_392), .B(n_5), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_434), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_430), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_386), .Y(n_567) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_438), .Y(n_568) );
AND2x6_ASAP7_75t_L g569 ( .A(n_378), .B(n_157), .Y(n_569) );
BUFx2_ASAP7_75t_L g570 ( .A(n_387), .Y(n_570) );
BUFx2_ASAP7_75t_L g571 ( .A(n_387), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_370), .B(n_5), .Y(n_572) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_438), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_395), .A2(n_9), .B1(n_6), .B2(n_7), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_443), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_395), .A2(n_9), .B1(n_6), .B2(n_7), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_366), .B(n_10), .Y(n_577) );
BUFx8_ASAP7_75t_L g578 ( .A(n_377), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_443), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_386), .Y(n_580) );
INVx3_ASAP7_75t_L g581 ( .A(n_382), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_453), .Y(n_582) );
NAND2xp33_ASAP7_75t_L g583 ( .A(n_390), .B(n_363), .Y(n_583) );
AND2x4_ASAP7_75t_L g584 ( .A(n_366), .B(n_10), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_453), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_475), .Y(n_586) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_438), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_475), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_460), .A2(n_13), .B1(n_11), .B2(n_12), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_446), .B(n_559), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_428), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_398), .B(n_11), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_477), .Y(n_593) );
BUFx3_ASAP7_75t_L g594 ( .A(n_378), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_405), .Y(n_595) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_485), .Y(n_596) );
INVx3_ASAP7_75t_L g597 ( .A(n_382), .Y(n_597) );
NOR2x1_ASAP7_75t_L g598 ( .A(n_501), .B(n_12), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_477), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_428), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_444), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_426), .B(n_14), .Y(n_602) );
INVx3_ASAP7_75t_L g603 ( .A(n_577), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_562), .Y(n_604) );
AND2x2_ASAP7_75t_SL g605 ( .A(n_577), .B(n_391), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_570), .B(n_425), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_567), .Y(n_607) );
INVx8_ASAP7_75t_L g608 ( .A(n_569), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_581), .B(n_405), .Y(n_609) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_562), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_562), .Y(n_611) );
BUFx3_ASAP7_75t_L g612 ( .A(n_569), .Y(n_612) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_570), .Y(n_613) );
CKINVDCx8_ASAP7_75t_R g614 ( .A(n_571), .Y(n_614) );
AO22x2_ASAP7_75t_L g615 ( .A1(n_574), .A2(n_532), .B1(n_551), .B2(n_502), .Y(n_615) );
BUFx4f_ASAP7_75t_L g616 ( .A(n_569), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_577), .A2(n_484), .B1(n_460), .B2(n_478), .Y(n_617) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_562), .Y(n_618) );
BUFx3_ASAP7_75t_L g619 ( .A(n_569), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_571), .B(n_465), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_562), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_562), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_567), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_578), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_580), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_580), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_581), .B(n_401), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_566), .B(n_492), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_577), .A2(n_484), .B1(n_557), .B2(n_536), .Y(n_629) );
BUFx4f_ASAP7_75t_L g630 ( .A(n_569), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_581), .B(n_382), .Y(n_631) );
INVxp33_ASAP7_75t_L g632 ( .A(n_595), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_591), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_591), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_568), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_568), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_581), .B(n_399), .Y(n_637) );
INVx4_ASAP7_75t_L g638 ( .A(n_569), .Y(n_638) );
INVx3_ASAP7_75t_L g639 ( .A(n_584), .Y(n_639) );
BUFx3_ASAP7_75t_L g640 ( .A(n_569), .Y(n_640) );
INVx2_ASAP7_75t_SL g641 ( .A(n_597), .Y(n_641) );
AND2x6_ASAP7_75t_L g642 ( .A(n_584), .B(n_598), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_597), .B(n_413), .Y(n_643) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_568), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_607), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_605), .A2(n_578), .B1(n_597), .B2(n_584), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_632), .B(n_590), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_642), .A2(n_584), .B1(n_601), .B2(n_600), .Y(n_648) );
O2A1O1Ixp5_ASAP7_75t_L g649 ( .A1(n_616), .A2(n_572), .B(n_592), .C(n_564), .Y(n_649) );
INVx4_ASAP7_75t_L g650 ( .A(n_608), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_607), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_637), .B(n_578), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_623), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_637), .B(n_578), .Y(n_654) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_612), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_605), .A2(n_602), .B1(n_583), .B2(n_576), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_628), .B(n_441), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_623), .Y(n_658) );
BUFx5_ASAP7_75t_L g659 ( .A(n_612), .Y(n_659) );
BUFx2_ASAP7_75t_L g660 ( .A(n_613), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_609), .B(n_594), .Y(n_661) );
INVx4_ASAP7_75t_L g662 ( .A(n_608), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_603), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_625), .Y(n_664) );
INVx3_ASAP7_75t_L g665 ( .A(n_603), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_627), .B(n_594), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_628), .B(n_441), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_643), .B(n_594), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_605), .B(n_368), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_603), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_617), .A2(n_458), .B1(n_481), .B2(n_424), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_638), .B(n_367), .Y(n_672) );
OAI22xp5_ASAP7_75t_SL g673 ( .A1(n_629), .A2(n_561), .B1(n_433), .B2(n_497), .Y(n_673) );
NOR2x2_ASAP7_75t_L g674 ( .A(n_614), .B(n_407), .Y(n_674) );
OR2x6_ASAP7_75t_L g675 ( .A(n_620), .B(n_561), .Y(n_675) );
AND2x6_ASAP7_75t_SL g676 ( .A(n_614), .B(n_371), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_638), .B(n_369), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_625), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_626), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_631), .B(n_563), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_642), .B(n_394), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_638), .B(n_372), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_638), .B(n_376), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_642), .B(n_394), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_603), .Y(n_685) );
INVx2_ASAP7_75t_SL g686 ( .A(n_620), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_639), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_639), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_626), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_639), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_642), .B(n_404), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_639), .Y(n_692) );
O2A1O1Ixp33_ASAP7_75t_L g693 ( .A1(n_606), .A2(n_601), .B(n_600), .C(n_565), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_642), .B(n_404), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_616), .B(n_379), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_642), .B(n_406), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_642), .B(n_406), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_633), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_642), .B(n_410), .Y(n_699) );
BUFx12f_ASAP7_75t_L g700 ( .A(n_624), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_629), .B(n_375), .Y(n_701) );
NAND2xp33_ASAP7_75t_L g702 ( .A(n_608), .B(n_412), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_633), .Y(n_703) );
BUFx3_ASAP7_75t_L g704 ( .A(n_612), .Y(n_704) );
INVx2_ASAP7_75t_SL g705 ( .A(n_641), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_634), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_634), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_615), .A2(n_565), .B1(n_575), .B2(n_563), .Y(n_708) );
INVx2_ASAP7_75t_SL g709 ( .A(n_641), .Y(n_709) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_616), .B(n_381), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_617), .A2(n_458), .B1(n_481), .B2(n_424), .Y(n_711) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_630), .B(n_383), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_615), .A2(n_579), .B1(n_582), .B2(n_575), .Y(n_713) );
BUFx3_ASAP7_75t_L g714 ( .A(n_619), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_630), .B(n_384), .Y(n_715) );
AND3x1_ASAP7_75t_L g716 ( .A(n_615), .B(n_589), .C(n_598), .Y(n_716) );
AND2x4_ASAP7_75t_L g717 ( .A(n_619), .B(n_589), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_619), .B(n_410), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_630), .B(n_388), .Y(n_719) );
NOR3x1_ASAP7_75t_L g720 ( .A(n_615), .B(n_497), .C(n_433), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_640), .B(n_462), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_640), .Y(n_722) );
AND2x4_ASAP7_75t_L g723 ( .A(n_640), .B(n_579), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_630), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_608), .A2(n_585), .B1(n_586), .B2(n_582), .Y(n_725) );
NOR2xp67_ASAP7_75t_L g726 ( .A(n_611), .B(n_585), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_608), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_611), .B(n_375), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_611), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_622), .Y(n_730) );
BUFx2_ASAP7_75t_L g731 ( .A(n_622), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_622), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_672), .A2(n_409), .B(n_374), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_672), .A2(n_523), .B(n_507), .Y(n_734) );
INVx3_ASAP7_75t_L g735 ( .A(n_665), .Y(n_735) );
NAND2xp5_ASAP7_75t_SL g736 ( .A(n_704), .B(n_462), .Y(n_736) );
OR2x2_ASAP7_75t_L g737 ( .A(n_647), .B(n_454), .Y(n_737) );
BUFx12f_ASAP7_75t_L g738 ( .A(n_676), .Y(n_738) );
O2A1O1Ixp33_ASAP7_75t_L g739 ( .A1(n_657), .A2(n_397), .B(n_403), .C(n_389), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_665), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_669), .B(n_455), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_648), .A2(n_511), .B1(n_527), .B2(n_525), .Y(n_742) );
NOR3xp33_ASAP7_75t_L g743 ( .A(n_673), .B(n_495), .C(n_396), .Y(n_743) );
AOI31xp33_ASAP7_75t_L g744 ( .A1(n_716), .A2(n_517), .A3(n_518), .B(n_455), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_648), .A2(n_525), .B1(n_527), .B2(n_511), .Y(n_745) );
NOR2xp33_ASAP7_75t_R g746 ( .A(n_700), .B(n_548), .Y(n_746) );
BUFx2_ASAP7_75t_L g747 ( .A(n_660), .Y(n_747) );
AND2x4_ASAP7_75t_L g748 ( .A(n_717), .B(n_548), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_663), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_646), .A2(n_556), .B1(n_555), .B2(n_518), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_717), .A2(n_556), .B1(n_555), .B2(n_553), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_717), .A2(n_553), .B1(n_560), .B2(n_549), .Y(n_752) );
BUFx6f_ASAP7_75t_SL g753 ( .A(n_675), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_656), .A2(n_560), .B1(n_549), .B2(n_419), .Y(n_754) );
INVx4_ASAP7_75t_L g755 ( .A(n_700), .Y(n_755) );
BUFx3_ASAP7_75t_L g756 ( .A(n_707), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_708), .A2(n_416), .B1(n_429), .B2(n_422), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_686), .B(n_667), .Y(n_758) );
O2A1O1Ixp33_ASAP7_75t_L g759 ( .A1(n_708), .A2(n_439), .B(n_448), .C(n_437), .Y(n_759) );
CKINVDCx5p33_ASAP7_75t_R g760 ( .A(n_671), .Y(n_760) );
A2O1A1Ixp33_ASAP7_75t_L g761 ( .A1(n_649), .A2(n_539), .B(n_554), .C(n_501), .Y(n_761) );
AO32x2_ASAP7_75t_L g762 ( .A1(n_705), .A2(n_408), .A3(n_482), .B1(n_457), .B2(n_568), .Y(n_762) );
NOR3xp33_ASAP7_75t_SL g763 ( .A(n_674), .B(n_385), .C(n_373), .Y(n_763) );
NOR3xp33_ASAP7_75t_SL g764 ( .A(n_674), .B(n_514), .C(n_500), .Y(n_764) );
A2O1A1Ixp33_ASAP7_75t_L g765 ( .A1(n_663), .A2(n_554), .B(n_539), .C(n_450), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_677), .A2(n_402), .B(n_393), .Y(n_766) );
O2A1O1Ixp33_ASAP7_75t_L g767 ( .A1(n_713), .A2(n_452), .B(n_461), .C(n_449), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_652), .B(n_521), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_654), .B(n_533), .Y(n_769) );
A2O1A1Ixp33_ASAP7_75t_L g770 ( .A1(n_670), .A2(n_464), .B(n_467), .C(n_463), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_682), .A2(n_417), .B(n_415), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_701), .B(n_375), .Y(n_772) );
AOI21xp5_ASAP7_75t_L g773 ( .A1(n_683), .A2(n_436), .B(n_431), .Y(n_773) );
BUFx6f_ASAP7_75t_L g774 ( .A(n_704), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g775 ( .A1(n_683), .A2(n_447), .B(n_440), .Y(n_775) );
NAND3xp33_ASAP7_75t_SL g776 ( .A(n_713), .B(n_442), .C(n_411), .Y(n_776) );
AOI221xp5_ASAP7_75t_L g777 ( .A1(n_711), .A2(n_489), .B1(n_494), .B2(n_486), .C(n_476), .Y(n_777) );
O2A1O1Ixp33_ASAP7_75t_L g778 ( .A1(n_675), .A2(n_498), .B(n_510), .C(n_496), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_661), .A2(n_668), .B(n_666), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_681), .B(n_400), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_684), .B(n_400), .Y(n_781) );
OAI22x1_ASAP7_75t_L g782 ( .A1(n_675), .A2(n_519), .B1(n_543), .B2(n_542), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_702), .A2(n_400), .B1(n_534), .B2(n_547), .Y(n_783) );
OAI21xp5_ASAP7_75t_L g784 ( .A1(n_670), .A2(n_466), .B(n_459), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_685), .Y(n_785) );
A2O1A1Ixp33_ASAP7_75t_L g786 ( .A1(n_685), .A2(n_552), .B(n_593), .C(n_588), .Y(n_786) );
OR2x6_ASAP7_75t_L g787 ( .A(n_650), .B(n_502), .Y(n_787) );
INVx4_ASAP7_75t_L g788 ( .A(n_650), .Y(n_788) );
O2A1O1Ixp33_ASAP7_75t_L g789 ( .A1(n_645), .A2(n_551), .B(n_532), .C(n_599), .Y(n_789) );
A2O1A1Ixp33_ASAP7_75t_L g790 ( .A1(n_687), .A2(n_599), .B(n_469), .C(n_470), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_720), .B(n_534), .Y(n_791) );
NOR2xp33_ASAP7_75t_R g792 ( .A(n_691), .B(n_534), .Y(n_792) );
NAND2x1p5_ASAP7_75t_L g793 ( .A(n_662), .B(n_508), .Y(n_793) );
BUFx8_ASAP7_75t_L g794 ( .A(n_728), .Y(n_794) );
NAND2xp5_ASAP7_75t_SL g795 ( .A(n_714), .B(n_380), .Y(n_795) );
BUFx2_ASAP7_75t_L g796 ( .A(n_723), .Y(n_796) );
O2A1O1Ixp33_ASAP7_75t_L g797 ( .A1(n_651), .A2(n_420), .B(n_512), .C(n_414), .Y(n_797) );
AOI21x1_ASAP7_75t_L g798 ( .A1(n_695), .A2(n_621), .B(n_604), .Y(n_798) );
BUFx6f_ASAP7_75t_L g799 ( .A(n_714), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_687), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_707), .B(n_418), .Y(n_801) );
AOI21xp5_ASAP7_75t_L g802 ( .A1(n_695), .A2(n_712), .B(n_710), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_688), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_694), .A2(n_472), .B1(n_473), .B2(n_468), .Y(n_804) );
AND2x4_ASAP7_75t_L g805 ( .A(n_662), .B(n_474), .Y(n_805) );
O2A1O1Ixp5_ASAP7_75t_L g806 ( .A1(n_710), .A2(n_444), .B(n_456), .C(n_445), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_680), .B(n_423), .Y(n_807) );
BUFx2_ASAP7_75t_L g808 ( .A(n_723), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_688), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_725), .B(n_427), .Y(n_810) );
O2A1O1Ixp33_ASAP7_75t_L g811 ( .A1(n_653), .A2(n_480), .B(n_483), .C(n_479), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_725), .B(n_432), .Y(n_812) );
OAI21xp5_ASAP7_75t_L g813 ( .A1(n_690), .A2(n_488), .B(n_487), .Y(n_813) );
INVx4_ASAP7_75t_L g814 ( .A(n_723), .Y(n_814) );
NOR2xp67_ASAP7_75t_L g815 ( .A(n_696), .B(n_14), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_697), .B(n_435), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_712), .A2(n_499), .B(n_491), .Y(n_817) );
OAI22xp5_ASAP7_75t_SL g818 ( .A1(n_699), .A2(n_490), .B1(n_493), .B2(n_471), .Y(n_818) );
INVxp67_ASAP7_75t_SL g819 ( .A(n_655), .Y(n_819) );
BUFx2_ASAP7_75t_SL g820 ( .A(n_709), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_658), .B(n_505), .Y(n_821) );
NAND2xp5_ASAP7_75t_SL g822 ( .A(n_655), .B(n_506), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_664), .B(n_508), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_678), .A2(n_504), .B1(n_513), .B2(n_503), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_690), .Y(n_825) );
NAND2xp5_ASAP7_75t_SL g826 ( .A(n_655), .B(n_509), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_679), .B(n_528), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_689), .A2(n_508), .B1(n_516), .B2(n_515), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_698), .B(n_529), .Y(n_829) );
A2O1A1Ixp33_ASAP7_75t_L g830 ( .A1(n_692), .A2(n_522), .B(n_526), .C(n_520), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_703), .B(n_530), .Y(n_831) );
O2A1O1Ixp33_ASAP7_75t_SL g832 ( .A1(n_724), .A2(n_537), .B(n_540), .C(n_535), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_692), .Y(n_833) );
AND2x4_ASAP7_75t_L g834 ( .A(n_727), .B(n_541), .Y(n_834) );
BUFx2_ASAP7_75t_L g835 ( .A(n_706), .Y(n_835) );
NOR2xp33_ASAP7_75t_L g836 ( .A(n_715), .B(n_544), .Y(n_836) );
INVx3_ASAP7_75t_SL g837 ( .A(n_715), .Y(n_837) );
NAND2xp5_ASAP7_75t_SL g838 ( .A(n_659), .B(n_546), .Y(n_838) );
BUFx6f_ASAP7_75t_L g839 ( .A(n_731), .Y(n_839) );
BUFx2_ASAP7_75t_L g840 ( .A(n_718), .Y(n_840) );
NAND3xp33_ASAP7_75t_L g841 ( .A(n_693), .B(n_508), .C(n_550), .Y(n_841) );
AOI21xp5_ASAP7_75t_L g842 ( .A1(n_719), .A2(n_558), .B(n_456), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_726), .A2(n_445), .B1(n_451), .B2(n_421), .Y(n_843) );
A2O1A1Ixp33_ASAP7_75t_L g844 ( .A1(n_722), .A2(n_524), .B(n_451), .C(n_421), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_732), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_721), .B(n_15), .Y(n_846) );
INVx3_ASAP7_75t_L g847 ( .A(n_659), .Y(n_847) );
NAND2xp5_ASAP7_75t_SL g848 ( .A(n_659), .B(n_485), .Y(n_848) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_659), .B(n_15), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_659), .B(n_17), .Y(n_850) );
BUFx3_ASAP7_75t_L g851 ( .A(n_729), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_730), .Y(n_852) );
O2A1O1Ixp5_ASAP7_75t_L g853 ( .A1(n_659), .A2(n_636), .B(n_635), .C(n_531), .Y(n_853) );
O2A1O1Ixp33_ASAP7_75t_SL g854 ( .A1(n_724), .A2(n_636), .B(n_635), .C(n_162), .Y(n_854) );
CKINVDCx6p67_ASAP7_75t_R g855 ( .A(n_700), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_665), .Y(n_856) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_660), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_665), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g859 ( .A(n_657), .B(n_17), .Y(n_859) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_657), .B(n_18), .Y(n_860) );
INVx2_ASAP7_75t_L g861 ( .A(n_665), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_665), .Y(n_862) );
AOI21xp5_ASAP7_75t_L g863 ( .A1(n_672), .A2(n_618), .B(n_610), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_657), .B(n_19), .Y(n_864) );
OAI22xp5_ASAP7_75t_SL g865 ( .A1(n_673), .A2(n_531), .B1(n_538), .B2(n_485), .Y(n_865) );
INVx2_ASAP7_75t_L g866 ( .A(n_665), .Y(n_866) );
OAI21xp5_ASAP7_75t_L g867 ( .A1(n_649), .A2(n_618), .B(n_610), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_835), .Y(n_868) );
AOI21xp5_ASAP7_75t_L g869 ( .A1(n_867), .A2(n_618), .B(n_610), .Y(n_869) );
AOI21xp5_ASAP7_75t_L g870 ( .A1(n_867), .A2(n_618), .B(n_610), .Y(n_870) );
INVx3_ASAP7_75t_L g871 ( .A(n_788), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_758), .B(n_19), .Y(n_872) );
AOI21xp5_ASAP7_75t_L g873 ( .A1(n_779), .A2(n_618), .B(n_610), .Y(n_873) );
AOI21xp5_ASAP7_75t_L g874 ( .A1(n_802), .A2(n_618), .B(n_610), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_748), .A2(n_531), .B1(n_538), .B2(n_485), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_748), .A2(n_538), .B1(n_545), .B2(n_531), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_823), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_834), .Y(n_878) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_760), .B(n_20), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_745), .A2(n_545), .B1(n_538), .B2(n_568), .Y(n_880) );
OAI21xp5_ASAP7_75t_L g881 ( .A1(n_761), .A2(n_573), .B(n_568), .Y(n_881) );
AOI221x1_ASAP7_75t_L g882 ( .A1(n_844), .A2(n_587), .B1(n_596), .B2(n_573), .C(n_545), .Y(n_882) );
AND2x4_ASAP7_75t_L g883 ( .A(n_788), .B(n_20), .Y(n_883) );
OAI21xp5_ASAP7_75t_L g884 ( .A1(n_841), .A2(n_587), .B(n_573), .Y(n_884) );
CKINVDCx12_ASAP7_75t_R g885 ( .A(n_787), .Y(n_885) );
A2O1A1Ixp33_ASAP7_75t_L g886 ( .A1(n_789), .A2(n_545), .B(n_587), .C(n_573), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_756), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g888 ( .A(n_751), .B(n_21), .Y(n_888) );
NAND2xp33_ASAP7_75t_SL g889 ( .A(n_745), .B(n_21), .Y(n_889) );
AOI21xp5_ASAP7_75t_L g890 ( .A1(n_863), .A2(n_644), .B(n_587), .Y(n_890) );
OR2x2_ASAP7_75t_L g891 ( .A(n_747), .B(n_22), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_834), .Y(n_892) );
BUFx2_ASAP7_75t_L g893 ( .A(n_857), .Y(n_893) );
NOR2xp33_ASAP7_75t_L g894 ( .A(n_772), .B(n_23), .Y(n_894) );
AND2x6_ASAP7_75t_L g895 ( .A(n_850), .B(n_573), .Y(n_895) );
AOI22xp33_ASAP7_75t_SL g896 ( .A1(n_742), .A2(n_26), .B1(n_24), .B2(n_25), .Y(n_896) );
O2A1O1Ixp33_ASAP7_75t_L g897 ( .A1(n_739), .A2(n_28), .B(n_26), .C(n_27), .Y(n_897) );
CKINVDCx5p33_ASAP7_75t_R g898 ( .A(n_855), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_746), .A2(n_29), .B1(n_27), .B2(n_28), .Y(n_899) );
OR2x6_ASAP7_75t_L g900 ( .A(n_755), .B(n_29), .Y(n_900) );
INVx5_ASAP7_75t_L g901 ( .A(n_787), .Y(n_901) );
A2O1A1Ixp33_ASAP7_75t_L g902 ( .A1(n_859), .A2(n_587), .B(n_596), .C(n_573), .Y(n_902) );
OAI21x1_ASAP7_75t_L g903 ( .A1(n_798), .A2(n_596), .B(n_587), .Y(n_903) );
AND2x6_ASAP7_75t_L g904 ( .A(n_774), .B(n_596), .Y(n_904) );
AO31x2_ASAP7_75t_L g905 ( .A1(n_849), .A2(n_596), .A3(n_644), .B(n_32), .Y(n_905) );
HB1xp67_ASAP7_75t_L g906 ( .A(n_839), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_786), .Y(n_907) );
BUFx6f_ASAP7_75t_L g908 ( .A(n_839), .Y(n_908) );
INVx1_ASAP7_75t_SL g909 ( .A(n_737), .Y(n_909) );
OAI21x1_ASAP7_75t_L g910 ( .A1(n_853), .A2(n_163), .B(n_160), .Y(n_910) );
A2O1A1Ixp33_ASAP7_75t_L g911 ( .A1(n_860), .A2(n_644), .B(n_35), .C(n_30), .Y(n_911) );
AO32x2_ASAP7_75t_L g912 ( .A1(n_757), .A2(n_31), .A3(n_35), .B1(n_36), .B2(n_37), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_765), .Y(n_913) );
BUFx8_ASAP7_75t_L g914 ( .A(n_753), .Y(n_914) );
A2O1A1Ixp33_ASAP7_75t_L g915 ( .A1(n_864), .A2(n_644), .B(n_37), .C(n_31), .Y(n_915) );
AND2x6_ASAP7_75t_L g916 ( .A(n_774), .B(n_36), .Y(n_916) );
AOI21xp5_ASAP7_75t_L g917 ( .A1(n_852), .A2(n_644), .B(n_168), .Y(n_917) );
A2O1A1Ixp33_ASAP7_75t_L g918 ( .A1(n_811), .A2(n_41), .B(n_38), .C(n_40), .Y(n_918) );
NAND2xp5_ASAP7_75t_SL g919 ( .A(n_839), .B(n_38), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_777), .B(n_40), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_770), .Y(n_921) );
OR2x2_ASAP7_75t_L g922 ( .A(n_752), .B(n_42), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_794), .B(n_42), .Y(n_923) );
CKINVDCx5p33_ASAP7_75t_R g924 ( .A(n_738), .Y(n_924) );
OAI21xp5_ASAP7_75t_L g925 ( .A1(n_841), .A2(n_173), .B(n_166), .Y(n_925) );
NOR2x1_ASAP7_75t_SL g926 ( .A(n_787), .B(n_43), .Y(n_926) );
INVx2_ASAP7_75t_SL g927 ( .A(n_755), .Y(n_927) );
AO31x2_ASAP7_75t_L g928 ( .A1(n_757), .A2(n_45), .A3(n_43), .B(n_44), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_794), .B(n_44), .Y(n_929) );
INVxp67_ASAP7_75t_SL g930 ( .A(n_796), .Y(n_930) );
INVx4_ASAP7_75t_L g931 ( .A(n_814), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_750), .B(n_45), .Y(n_932) );
AO31x2_ASAP7_75t_L g933 ( .A1(n_790), .A2(n_48), .A3(n_46), .B(n_47), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_743), .A2(n_50), .B1(n_48), .B2(n_49), .Y(n_934) );
BUFx6f_ASAP7_75t_L g935 ( .A(n_774), .Y(n_935) );
AND2x2_ASAP7_75t_L g936 ( .A(n_763), .B(n_51), .Y(n_936) );
OAI21x1_ASAP7_75t_L g937 ( .A1(n_848), .A2(n_184), .B(n_183), .Y(n_937) );
AOI22xp33_ASAP7_75t_SL g938 ( .A1(n_865), .A2(n_753), .B1(n_791), .B2(n_820), .Y(n_938) );
INVx4_ASAP7_75t_L g939 ( .A(n_814), .Y(n_939) );
NOR2xp67_ASAP7_75t_SL g940 ( .A(n_799), .B(n_51), .Y(n_940) );
INVx4_ASAP7_75t_L g941 ( .A(n_793), .Y(n_941) );
CKINVDCx11_ASAP7_75t_R g942 ( .A(n_837), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_759), .Y(n_943) );
NOR2xp33_ASAP7_75t_L g944 ( .A(n_744), .B(n_52), .Y(n_944) );
A2O1A1Ixp33_ASAP7_75t_L g945 ( .A1(n_836), .A2(n_56), .B(n_53), .C(n_54), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_764), .B(n_54), .Y(n_946) );
NOR2xp33_ASAP7_75t_L g947 ( .A(n_768), .B(n_56), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_741), .B(n_58), .Y(n_948) );
AOI21xp5_ASAP7_75t_L g949 ( .A1(n_838), .A2(n_189), .B(n_188), .Y(n_949) );
NOR2xp33_ASAP7_75t_SL g950 ( .A(n_776), .B(n_59), .Y(n_950) );
AOI21xp5_ASAP7_75t_L g951 ( .A1(n_769), .A2(n_197), .B(n_192), .Y(n_951) );
NOR3xp33_ASAP7_75t_L g952 ( .A(n_778), .B(n_60), .C(n_62), .Y(n_952) );
AO32x2_ASAP7_75t_L g953 ( .A1(n_843), .A2(n_62), .A3(n_63), .B1(n_65), .B2(n_67), .Y(n_953) );
HB1xp67_ASAP7_75t_L g954 ( .A(n_808), .Y(n_954) );
BUFx2_ASAP7_75t_SL g955 ( .A(n_805), .Y(n_955) );
AND2x4_ASAP7_75t_L g956 ( .A(n_840), .B(n_63), .Y(n_956) );
AOI21xp5_ASAP7_75t_L g957 ( .A1(n_801), .A2(n_203), .B(n_198), .Y(n_957) );
NOR2xp33_ASAP7_75t_L g958 ( .A(n_754), .B(n_65), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_782), .B(n_67), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_805), .B(n_68), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_783), .B(n_68), .Y(n_961) );
NOR2x1_ASAP7_75t_L g962 ( .A(n_767), .B(n_736), .Y(n_962) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_797), .B(n_69), .Y(n_963) );
INVx2_ASAP7_75t_L g964 ( .A(n_749), .Y(n_964) );
INVx2_ASAP7_75t_SL g965 ( .A(n_792), .Y(n_965) );
INVx4_ASAP7_75t_L g966 ( .A(n_799), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_803), .Y(n_967) );
AO31x2_ASAP7_75t_L g968 ( .A1(n_843), .A2(n_69), .A3(n_70), .B(n_71), .Y(n_968) );
INVx2_ASAP7_75t_L g969 ( .A(n_785), .Y(n_969) );
OAI21xp5_ASAP7_75t_L g970 ( .A1(n_806), .A2(n_206), .B(n_205), .Y(n_970) );
OAI21xp5_ASAP7_75t_L g971 ( .A1(n_784), .A2(n_209), .B(n_208), .Y(n_971) );
AOI21xp5_ASAP7_75t_L g972 ( .A1(n_821), .A2(n_215), .B(n_214), .Y(n_972) );
A2O1A1Ixp33_ASAP7_75t_L g973 ( .A1(n_842), .A2(n_70), .B(n_71), .C(n_72), .Y(n_973) );
BUFx3_ASAP7_75t_L g974 ( .A(n_799), .Y(n_974) );
AO31x2_ASAP7_75t_L g975 ( .A1(n_824), .A2(n_72), .A3(n_73), .B(n_74), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_780), .A2(n_781), .B1(n_818), .B2(n_812), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_810), .A2(n_73), .B1(n_74), .B2(n_75), .Y(n_977) );
BUFx3_ASAP7_75t_L g978 ( .A(n_851), .Y(n_978) );
BUFx12f_ASAP7_75t_L g979 ( .A(n_762), .Y(n_979) );
O2A1O1Ixp33_ASAP7_75t_SL g980 ( .A1(n_846), .A2(n_233), .B(n_360), .C(n_359), .Y(n_980) );
OAI22xp33_ASAP7_75t_L g981 ( .A1(n_827), .A2(n_76), .B1(n_78), .B2(n_79), .Y(n_981) );
OAI21xp5_ASAP7_75t_L g982 ( .A1(n_784), .A2(n_217), .B(n_216), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_825), .Y(n_983) );
INVx1_ASAP7_75t_L g984 ( .A(n_833), .Y(n_984) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_829), .B(n_76), .Y(n_985) );
A2O1A1Ixp33_ASAP7_75t_L g986 ( .A1(n_813), .A2(n_79), .B(n_81), .C(n_83), .Y(n_986) );
INVx2_ASAP7_75t_SL g987 ( .A(n_795), .Y(n_987) );
BUFx6f_ASAP7_75t_L g988 ( .A(n_847), .Y(n_988) );
INVx2_ASAP7_75t_SL g989 ( .A(n_735), .Y(n_989) );
INVxp67_ASAP7_75t_L g990 ( .A(n_824), .Y(n_990) );
INVx2_ASAP7_75t_L g991 ( .A(n_800), .Y(n_991) );
O2A1O1Ixp33_ASAP7_75t_SL g992 ( .A1(n_830), .A2(n_235), .B(n_358), .C(n_357), .Y(n_992) );
AOI21xp5_ASAP7_75t_L g993 ( .A1(n_831), .A2(n_227), .B(n_224), .Y(n_993) );
BUFx6f_ASAP7_75t_L g994 ( .A(n_847), .Y(n_994) );
AOI221x1_ASAP7_75t_L g995 ( .A1(n_813), .A2(n_81), .B1(n_84), .B2(n_85), .C(n_86), .Y(n_995) );
CKINVDCx5p33_ASAP7_75t_R g996 ( .A(n_804), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_762), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_762), .Y(n_998) );
AOI21xp5_ASAP7_75t_L g999 ( .A1(n_845), .A2(n_230), .B(n_228), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_807), .B(n_85), .Y(n_1000) );
INVx2_ASAP7_75t_L g1001 ( .A(n_809), .Y(n_1001) );
AOI221xp5_ASAP7_75t_L g1002 ( .A1(n_832), .A2(n_87), .B1(n_88), .B2(n_89), .C(n_90), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_740), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_735), .B(n_87), .Y(n_1004) );
OAI22x1_ASAP7_75t_L g1005 ( .A1(n_856), .A2(n_89), .B1(n_91), .B2(n_92), .Y(n_1005) );
AO31x2_ASAP7_75t_L g1006 ( .A1(n_828), .A2(n_93), .A3(n_94), .B(n_95), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_858), .B(n_95), .Y(n_1007) );
OAI221xp5_ASAP7_75t_L g1008 ( .A1(n_733), .A2(n_96), .B1(n_97), .B2(n_98), .C(n_99), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_734), .B(n_96), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_861), .Y(n_1010) );
AOI22xp33_ASAP7_75t_SL g1011 ( .A1(n_816), .A2(n_97), .B1(n_99), .B2(n_100), .Y(n_1011) );
AOI21xp5_ASAP7_75t_L g1012 ( .A1(n_819), .A2(n_234), .B(n_232), .Y(n_1012) );
HB1xp67_ASAP7_75t_L g1013 ( .A(n_815), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_862), .Y(n_1014) );
NOR2xp33_ASAP7_75t_L g1015 ( .A(n_866), .B(n_101), .Y(n_1015) );
AOI21xp5_ASAP7_75t_L g1016 ( .A1(n_854), .A2(n_239), .B(n_238), .Y(n_1016) );
INVx2_ASAP7_75t_L g1017 ( .A(n_822), .Y(n_1017) );
AO31x2_ASAP7_75t_L g1018 ( .A1(n_817), .A2(n_101), .A3(n_102), .B(n_103), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_766), .A2(n_102), .B1(n_104), .B2(n_105), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_771), .B(n_104), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_773), .B(n_105), .Y(n_1021) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_775), .A2(n_106), .B1(n_107), .B2(n_108), .Y(n_1022) );
CKINVDCx5p33_ASAP7_75t_R g1023 ( .A(n_826), .Y(n_1023) );
OA21x2_ASAP7_75t_L g1024 ( .A1(n_867), .A2(n_259), .B(n_353), .Y(n_1024) );
AOI21xp5_ASAP7_75t_L g1025 ( .A1(n_867), .A2(n_263), .B(n_351), .Y(n_1025) );
BUFx2_ASAP7_75t_L g1026 ( .A(n_747), .Y(n_1026) );
AOI21x1_ASAP7_75t_L g1027 ( .A1(n_867), .A2(n_257), .B(n_349), .Y(n_1027) );
BUFx3_ASAP7_75t_L g1028 ( .A(n_855), .Y(n_1028) );
BUFx3_ASAP7_75t_L g1029 ( .A(n_855), .Y(n_1029) );
OAI22xp33_ASAP7_75t_L g1030 ( .A1(n_745), .A2(n_109), .B1(n_110), .B2(n_111), .Y(n_1030) );
AOI222xp33_ASAP7_75t_L g1031 ( .A1(n_777), .A2(n_109), .B1(n_110), .B2(n_112), .C1(n_113), .C2(n_114), .Y(n_1031) );
INVx2_ASAP7_75t_L g1032 ( .A(n_756), .Y(n_1032) );
O2A1O1Ixp33_ASAP7_75t_L g1033 ( .A1(n_739), .A2(n_112), .B(n_113), .C(n_115), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_943), .B(n_116), .Y(n_1034) );
BUFx6f_ASAP7_75t_L g1035 ( .A(n_908), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_868), .Y(n_1036) );
AO31x2_ASAP7_75t_L g1037 ( .A1(n_997), .A2(n_118), .A3(n_119), .B(n_120), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_990), .B(n_120), .Y(n_1038) );
AND2x2_ASAP7_75t_SL g1039 ( .A(n_883), .B(n_956), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_909), .B(n_121), .Y(n_1040) );
OR2x6_ASAP7_75t_L g1041 ( .A(n_955), .B(n_121), .Y(n_1041) );
INVx8_ASAP7_75t_L g1042 ( .A(n_901), .Y(n_1042) );
AO31x2_ASAP7_75t_L g1043 ( .A1(n_998), .A2(n_122), .A3(n_123), .B(n_124), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_883), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_967), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_996), .B(n_125), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_983), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_984), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_921), .B(n_126), .Y(n_1049) );
INVxp67_ASAP7_75t_L g1050 ( .A(n_1026), .Y(n_1050) );
AND2x4_ASAP7_75t_L g1051 ( .A(n_901), .B(n_126), .Y(n_1051) );
OR2x2_ASAP7_75t_L g1052 ( .A(n_893), .B(n_127), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_872), .Y(n_1053) );
AOI21xp5_ASAP7_75t_L g1054 ( .A1(n_873), .A2(n_274), .B(n_347), .Y(n_1054) );
AOI21xp5_ASAP7_75t_L g1055 ( .A1(n_870), .A2(n_271), .B(n_345), .Y(n_1055) );
INVx2_ASAP7_75t_L g1056 ( .A(n_964), .Y(n_1056) );
OAI21xp5_ASAP7_75t_L g1057 ( .A1(n_913), .A2(n_127), .B(n_128), .Y(n_1057) );
OAI21x1_ASAP7_75t_L g1058 ( .A1(n_903), .A2(n_890), .B(n_1027), .Y(n_1058) );
AOI21xp5_ASAP7_75t_L g1059 ( .A1(n_874), .A2(n_270), .B(n_344), .Y(n_1059) );
NOR2xp33_ASAP7_75t_L g1060 ( .A(n_885), .B(n_128), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_960), .Y(n_1061) );
INVx8_ASAP7_75t_L g1062 ( .A(n_901), .Y(n_1062) );
A2O1A1Ixp33_ASAP7_75t_L g1063 ( .A1(n_947), .A2(n_129), .B(n_130), .C(n_131), .Y(n_1063) );
OAI21xp5_ASAP7_75t_SL g1064 ( .A1(n_944), .A2(n_129), .B(n_132), .Y(n_1064) );
OAI22xp33_ASAP7_75t_L g1065 ( .A1(n_922), .A2(n_133), .B1(n_135), .B2(n_136), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_926), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_878), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_920), .B(n_133), .Y(n_1068) );
AOI221xp5_ASAP7_75t_L g1069 ( .A1(n_963), .A2(n_137), .B1(n_138), .B2(n_139), .C(n_140), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_956), .B(n_139), .Y(n_1070) );
OAI21xp5_ASAP7_75t_L g1071 ( .A1(n_907), .A2(n_140), .B(n_141), .Y(n_1071) );
INVx2_ASAP7_75t_L g1072 ( .A(n_969), .Y(n_1072) );
OAI21x1_ASAP7_75t_SL g1073 ( .A1(n_941), .A2(n_142), .B(n_143), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_892), .Y(n_1074) );
AO21x2_ASAP7_75t_L g1075 ( .A1(n_884), .A2(n_288), .B(n_343), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_894), .B(n_143), .Y(n_1076) );
CKINVDCx9p33_ASAP7_75t_R g1077 ( .A(n_888), .Y(n_1077) );
INVx1_ASAP7_75t_SL g1078 ( .A(n_978), .Y(n_1078) );
AO31x2_ASAP7_75t_L g1079 ( .A1(n_1025), .A2(n_995), .A3(n_1016), .B(n_886), .Y(n_1079) );
CKINVDCx5p33_ASAP7_75t_R g1080 ( .A(n_898), .Y(n_1080) );
INVx2_ASAP7_75t_L g1081 ( .A(n_991), .Y(n_1081) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_930), .B(n_144), .Y(n_1082) );
OAI21xp5_ASAP7_75t_L g1083 ( .A1(n_1009), .A2(n_144), .B(n_145), .Y(n_1083) );
OAI21x1_ASAP7_75t_L g1084 ( .A1(n_910), .A2(n_282), .B(n_340), .Y(n_1084) );
AND2x4_ASAP7_75t_L g1085 ( .A(n_941), .B(n_145), .Y(n_1085) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_979), .A2(n_146), .B1(n_147), .B2(n_148), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_958), .B(n_148), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_959), .Y(n_1088) );
AOI22xp5_ASAP7_75t_L g1089 ( .A1(n_889), .A2(n_149), .B1(n_150), .B2(n_151), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1005), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_976), .B(n_150), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_879), .B(n_151), .Y(n_1092) );
AOI221xp5_ASAP7_75t_L g1093 ( .A1(n_1030), .A2(n_152), .B1(n_153), .B2(n_154), .C(n_155), .Y(n_1093) );
A2O1A1Ixp33_ASAP7_75t_L g1094 ( .A1(n_985), .A2(n_152), .B(n_153), .C(n_154), .Y(n_1094) );
INVx3_ASAP7_75t_L g1095 ( .A(n_908), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_954), .B(n_242), .Y(n_1096) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1001), .Y(n_1097) );
AOI21xp5_ASAP7_75t_L g1098 ( .A1(n_1000), .A2(n_243), .B(n_245), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_938), .B(n_361), .Y(n_1099) );
INVx3_ASAP7_75t_L g1100 ( .A(n_908), .Y(n_1100) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1003), .Y(n_1101) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_891), .B(n_246), .Y(n_1102) );
BUFx3_ASAP7_75t_L g1103 ( .A(n_1028), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_952), .A2(n_247), .B1(n_248), .B2(n_250), .Y(n_1104) );
BUFx6f_ASAP7_75t_SL g1105 ( .A(n_1029), .Y(n_1105) );
OR2x2_ASAP7_75t_L g1106 ( .A(n_965), .B(n_252), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_932), .B(n_338), .Y(n_1107) );
INVx2_ASAP7_75t_L g1108 ( .A(n_1007), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_975), .Y(n_1109) );
BUFx3_ASAP7_75t_L g1110 ( .A(n_942), .Y(n_1110) );
AO21x2_ASAP7_75t_L g1111 ( .A1(n_925), .A2(n_253), .B(n_266), .Y(n_1111) );
OR2x6_ASAP7_75t_L g1112 ( .A(n_900), .B(n_268), .Y(n_1112) );
INVx2_ASAP7_75t_L g1113 ( .A(n_1010), .Y(n_1113) );
BUFx2_ASAP7_75t_L g1114 ( .A(n_900), .Y(n_1114) );
INVx1_ASAP7_75t_L g1115 ( .A(n_975), .Y(n_1115) );
CKINVDCx20_ASAP7_75t_R g1116 ( .A(n_914), .Y(n_1116) );
INVx2_ASAP7_75t_L g1117 ( .A(n_1014), .Y(n_1117) );
NOR2xp33_ASAP7_75t_L g1118 ( .A(n_927), .B(n_269), .Y(n_1118) );
AO31x2_ASAP7_75t_L g1119 ( .A1(n_902), .A2(n_277), .A3(n_278), .B(n_280), .Y(n_1119) );
AO21x2_ASAP7_75t_L g1120 ( .A1(n_970), .A2(n_281), .B(n_294), .Y(n_1120) );
BUFx8_ASAP7_75t_L g1121 ( .A(n_916), .Y(n_1121) );
INVx2_ASAP7_75t_L g1122 ( .A(n_935), .Y(n_1122) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_880), .A2(n_301), .B1(n_302), .B2(n_303), .Y(n_1123) );
INVx1_ASAP7_75t_SL g1124 ( .A(n_906), .Y(n_1124) );
O2A1O1Ixp33_ASAP7_75t_L g1125 ( .A1(n_897), .A2(n_306), .B(n_308), .C(n_309), .Y(n_1125) );
OAI22xp33_ASAP7_75t_L g1126 ( .A1(n_950), .A2(n_929), .B1(n_923), .B2(n_961), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_975), .Y(n_1127) );
BUFx2_ASAP7_75t_L g1128 ( .A(n_916), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1031), .B(n_313), .Y(n_1129) );
AOI22xp33_ASAP7_75t_SL g1130 ( .A1(n_916), .A2(n_322), .B1(n_324), .B2(n_325), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_962), .A2(n_326), .B1(n_328), .B2(n_331), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_931), .B(n_939), .Y(n_1132) );
AND2x4_ASAP7_75t_L g1133 ( .A(n_871), .B(n_334), .Y(n_1133) );
BUFx6f_ASAP7_75t_L g1134 ( .A(n_935), .Y(n_1134) );
BUFx2_ASAP7_75t_L g1135 ( .A(n_916), .Y(n_1135) );
OR2x6_ASAP7_75t_L g1136 ( .A(n_931), .B(n_335), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_928), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_928), .Y(n_1138) );
AND2x4_ASAP7_75t_L g1139 ( .A(n_871), .B(n_337), .Y(n_1139) );
INVx2_ASAP7_75t_L g1140 ( .A(n_935), .Y(n_1140) );
OAI221xp5_ASAP7_75t_SL g1141 ( .A1(n_934), .A2(n_1033), .B1(n_899), .B2(n_918), .C(n_875), .Y(n_1141) );
A2O1A1Ixp33_ASAP7_75t_L g1142 ( .A1(n_911), .A2(n_915), .B(n_1015), .C(n_948), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_939), .B(n_987), .Y(n_1143) );
OAI21x1_ASAP7_75t_L g1144 ( .A1(n_917), .A2(n_937), .B(n_1024), .Y(n_1144) );
AOI21xp5_ASAP7_75t_L g1145 ( .A1(n_1024), .A2(n_980), .B(n_951), .Y(n_1145) );
A2O1A1Ixp33_ASAP7_75t_L g1146 ( .A1(n_986), .A2(n_1021), .B(n_1020), .C(n_945), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_936), .B(n_946), .Y(n_1147) );
NOR2x1_ASAP7_75t_SL g1148 ( .A(n_966), .B(n_988), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_887), .B(n_1032), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_896), .B(n_876), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_928), .Y(n_1151) );
AOI21xp5_ASAP7_75t_L g1152 ( .A1(n_971), .A2(n_982), .B(n_992), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1023), .B(n_877), .Y(n_1153) );
NAND2x1p5_ASAP7_75t_L g1154 ( .A(n_966), .B(n_974), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_968), .Y(n_1155) );
AOI222xp33_ASAP7_75t_L g1156 ( .A1(n_914), .A2(n_1002), .B1(n_1008), .B2(n_1022), .C1(n_981), .C2(n_977), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1017), .B(n_989), .Y(n_1157) );
BUFx8_ASAP7_75t_L g1158 ( .A(n_912), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1004), .B(n_1011), .Y(n_1159) );
OA21x2_ASAP7_75t_L g1160 ( .A1(n_957), .A2(n_972), .B(n_993), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g1161 ( .A1(n_919), .A2(n_1013), .B1(n_895), .B2(n_1019), .Y(n_1161) );
INVx2_ASAP7_75t_L g1162 ( .A(n_905), .Y(n_1162) );
CKINVDCx5p33_ASAP7_75t_R g1163 ( .A(n_924), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_973), .B(n_968), .Y(n_1164) );
INVx2_ASAP7_75t_L g1165 ( .A(n_905), .Y(n_1165) );
OAI21xp5_ASAP7_75t_L g1166 ( .A1(n_1012), .A2(n_949), .B(n_999), .Y(n_1166) );
OA21x2_ASAP7_75t_L g1167 ( .A1(n_933), .A2(n_895), .B(n_1018), .Y(n_1167) );
INVx1_ASAP7_75t_L g1168 ( .A(n_933), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_933), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_895), .B(n_1006), .Y(n_1170) );
BUFx3_ASAP7_75t_L g1171 ( .A(n_904), .Y(n_1171) );
AOI221xp5_ASAP7_75t_L g1172 ( .A1(n_940), .A2(n_988), .B1(n_994), .B2(n_912), .C(n_953), .Y(n_1172) );
OA21x2_ASAP7_75t_L g1173 ( .A1(n_1018), .A2(n_953), .B(n_912), .Y(n_1173) );
INVx5_ASAP7_75t_L g1174 ( .A(n_904), .Y(n_1174) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_953), .A2(n_1006), .B1(n_1018), .B2(n_904), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1006), .Y(n_1176) );
INVx2_ASAP7_75t_L g1177 ( .A(n_904), .Y(n_1177) );
A2O1A1Ixp33_ASAP7_75t_L g1178 ( .A1(n_947), .A2(n_889), .B(n_985), .C(n_646), .Y(n_1178) );
CKINVDCx11_ASAP7_75t_R g1179 ( .A(n_1028), .Y(n_1179) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_889), .A2(n_675), .B1(n_673), .B2(n_753), .Y(n_1180) );
AOI21xp5_ASAP7_75t_L g1181 ( .A1(n_873), .A2(n_870), .B(n_869), .Y(n_1181) );
AND2x4_ASAP7_75t_L g1182 ( .A(n_901), .B(n_941), .Y(n_1182) );
BUFx2_ASAP7_75t_L g1183 ( .A(n_1026), .Y(n_1183) );
A2O1A1Ixp33_ASAP7_75t_L g1184 ( .A1(n_947), .A2(n_889), .B(n_985), .C(n_646), .Y(n_1184) );
AOI21xp5_ASAP7_75t_L g1185 ( .A1(n_873), .A2(n_870), .B(n_869), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_909), .B(n_748), .Y(n_1186) );
AO31x2_ASAP7_75t_L g1187 ( .A1(n_997), .A2(n_998), .A3(n_761), .B(n_882), .Y(n_1187) );
NOR2xp33_ASAP7_75t_L g1188 ( .A(n_996), .B(n_760), .Y(n_1188) );
INVx2_ASAP7_75t_L g1189 ( .A(n_967), .Y(n_1189) );
BUFx12f_ASAP7_75t_L g1190 ( .A(n_898), .Y(n_1190) );
AO21x2_ASAP7_75t_L g1191 ( .A1(n_997), .A2(n_998), .B(n_881), .Y(n_1191) );
NOR2x1_ASAP7_75t_SL g1192 ( .A(n_901), .B(n_787), .Y(n_1192) );
NOR2xp33_ASAP7_75t_L g1193 ( .A(n_996), .B(n_760), .Y(n_1193) );
OAI21x1_ASAP7_75t_L g1194 ( .A1(n_903), .A2(n_870), .B(n_869), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_868), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_909), .B(n_748), .Y(n_1196) );
OA21x2_ASAP7_75t_L g1197 ( .A1(n_1181), .A2(n_1185), .B(n_1162), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1176), .Y(n_1198) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1189), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1109), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1036), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1195), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1115), .Y(n_1203) );
AOI21x1_ASAP7_75t_L g1204 ( .A1(n_1170), .A2(n_1175), .B(n_1164), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1045), .Y(n_1205) );
OR2x6_ASAP7_75t_L g1206 ( .A(n_1136), .B(n_1128), .Y(n_1206) );
BUFx2_ASAP7_75t_L g1207 ( .A(n_1135), .Y(n_1207) );
BUFx3_ASAP7_75t_L g1208 ( .A(n_1182), .Y(n_1208) );
INVx2_ASAP7_75t_L g1209 ( .A(n_1165), .Y(n_1209) );
AO21x2_ASAP7_75t_L g1210 ( .A1(n_1175), .A2(n_1138), .B(n_1137), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1047), .Y(n_1211) );
HB1xp67_ASAP7_75t_L g1212 ( .A(n_1183), .Y(n_1212) );
OAI21x1_ASAP7_75t_L g1213 ( .A1(n_1058), .A2(n_1194), .B(n_1144), .Y(n_1213) );
INVxp67_ASAP7_75t_L g1214 ( .A(n_1052), .Y(n_1214) );
NAND4xp25_ASAP7_75t_L g1215 ( .A(n_1180), .B(n_1090), .C(n_1064), .D(n_1088), .Y(n_1215) );
OA21x2_ASAP7_75t_L g1216 ( .A1(n_1168), .A2(n_1169), .B(n_1151), .Y(n_1216) );
INVx3_ASAP7_75t_SL g1217 ( .A(n_1116), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1127), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1056), .B(n_1072), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1155), .Y(n_1220) );
INVx3_ASAP7_75t_L g1221 ( .A(n_1174), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1048), .Y(n_1222) );
OR2x2_ASAP7_75t_L g1223 ( .A(n_1124), .B(n_1196), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1101), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1081), .B(n_1097), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1173), .Y(n_1226) );
HB1xp67_ASAP7_75t_L g1227 ( .A(n_1041), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1173), .Y(n_1228) );
AO21x2_ASAP7_75t_L g1229 ( .A1(n_1191), .A2(n_1057), .B(n_1071), .Y(n_1229) );
AO21x2_ASAP7_75t_L g1230 ( .A1(n_1071), .A2(n_1142), .B(n_1146), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1037), .Y(n_1231) );
OR2x2_ASAP7_75t_L g1232 ( .A(n_1124), .B(n_1034), .Y(n_1232) );
INVx2_ASAP7_75t_L g1233 ( .A(n_1187), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1037), .Y(n_1234) );
INVx2_ASAP7_75t_L g1235 ( .A(n_1187), .Y(n_1235) );
INVx2_ASAP7_75t_L g1236 ( .A(n_1187), .Y(n_1236) );
HB1xp67_ASAP7_75t_L g1237 ( .A(n_1041), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1037), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1043), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1039), .B(n_1113), .Y(n_1240) );
AOI221xp5_ASAP7_75t_L g1241 ( .A1(n_1065), .A2(n_1064), .B1(n_1126), .B2(n_1053), .C(n_1069), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1117), .B(n_1147), .Y(n_1242) );
INVx1_ASAP7_75t_SL g1243 ( .A(n_1078), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1043), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1245 ( .A(n_1034), .B(n_1038), .Y(n_1245) );
OA21x2_ASAP7_75t_L g1246 ( .A1(n_1172), .A2(n_1166), .B(n_1084), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1083), .B(n_1067), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1186), .B(n_1061), .Y(n_1248) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1074), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1149), .Y(n_1250) );
AO21x2_ASAP7_75t_L g1251 ( .A1(n_1120), .A2(n_1111), .B(n_1184), .Y(n_1251) );
OR2x6_ASAP7_75t_L g1252 ( .A(n_1136), .B(n_1112), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1108), .B(n_1136), .Y(n_1253) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1134), .Y(n_1254) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1085), .Y(n_1255) );
INVxp67_ASAP7_75t_SL g1256 ( .A(n_1121), .Y(n_1256) );
OR2x6_ASAP7_75t_L g1257 ( .A(n_1112), .B(n_1042), .Y(n_1257) );
INVx2_ASAP7_75t_SL g1258 ( .A(n_1042), .Y(n_1258) );
INVx3_ASAP7_75t_L g1259 ( .A(n_1174), .Y(n_1259) );
AND2x4_ASAP7_75t_L g1260 ( .A(n_1182), .B(n_1174), .Y(n_1260) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1085), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1262 ( .A(n_1044), .B(n_1159), .Y(n_1262) );
INVx2_ASAP7_75t_L g1263 ( .A(n_1134), .Y(n_1263) );
OAI33xp33_ASAP7_75t_L g1264 ( .A1(n_1086), .A2(n_1087), .A3(n_1091), .B1(n_1046), .B2(n_1076), .B3(n_1082), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1043), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1167), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1041), .B(n_1049), .Y(n_1267) );
INVx3_ASAP7_75t_L g1268 ( .A(n_1171), .Y(n_1268) );
BUFx2_ASAP7_75t_L g1269 ( .A(n_1121), .Y(n_1269) );
OA21x2_ASAP7_75t_L g1270 ( .A1(n_1054), .A2(n_1055), .B(n_1059), .Y(n_1270) );
OAI22xp5_ASAP7_75t_L g1271 ( .A1(n_1112), .A2(n_1089), .B1(n_1114), .B2(n_1178), .Y(n_1271) );
OA21x2_ASAP7_75t_L g1272 ( .A1(n_1107), .A2(n_1098), .B(n_1131), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1188), .B(n_1193), .Y(n_1273) );
BUFx3_ASAP7_75t_L g1274 ( .A(n_1042), .Y(n_1274) );
OR2x6_ASAP7_75t_L g1275 ( .A(n_1062), .B(n_1051), .Y(n_1275) );
BUFx3_ASAP7_75t_L g1276 ( .A(n_1062), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1051), .Y(n_1277) );
BUFx3_ASAP7_75t_L g1278 ( .A(n_1062), .Y(n_1278) );
OR2x2_ASAP7_75t_L g1279 ( .A(n_1078), .B(n_1050), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1167), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1281 ( .A(n_1129), .B(n_1068), .Y(n_1281) );
AND2x4_ASAP7_75t_L g1282 ( .A(n_1066), .B(n_1100), .Y(n_1282) );
AND2x4_ASAP7_75t_L g1283 ( .A(n_1095), .B(n_1100), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1070), .B(n_1086), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1158), .Y(n_1285) );
INVx2_ASAP7_75t_L g1286 ( .A(n_1035), .Y(n_1286) );
INVx1_ASAP7_75t_SL g1287 ( .A(n_1103), .Y(n_1287) );
INVx2_ASAP7_75t_L g1288 ( .A(n_1035), .Y(n_1288) );
OA21x2_ASAP7_75t_L g1289 ( .A1(n_1150), .A2(n_1094), .B(n_1063), .Y(n_1289) );
AND2x4_ASAP7_75t_L g1290 ( .A(n_1095), .B(n_1148), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1133), .B(n_1139), .Y(n_1291) );
OR2x2_ASAP7_75t_L g1292 ( .A(n_1102), .B(n_1153), .Y(n_1292) );
OR2x2_ASAP7_75t_L g1293 ( .A(n_1132), .B(n_1157), .Y(n_1293) );
INVxp67_ASAP7_75t_SL g1294 ( .A(n_1192), .Y(n_1294) );
OR2x2_ASAP7_75t_L g1295 ( .A(n_1143), .B(n_1154), .Y(n_1295) );
OAI221xp5_ASAP7_75t_L g1296 ( .A1(n_1141), .A2(n_1060), .B1(n_1161), .B2(n_1093), .C(n_1156), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1133), .B(n_1139), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1040), .B(n_1122), .Y(n_1298) );
AO21x2_ASAP7_75t_L g1299 ( .A1(n_1075), .A2(n_1073), .B(n_1125), .Y(n_1299) );
OAI21xp5_ASAP7_75t_L g1300 ( .A1(n_1156), .A2(n_1104), .B(n_1123), .Y(n_1300) );
INVx2_ASAP7_75t_L g1301 ( .A(n_1035), .Y(n_1301) );
INVx2_ASAP7_75t_L g1302 ( .A(n_1140), .Y(n_1302) );
AOI22xp33_ASAP7_75t_L g1303 ( .A1(n_1158), .A2(n_1092), .B1(n_1099), .B2(n_1118), .Y(n_1303) );
OAI22xp5_ASAP7_75t_L g1304 ( .A1(n_1130), .A2(n_1123), .B1(n_1096), .B2(n_1077), .Y(n_1304) );
AO21x2_ASAP7_75t_L g1305 ( .A1(n_1075), .A2(n_1177), .B(n_1079), .Y(n_1305) );
INVx2_ASAP7_75t_L g1306 ( .A(n_1119), .Y(n_1306) );
OA21x2_ASAP7_75t_L g1307 ( .A1(n_1079), .A2(n_1119), .B(n_1160), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1106), .B(n_1110), .Y(n_1308) );
OA21x2_ASAP7_75t_L g1309 ( .A1(n_1080), .A2(n_1163), .B(n_1105), .Y(n_1309) );
HB1xp67_ASAP7_75t_L g1310 ( .A(n_1105), .Y(n_1310) );
OAI21xp5_ASAP7_75t_L g1311 ( .A1(n_1179), .A2(n_1184), .B(n_1178), .Y(n_1311) );
AOI21xp5_ASAP7_75t_L g1312 ( .A1(n_1190), .A2(n_1152), .B(n_1145), .Y(n_1312) );
INVx3_ASAP7_75t_L g1313 ( .A(n_1174), .Y(n_1313) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_1186), .B(n_990), .Y(n_1314) );
AO21x2_ASAP7_75t_L g1315 ( .A1(n_1181), .A2(n_1185), .B(n_1170), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g1316 ( .A1(n_1129), .A2(n_753), .B1(n_1180), .B2(n_889), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1056), .B(n_1072), .Y(n_1317) );
INVxp67_ASAP7_75t_L g1318 ( .A(n_1183), .Y(n_1318) );
OR2x6_ASAP7_75t_L g1319 ( .A(n_1136), .B(n_1128), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1176), .Y(n_1320) );
BUFx3_ASAP7_75t_L g1321 ( .A(n_1182), .Y(n_1321) );
INVx3_ASAP7_75t_L g1322 ( .A(n_1174), .Y(n_1322) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1176), .Y(n_1323) );
AND2x4_ASAP7_75t_L g1324 ( .A(n_1252), .B(n_1285), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1242), .B(n_1199), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1242), .B(n_1199), .Y(n_1326) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1198), .Y(n_1327) );
AOI22xp33_ASAP7_75t_L g1328 ( .A1(n_1296), .A2(n_1252), .B1(n_1271), .B2(n_1311), .Y(n_1328) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1198), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1200), .B(n_1203), .Y(n_1330) );
AND2x4_ASAP7_75t_L g1331 ( .A(n_1252), .B(n_1285), .Y(n_1331) );
NOR2xp33_ASAP7_75t_L g1332 ( .A(n_1273), .B(n_1215), .Y(n_1332) );
NAND2xp5_ASAP7_75t_SL g1333 ( .A(n_1304), .B(n_1291), .Y(n_1333) );
OR2x6_ASAP7_75t_L g1334 ( .A(n_1252), .B(n_1206), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1200), .B(n_1203), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1218), .B(n_1220), .Y(n_1336) );
NOR2xp33_ASAP7_75t_L g1337 ( .A(n_1292), .B(n_1287), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1218), .B(n_1220), .Y(n_1338) );
BUFx3_ASAP7_75t_L g1339 ( .A(n_1274), .Y(n_1339) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1320), .Y(n_1340) );
NAND2xp5_ASAP7_75t_L g1341 ( .A(n_1314), .B(n_1250), .Y(n_1341) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_1201), .B(n_1202), .Y(n_1342) );
AND2x4_ASAP7_75t_L g1343 ( .A(n_1206), .B(n_1319), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1320), .B(n_1323), .Y(n_1344) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1323), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1205), .B(n_1211), .Y(n_1346) );
HB1xp67_ASAP7_75t_L g1347 ( .A(n_1293), .Y(n_1347) );
NOR2x1_ASAP7_75t_R g1348 ( .A(n_1269), .B(n_1256), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1222), .B(n_1224), .Y(n_1349) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1216), .Y(n_1350) );
INVxp67_ASAP7_75t_R g1351 ( .A(n_1291), .Y(n_1351) );
BUFx3_ASAP7_75t_L g1352 ( .A(n_1274), .Y(n_1352) );
NAND2xp5_ASAP7_75t_L g1353 ( .A(n_1219), .B(n_1225), .Y(n_1353) );
BUFx6f_ASAP7_75t_L g1354 ( .A(n_1213), .Y(n_1354) );
HB1xp67_ASAP7_75t_L g1355 ( .A(n_1293), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_1219), .B(n_1225), .Y(n_1356) );
NOR2xp33_ASAP7_75t_L g1357 ( .A(n_1292), .B(n_1248), .Y(n_1357) );
NAND2xp5_ASAP7_75t_L g1358 ( .A(n_1317), .B(n_1223), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1317), .B(n_1247), .Y(n_1359) );
AND2x4_ASAP7_75t_L g1360 ( .A(n_1206), .B(n_1319), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1223), .B(n_1284), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1247), .B(n_1230), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1284), .B(n_1249), .Y(n_1363) );
BUFx3_ASAP7_75t_L g1364 ( .A(n_1276), .Y(n_1364) );
NAND2xp5_ASAP7_75t_L g1365 ( .A(n_1240), .B(n_1298), .Y(n_1365) );
AND2x4_ASAP7_75t_L g1366 ( .A(n_1206), .B(n_1319), .Y(n_1366) );
OR2x2_ASAP7_75t_L g1367 ( .A(n_1232), .B(n_1262), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1230), .B(n_1210), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1230), .B(n_1210), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1240), .B(n_1298), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1210), .B(n_1231), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1372 ( .A(n_1262), .B(n_1214), .Y(n_1372) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1226), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1226), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1231), .B(n_1234), .Y(n_1375) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1228), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_1234), .B(n_1238), .Y(n_1377) );
INVxp67_ASAP7_75t_SL g1378 ( .A(n_1297), .Y(n_1378) );
AND2x4_ASAP7_75t_L g1379 ( .A(n_1319), .B(n_1257), .Y(n_1379) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1228), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1238), .B(n_1239), .Y(n_1381) );
NAND2xp5_ASAP7_75t_L g1382 ( .A(n_1267), .B(n_1241), .Y(n_1382) );
AND2x2_ASAP7_75t_L g1383 ( .A(n_1239), .B(n_1244), .Y(n_1383) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1244), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1265), .B(n_1302), .Y(n_1385) );
BUFx3_ASAP7_75t_L g1386 ( .A(n_1276), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1302), .B(n_1209), .Y(n_1387) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1266), .Y(n_1388) );
INVx2_ASAP7_75t_SL g1389 ( .A(n_1260), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1266), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1280), .Y(n_1391) );
INVx2_ASAP7_75t_L g1392 ( .A(n_1280), .Y(n_1392) );
OR2x2_ASAP7_75t_L g1393 ( .A(n_1232), .B(n_1245), .Y(n_1393) );
INVx5_ASAP7_75t_L g1394 ( .A(n_1257), .Y(n_1394) );
OR2x2_ASAP7_75t_L g1395 ( .A(n_1245), .B(n_1257), .Y(n_1395) );
OR2x2_ASAP7_75t_L g1396 ( .A(n_1257), .B(n_1297), .Y(n_1396) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1204), .B(n_1315), .Y(n_1397) );
INVx2_ASAP7_75t_SL g1398 ( .A(n_1260), .Y(n_1398) );
INVx2_ASAP7_75t_SL g1399 ( .A(n_1260), .Y(n_1399) );
INVx4_ASAP7_75t_L g1400 ( .A(n_1275), .Y(n_1400) );
NAND2xp33_ASAP7_75t_SL g1401 ( .A(n_1269), .B(n_1227), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1204), .B(n_1315), .Y(n_1402) );
NAND2xp5_ASAP7_75t_L g1403 ( .A(n_1267), .B(n_1253), .Y(n_1403) );
HB1xp67_ASAP7_75t_L g1404 ( .A(n_1212), .Y(n_1404) );
NAND2xp5_ASAP7_75t_SL g1405 ( .A(n_1294), .B(n_1290), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1253), .B(n_1243), .Y(n_1406) );
HB1xp67_ASAP7_75t_L g1407 ( .A(n_1347), .Y(n_1407) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1355), .Y(n_1408) );
NAND2xp5_ASAP7_75t_L g1409 ( .A(n_1325), .B(n_1237), .Y(n_1409) );
OR2x2_ASAP7_75t_L g1410 ( .A(n_1393), .B(n_1361), .Y(n_1410) );
HB1xp67_ASAP7_75t_L g1411 ( .A(n_1404), .Y(n_1411) );
AND2x2_ASAP7_75t_L g1412 ( .A(n_1359), .B(n_1315), .Y(n_1412) );
INVx2_ASAP7_75t_L g1413 ( .A(n_1392), .Y(n_1413) );
OR2x2_ASAP7_75t_L g1414 ( .A(n_1393), .B(n_1279), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1415 ( .A(n_1325), .B(n_1318), .Y(n_1415) );
INVx3_ASAP7_75t_SL g1416 ( .A(n_1339), .Y(n_1416) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1342), .Y(n_1417) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1346), .Y(n_1418) );
NAND2xp5_ASAP7_75t_L g1419 ( .A(n_1326), .B(n_1255), .Y(n_1419) );
AND2x2_ASAP7_75t_L g1420 ( .A(n_1359), .B(n_1362), .Y(n_1420) );
NAND4xp25_ASAP7_75t_SL g1421 ( .A(n_1348), .B(n_1316), .C(n_1303), .D(n_1308), .Y(n_1421) );
NAND2xp5_ASAP7_75t_L g1422 ( .A(n_1326), .B(n_1261), .Y(n_1422) );
INVxp67_ASAP7_75t_L g1423 ( .A(n_1348), .Y(n_1423) );
HB1xp67_ASAP7_75t_L g1424 ( .A(n_1356), .Y(n_1424) );
INVx2_ASAP7_75t_L g1425 ( .A(n_1392), .Y(n_1425) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_1362), .B(n_1197), .Y(n_1426) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1349), .Y(n_1427) );
AND2x4_ASAP7_75t_SL g1428 ( .A(n_1400), .B(n_1275), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1330), .B(n_1197), .Y(n_1429) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1327), .Y(n_1430) );
OR2x2_ASAP7_75t_L g1431 ( .A(n_1367), .B(n_1279), .Y(n_1431) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1327), .Y(n_1432) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1330), .B(n_1197), .Y(n_1433) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1329), .Y(n_1434) );
NAND2x1_ASAP7_75t_SL g1435 ( .A(n_1379), .B(n_1217), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1335), .B(n_1197), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_1356), .B(n_1277), .Y(n_1437) );
OAI221xp5_ASAP7_75t_L g1438 ( .A1(n_1328), .A2(n_1332), .B1(n_1382), .B2(n_1281), .C(n_1333), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_1358), .B(n_1308), .Y(n_1439) );
OR2x2_ASAP7_75t_L g1440 ( .A(n_1367), .B(n_1235), .Y(n_1440) );
AND2x4_ASAP7_75t_L g1441 ( .A(n_1334), .B(n_1312), .Y(n_1441) );
OR2x2_ASAP7_75t_L g1442 ( .A(n_1403), .B(n_1207), .Y(n_1442) );
OR2x2_ASAP7_75t_L g1443 ( .A(n_1365), .B(n_1207), .Y(n_1443) );
NAND2x1_ASAP7_75t_SL g1444 ( .A(n_1379), .B(n_1217), .Y(n_1444) );
NOR2xp33_ASAP7_75t_L g1445 ( .A(n_1395), .B(n_1264), .Y(n_1445) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_1341), .B(n_1208), .Y(n_1446) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1329), .Y(n_1447) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1340), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1336), .B(n_1236), .Y(n_1449) );
OR2x2_ASAP7_75t_L g1450 ( .A(n_1370), .B(n_1295), .Y(n_1450) );
NAND2xp5_ASAP7_75t_L g1451 ( .A(n_1353), .B(n_1208), .Y(n_1451) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_1336), .B(n_1235), .Y(n_1452) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1338), .B(n_1233), .Y(n_1453) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1340), .Y(n_1454) );
OR2x2_ASAP7_75t_L g1455 ( .A(n_1363), .B(n_1229), .Y(n_1455) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_1338), .B(n_1307), .Y(n_1456) );
NAND2xp5_ASAP7_75t_L g1457 ( .A(n_1357), .B(n_1321), .Y(n_1457) );
OR2x2_ASAP7_75t_L g1458 ( .A(n_1372), .B(n_1229), .Y(n_1458) );
NAND2xp5_ASAP7_75t_L g1459 ( .A(n_1378), .B(n_1321), .Y(n_1459) );
AND2x2_ASAP7_75t_L g1460 ( .A(n_1344), .B(n_1307), .Y(n_1460) );
AND2x2_ASAP7_75t_L g1461 ( .A(n_1344), .B(n_1307), .Y(n_1461) );
BUFx2_ASAP7_75t_L g1462 ( .A(n_1339), .Y(n_1462) );
OR2x2_ASAP7_75t_L g1463 ( .A(n_1395), .B(n_1229), .Y(n_1463) );
HB1xp67_ASAP7_75t_L g1464 ( .A(n_1387), .Y(n_1464) );
OR2x2_ASAP7_75t_L g1465 ( .A(n_1406), .B(n_1295), .Y(n_1465) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1345), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1467 ( .A(n_1368), .B(n_1307), .Y(n_1467) );
NOR2x1_ASAP7_75t_L g1468 ( .A(n_1352), .B(n_1275), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1368), .B(n_1306), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1369), .B(n_1306), .Y(n_1470) );
NAND2xp5_ASAP7_75t_L g1471 ( .A(n_1337), .B(n_1289), .Y(n_1471) );
INVx1_ASAP7_75t_SL g1472 ( .A(n_1352), .Y(n_1472) );
AOI22xp33_ASAP7_75t_L g1473 ( .A1(n_1334), .A2(n_1300), .B1(n_1289), .B2(n_1275), .Y(n_1473) );
NOR2x1p5_ASAP7_75t_L g1474 ( .A(n_1364), .B(n_1278), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_1369), .B(n_1305), .Y(n_1475) );
INVx1_ASAP7_75t_SL g1476 ( .A(n_1364), .Y(n_1476) );
NAND2xp5_ASAP7_75t_L g1477 ( .A(n_1345), .B(n_1324), .Y(n_1477) );
HB1xp67_ASAP7_75t_L g1478 ( .A(n_1387), .Y(n_1478) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_1385), .B(n_1305), .Y(n_1479) );
AND2x4_ASAP7_75t_L g1480 ( .A(n_1334), .B(n_1305), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1481 ( .A(n_1385), .B(n_1246), .Y(n_1481) );
NAND2xp5_ASAP7_75t_L g1482 ( .A(n_1324), .B(n_1289), .Y(n_1482) );
AND2x4_ASAP7_75t_SL g1483 ( .A(n_1400), .B(n_1322), .Y(n_1483) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1373), .Y(n_1484) );
INVxp67_ASAP7_75t_L g1485 ( .A(n_1386), .Y(n_1485) );
OR2x2_ASAP7_75t_L g1486 ( .A(n_1396), .B(n_1258), .Y(n_1486) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1373), .Y(n_1487) );
NAND2xp5_ASAP7_75t_L g1488 ( .A(n_1324), .B(n_1289), .Y(n_1488) );
AND4x1_ASAP7_75t_L g1489 ( .A(n_1394), .B(n_1309), .C(n_1278), .D(n_1310), .Y(n_1489) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1420), .B(n_1371), .Y(n_1490) );
AND2x4_ASAP7_75t_L g1491 ( .A(n_1480), .B(n_1343), .Y(n_1491) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1424), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1420), .B(n_1371), .Y(n_1493) );
INVx2_ASAP7_75t_SL g1494 ( .A(n_1474), .Y(n_1494) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1430), .Y(n_1495) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_1412), .B(n_1375), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1497 ( .A(n_1464), .B(n_1374), .Y(n_1497) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1407), .Y(n_1498) );
NAND2xp5_ASAP7_75t_L g1499 ( .A(n_1408), .B(n_1331), .Y(n_1499) );
NAND2xp5_ASAP7_75t_L g1500 ( .A(n_1445), .B(n_1331), .Y(n_1500) );
NOR2x1p5_ASAP7_75t_L g1501 ( .A(n_1471), .B(n_1386), .Y(n_1501) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1411), .Y(n_1502) );
OR2x2_ASAP7_75t_L g1503 ( .A(n_1478), .B(n_1374), .Y(n_1503) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1432), .Y(n_1504) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_1412), .B(n_1375), .Y(n_1505) );
NAND2xp5_ASAP7_75t_L g1506 ( .A(n_1445), .B(n_1331), .Y(n_1506) );
OR2x2_ASAP7_75t_L g1507 ( .A(n_1431), .B(n_1376), .Y(n_1507) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1431), .Y(n_1508) );
NAND2xp5_ASAP7_75t_L g1509 ( .A(n_1417), .B(n_1377), .Y(n_1509) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1434), .Y(n_1510) );
INVx2_ASAP7_75t_L g1511 ( .A(n_1413), .Y(n_1511) );
INVx4_ASAP7_75t_L g1512 ( .A(n_1416), .Y(n_1512) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1447), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1426), .B(n_1377), .Y(n_1514) );
OR2x2_ASAP7_75t_L g1515 ( .A(n_1458), .B(n_1376), .Y(n_1515) );
NAND2xp5_ASAP7_75t_L g1516 ( .A(n_1418), .B(n_1381), .Y(n_1516) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1448), .Y(n_1517) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1454), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1519 ( .A(n_1426), .B(n_1381), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_1456), .B(n_1383), .Y(n_1520) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1466), .Y(n_1521) );
INVxp67_ASAP7_75t_L g1522 ( .A(n_1462), .Y(n_1522) );
AND2x2_ASAP7_75t_L g1523 ( .A(n_1456), .B(n_1383), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1460), .B(n_1397), .Y(n_1524) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1414), .Y(n_1525) );
NAND2xp5_ASAP7_75t_L g1526 ( .A(n_1427), .B(n_1380), .Y(n_1526) );
INVxp67_ASAP7_75t_L g1527 ( .A(n_1472), .Y(n_1527) );
OR2x2_ASAP7_75t_L g1528 ( .A(n_1458), .B(n_1380), .Y(n_1528) );
AOI222xp33_ASAP7_75t_L g1529 ( .A1(n_1438), .A2(n_1401), .B1(n_1379), .B2(n_1360), .C1(n_1366), .C2(n_1343), .Y(n_1529) );
NAND2xp5_ASAP7_75t_L g1530 ( .A(n_1410), .B(n_1388), .Y(n_1530) );
AND2x2_ASAP7_75t_SL g1531 ( .A(n_1428), .B(n_1343), .Y(n_1531) );
INVxp67_ASAP7_75t_SL g1532 ( .A(n_1485), .Y(n_1532) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_1460), .B(n_1397), .Y(n_1533) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1484), .Y(n_1534) );
NOR2xp33_ASAP7_75t_L g1535 ( .A(n_1423), .B(n_1309), .Y(n_1535) );
OR2x2_ASAP7_75t_L g1536 ( .A(n_1440), .B(n_1388), .Y(n_1536) );
NAND2xp5_ASAP7_75t_L g1537 ( .A(n_1419), .B(n_1390), .Y(n_1537) );
NAND2xp5_ASAP7_75t_L g1538 ( .A(n_1422), .B(n_1390), .Y(n_1538) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1461), .B(n_1402), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1540 ( .A(n_1461), .B(n_1402), .Y(n_1540) );
INVx2_ASAP7_75t_L g1541 ( .A(n_1425), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_1429), .B(n_1350), .Y(n_1542) );
OR2x2_ASAP7_75t_L g1543 ( .A(n_1440), .B(n_1391), .Y(n_1543) );
INVx1_ASAP7_75t_SL g1544 ( .A(n_1416), .Y(n_1544) );
NAND2xp5_ASAP7_75t_L g1545 ( .A(n_1437), .B(n_1409), .Y(n_1545) );
OR2x2_ASAP7_75t_L g1546 ( .A(n_1455), .B(n_1391), .Y(n_1546) );
AND2x2_ASAP7_75t_L g1547 ( .A(n_1429), .B(n_1350), .Y(n_1547) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1492), .Y(n_1548) );
OR2x2_ASAP7_75t_L g1549 ( .A(n_1490), .B(n_1463), .Y(n_1549) );
OR2x2_ASAP7_75t_L g1550 ( .A(n_1490), .B(n_1463), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1551 ( .A(n_1493), .B(n_1467), .Y(n_1551) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1507), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1553 ( .A(n_1493), .B(n_1467), .Y(n_1553) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1507), .Y(n_1554) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1495), .Y(n_1555) );
NAND2xp5_ASAP7_75t_SL g1556 ( .A(n_1512), .B(n_1489), .Y(n_1556) );
NAND2xp5_ASAP7_75t_L g1557 ( .A(n_1496), .B(n_1433), .Y(n_1557) );
AND2x2_ASAP7_75t_L g1558 ( .A(n_1524), .B(n_1475), .Y(n_1558) );
OR2x2_ASAP7_75t_L g1559 ( .A(n_1542), .B(n_1455), .Y(n_1559) );
OAI21xp33_ASAP7_75t_SL g1560 ( .A1(n_1512), .A2(n_1444), .B(n_1435), .Y(n_1560) );
BUFx2_ASAP7_75t_L g1561 ( .A(n_1512), .Y(n_1561) );
HB1xp67_ASAP7_75t_L g1562 ( .A(n_1542), .Y(n_1562) );
OR2x2_ASAP7_75t_L g1563 ( .A(n_1547), .B(n_1475), .Y(n_1563) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1495), .Y(n_1564) );
AO21x1_ASAP7_75t_L g1565 ( .A1(n_1532), .A2(n_1459), .B(n_1428), .Y(n_1565) );
NOR2xp33_ASAP7_75t_L g1566 ( .A(n_1544), .B(n_1421), .Y(n_1566) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_1496), .B(n_1433), .Y(n_1567) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1547), .Y(n_1568) );
AND2x2_ASAP7_75t_L g1569 ( .A(n_1524), .B(n_1533), .Y(n_1569) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_1505), .B(n_1508), .Y(n_1570) );
AOI222xp33_ASAP7_75t_L g1571 ( .A1(n_1502), .A2(n_1473), .B1(n_1415), .B2(n_1439), .C1(n_1446), .C2(n_1477), .Y(n_1571) );
NAND2xp5_ASAP7_75t_L g1572 ( .A(n_1505), .B(n_1436), .Y(n_1572) );
INVx2_ASAP7_75t_L g1573 ( .A(n_1511), .Y(n_1573) );
NOR2xp33_ASAP7_75t_L g1574 ( .A(n_1527), .B(n_1309), .Y(n_1574) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1504), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1576 ( .A(n_1533), .B(n_1436), .Y(n_1576) );
AOI21xp33_ASAP7_75t_L g1577 ( .A1(n_1535), .A2(n_1476), .B(n_1334), .Y(n_1577) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1520), .B(n_1469), .Y(n_1578) );
NAND2xp5_ASAP7_75t_L g1579 ( .A(n_1520), .B(n_1469), .Y(n_1579) );
NAND2xp5_ASAP7_75t_L g1580 ( .A(n_1523), .B(n_1470), .Y(n_1580) );
NAND2xp5_ASAP7_75t_L g1581 ( .A(n_1523), .B(n_1470), .Y(n_1581) );
INVx2_ASAP7_75t_SL g1582 ( .A(n_1494), .Y(n_1582) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1504), .Y(n_1583) );
NAND2xp5_ASAP7_75t_L g1584 ( .A(n_1514), .B(n_1465), .Y(n_1584) );
INVxp67_ASAP7_75t_L g1585 ( .A(n_1500), .Y(n_1585) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1513), .Y(n_1586) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1513), .Y(n_1587) );
AOI21xp5_ASAP7_75t_L g1588 ( .A1(n_1556), .A2(n_1531), .B(n_1494), .Y(n_1588) );
AOI22xp5_ASAP7_75t_L g1589 ( .A1(n_1566), .A2(n_1529), .B1(n_1506), .B2(n_1473), .Y(n_1589) );
OAI22xp33_ASAP7_75t_L g1590 ( .A1(n_1561), .A2(n_1394), .B1(n_1351), .B2(n_1400), .Y(n_1590) );
AOI222xp33_ASAP7_75t_L g1591 ( .A1(n_1556), .A2(n_1498), .B1(n_1525), .B2(n_1522), .C1(n_1509), .C2(n_1516), .Y(n_1591) );
NAND2x1_ASAP7_75t_L g1592 ( .A(n_1561), .B(n_1468), .Y(n_1592) );
NAND2xp5_ASAP7_75t_L g1593 ( .A(n_1571), .B(n_1539), .Y(n_1593) );
OA21x2_ASAP7_75t_L g1594 ( .A1(n_1565), .A2(n_1499), .B(n_1526), .Y(n_1594) );
AOI322xp5_ASAP7_75t_L g1595 ( .A1(n_1574), .A2(n_1514), .A3(n_1519), .B1(n_1531), .B2(n_1539), .C1(n_1540), .C2(n_1545), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_1569), .B(n_1519), .Y(n_1596) );
INVxp67_ASAP7_75t_L g1597 ( .A(n_1548), .Y(n_1597) );
AOI22xp33_ASAP7_75t_L g1598 ( .A1(n_1585), .A2(n_1360), .B1(n_1366), .B2(n_1491), .Y(n_1598) );
OAI211xp5_ASAP7_75t_L g1599 ( .A1(n_1560), .A2(n_1394), .B(n_1457), .C(n_1405), .Y(n_1599) );
INVx1_ASAP7_75t_SL g1600 ( .A(n_1582), .Y(n_1600) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1562), .Y(n_1601) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1555), .Y(n_1602) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1564), .Y(n_1603) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1575), .Y(n_1604) );
NAND2xp5_ASAP7_75t_L g1605 ( .A(n_1568), .B(n_1540), .Y(n_1605) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1583), .Y(n_1606) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1586), .Y(n_1607) );
OAI22xp33_ASAP7_75t_L g1608 ( .A1(n_1582), .A2(n_1394), .B1(n_1351), .B2(n_1396), .Y(n_1608) );
A2O1A1Ixp33_ASAP7_75t_L g1609 ( .A1(n_1577), .A2(n_1501), .B(n_1483), .C(n_1366), .Y(n_1609) );
NOR3xp33_ASAP7_75t_L g1610 ( .A(n_1587), .B(n_1258), .C(n_1530), .Y(n_1610) );
AOI221x1_ASAP7_75t_L g1611 ( .A1(n_1552), .A2(n_1360), .B1(n_1491), .B2(n_1441), .C(n_1517), .Y(n_1611) );
AOI221xp5_ASAP7_75t_L g1612 ( .A1(n_1554), .A2(n_1538), .B1(n_1537), .B2(n_1534), .C(n_1510), .Y(n_1612) );
OAI211xp5_ASAP7_75t_L g1613 ( .A1(n_1565), .A2(n_1394), .B(n_1482), .C(n_1488), .Y(n_1613) );
OAI22xp5_ASAP7_75t_L g1614 ( .A1(n_1563), .A2(n_1394), .B1(n_1491), .B2(n_1497), .Y(n_1614) );
INVxp67_ASAP7_75t_SL g1615 ( .A(n_1573), .Y(n_1615) );
AOI21xp5_ASAP7_75t_SL g1616 ( .A1(n_1594), .A2(n_1309), .B(n_1399), .Y(n_1616) );
AOI21xp33_ASAP7_75t_SL g1617 ( .A1(n_1594), .A2(n_1563), .B(n_1569), .Y(n_1617) );
NAND2xp5_ASAP7_75t_L g1618 ( .A(n_1593), .B(n_1568), .Y(n_1618) );
OAI32xp33_ASAP7_75t_L g1619 ( .A1(n_1600), .A2(n_1559), .A3(n_1550), .B1(n_1549), .B2(n_1584), .Y(n_1619) );
INVxp67_ASAP7_75t_L g1620 ( .A(n_1591), .Y(n_1620) );
AOI32xp33_ASAP7_75t_L g1621 ( .A1(n_1610), .A2(n_1551), .A3(n_1553), .B1(n_1576), .B2(n_1558), .Y(n_1621) );
OAI211xp5_ASAP7_75t_L g1622 ( .A1(n_1588), .A2(n_1486), .B(n_1549), .C(n_1550), .Y(n_1622) );
OAI21xp5_ASAP7_75t_SL g1623 ( .A1(n_1599), .A2(n_1483), .B(n_1441), .Y(n_1623) );
O2A1O1Ixp33_ASAP7_75t_L g1624 ( .A1(n_1613), .A2(n_1559), .B(n_1570), .C(n_1399), .Y(n_1624) );
AOI22xp33_ASAP7_75t_L g1625 ( .A1(n_1589), .A2(n_1441), .B1(n_1480), .B2(n_1389), .Y(n_1625) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1602), .Y(n_1626) );
AOI32xp33_ASAP7_75t_L g1627 ( .A1(n_1610), .A2(n_1551), .A3(n_1553), .B1(n_1576), .B2(n_1558), .Y(n_1627) );
OAI22xp5_ASAP7_75t_L g1628 ( .A1(n_1609), .A2(n_1581), .B1(n_1580), .B2(n_1579), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1629 ( .A(n_1596), .B(n_1557), .Y(n_1629) );
NAND2xp5_ASAP7_75t_L g1630 ( .A(n_1612), .B(n_1578), .Y(n_1630) );
INVxp67_ASAP7_75t_L g1631 ( .A(n_1603), .Y(n_1631) );
AOI221xp5_ASAP7_75t_L g1632 ( .A1(n_1597), .A2(n_1572), .B1(n_1567), .B2(n_1518), .C(n_1521), .Y(n_1632) );
NAND3xp33_ASAP7_75t_L g1633 ( .A(n_1595), .B(n_1528), .C(n_1515), .Y(n_1633) );
NAND2xp5_ASAP7_75t_L g1634 ( .A(n_1597), .B(n_1515), .Y(n_1634) );
OAI21xp5_ASAP7_75t_L g1635 ( .A1(n_1611), .A2(n_1503), .B(n_1497), .Y(n_1635) );
OAI221xp5_ASAP7_75t_SL g1636 ( .A1(n_1620), .A2(n_1621), .B1(n_1627), .B2(n_1622), .C(n_1625), .Y(n_1636) );
NAND4xp25_ASAP7_75t_SL g1637 ( .A(n_1624), .B(n_1598), .C(n_1605), .D(n_1601), .Y(n_1637) );
AOI211xp5_ASAP7_75t_L g1638 ( .A1(n_1617), .A2(n_1590), .B(n_1608), .C(n_1614), .Y(n_1638) );
AOI221x1_ASAP7_75t_L g1639 ( .A1(n_1616), .A2(n_1604), .B1(n_1606), .B2(n_1607), .C(n_1221), .Y(n_1639) );
INVx2_ASAP7_75t_L g1640 ( .A(n_1626), .Y(n_1640) );
O2A1O1Ixp5_ASAP7_75t_L g1641 ( .A1(n_1619), .A2(n_1618), .B(n_1628), .C(n_1630), .Y(n_1641) );
NAND4xp25_ASAP7_75t_L g1642 ( .A(n_1624), .B(n_1282), .C(n_1451), .D(n_1450), .Y(n_1642) );
OR2x2_ASAP7_75t_L g1643 ( .A(n_1633), .B(n_1615), .Y(n_1643) );
INVx2_ASAP7_75t_L g1644 ( .A(n_1631), .Y(n_1644) );
AOI211xp5_ASAP7_75t_SL g1645 ( .A1(n_1623), .A2(n_1259), .B(n_1221), .C(n_1313), .Y(n_1645) );
NOR2x1_ASAP7_75t_L g1646 ( .A(n_1635), .B(n_1592), .Y(n_1646) );
NOR3xp33_ASAP7_75t_L g1647 ( .A(n_1632), .B(n_1615), .C(n_1268), .Y(n_1647) );
OAI22xp5_ASAP7_75t_R g1648 ( .A1(n_1629), .A2(n_1521), .B1(n_1487), .B2(n_1389), .Y(n_1648) );
NAND2xp33_ASAP7_75t_R g1649 ( .A(n_1634), .B(n_1221), .Y(n_1649) );
OAI211xp5_ASAP7_75t_L g1650 ( .A1(n_1636), .A2(n_1398), .B(n_1503), .C(n_1259), .Y(n_1650) );
NOR2xp33_ASAP7_75t_L g1651 ( .A(n_1637), .B(n_1528), .Y(n_1651) );
AOI211x1_ASAP7_75t_L g1652 ( .A1(n_1642), .A2(n_1452), .B(n_1449), .C(n_1453), .Y(n_1652) );
NAND3xp33_ASAP7_75t_L g1653 ( .A(n_1641), .B(n_1573), .C(n_1546), .Y(n_1653) );
OAI321xp33_ASAP7_75t_L g1654 ( .A1(n_1642), .A2(n_1546), .A3(n_1543), .B1(n_1536), .B2(n_1398), .C(n_1443), .Y(n_1654) );
NOR2xp33_ASAP7_75t_L g1655 ( .A(n_1644), .B(n_1543), .Y(n_1655) );
NAND4xp75_ASAP7_75t_L g1656 ( .A(n_1646), .B(n_1272), .C(n_1270), .D(n_1246), .Y(n_1656) );
NOR4xp25_ASAP7_75t_L g1657 ( .A(n_1643), .B(n_1322), .C(n_1313), .D(n_1259), .Y(n_1657) );
NAND2xp5_ASAP7_75t_L g1658 ( .A(n_1640), .B(n_1536), .Y(n_1658) );
OAI221xp5_ASAP7_75t_SL g1659 ( .A1(n_1638), .A2(n_1442), .B1(n_1481), .B2(n_1479), .C(n_1449), .Y(n_1659) );
O2A1O1Ixp33_ASAP7_75t_L g1660 ( .A1(n_1650), .A2(n_1659), .B(n_1654), .C(n_1651), .Y(n_1660) );
NOR2x1_ASAP7_75t_L g1661 ( .A(n_1653), .B(n_1648), .Y(n_1661) );
NAND2xp5_ASAP7_75t_SL g1662 ( .A(n_1657), .B(n_1647), .Y(n_1662) );
NOR4xp75_ASAP7_75t_L g1663 ( .A(n_1656), .B(n_1645), .C(n_1649), .D(n_1639), .Y(n_1663) );
NAND4xp75_ASAP7_75t_L g1664 ( .A(n_1652), .B(n_1645), .C(n_1272), .D(n_1270), .Y(n_1664) );
NOR3xp33_ASAP7_75t_L g1665 ( .A(n_1655), .B(n_1313), .C(n_1322), .Y(n_1665) );
OAI21xp5_ASAP7_75t_L g1666 ( .A1(n_1658), .A2(n_1282), .B(n_1480), .Y(n_1666) );
INVx2_ASAP7_75t_L g1667 ( .A(n_1664), .Y(n_1667) );
INVx1_ASAP7_75t_L g1668 ( .A(n_1662), .Y(n_1668) );
NAND3xp33_ASAP7_75t_SL g1669 ( .A(n_1663), .B(n_1286), .C(n_1263), .Y(n_1669) );
INVx3_ASAP7_75t_L g1670 ( .A(n_1661), .Y(n_1670) );
INVx2_ASAP7_75t_L g1671 ( .A(n_1666), .Y(n_1671) );
INVx2_ASAP7_75t_L g1672 ( .A(n_1665), .Y(n_1672) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1668), .Y(n_1673) );
AOI22xp5_ASAP7_75t_L g1674 ( .A1(n_1670), .A2(n_1660), .B1(n_1282), .B2(n_1268), .Y(n_1674) );
AND2x2_ASAP7_75t_SL g1675 ( .A(n_1670), .B(n_1268), .Y(n_1675) );
AO22x2_ASAP7_75t_L g1676 ( .A1(n_1668), .A2(n_1290), .B1(n_1283), .B2(n_1541), .Y(n_1676) );
XOR2xp5_ASAP7_75t_L g1677 ( .A(n_1667), .B(n_1290), .Y(n_1677) );
AOI22xp5_ASAP7_75t_L g1678 ( .A1(n_1677), .A2(n_1672), .B1(n_1669), .B2(n_1671), .Y(n_1678) );
NOR2x1_ASAP7_75t_L g1679 ( .A(n_1673), .B(n_1299), .Y(n_1679) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1674), .Y(n_1680) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1676), .Y(n_1681) );
BUFx2_ASAP7_75t_L g1682 ( .A(n_1681), .Y(n_1682) );
OAI22x1_ASAP7_75t_L g1683 ( .A1(n_1678), .A2(n_1675), .B1(n_1283), .B2(n_1272), .Y(n_1683) );
BUFx8_ASAP7_75t_L g1684 ( .A(n_1680), .Y(n_1684) );
AOI22xp5_ASAP7_75t_L g1685 ( .A1(n_1679), .A2(n_1299), .B1(n_1283), .B2(n_1251), .Y(n_1685) );
AOI222xp33_ASAP7_75t_L g1686 ( .A1(n_1684), .A2(n_1682), .B1(n_1683), .B2(n_1685), .C1(n_1384), .C2(n_1354), .Y(n_1686) );
OAI21xp5_ASAP7_75t_L g1687 ( .A1(n_1686), .A2(n_1301), .B(n_1263), .Y(n_1687) );
AOI21xp5_ASAP7_75t_L g1688 ( .A1(n_1687), .A2(n_1254), .B(n_1288), .Y(n_1688) );
endmodule