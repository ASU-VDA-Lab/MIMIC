module fake_netlist_5_2208_n_767 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_767);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_767;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_443;
wire n_372;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_516;
wire n_385;
wire n_498;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_344;
wire n_287;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_432;
wire n_164;
wire n_553;
wire n_395;
wire n_727;
wire n_311;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_144;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_113),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_43),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_24),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_78),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_57),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_108),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_77),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_58),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_15),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_83),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_59),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_5),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_36),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_42),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_15),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_93),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_54),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_129),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_29),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_76),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_26),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_92),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_142),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_44),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_50),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_70),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_41),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_80),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_102),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

BUFx8_ASAP7_75t_SL g183 ( 
.A(n_27),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_17),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_62),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_109),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_141),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_3),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_137),
.Y(n_191)
);

BUFx8_ASAP7_75t_SL g192 ( 
.A(n_63),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_72),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_128),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_35),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_14),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_145),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

AND2x4_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_174),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_155),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_0),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_147),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_157),
.B(n_0),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_1),
.Y(n_214)
);

BUFx8_ASAP7_75t_SL g215 ( 
.A(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_171),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_1),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_146),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_148),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_153),
.B(n_143),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_159),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_164),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_162),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

BUFx8_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_186),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

CKINVDCx6p67_ASAP7_75t_R g235 ( 
.A(n_144),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_149),
.B(n_2),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

AO22x2_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_224),
.B1(n_217),
.B2(n_214),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_150),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_224),
.A2(n_144),
.B1(n_163),
.B2(n_191),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_233),
.A2(n_196),
.B1(n_151),
.B2(n_152),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_163),
.B1(n_191),
.B2(n_189),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_219),
.B(n_192),
.Y(n_245)
);

AO22x2_ASAP7_75t_L g246 ( 
.A1(n_206),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_233),
.A2(n_188),
.B1(n_187),
.B2(n_181),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_L g248 ( 
.A1(n_213),
.A2(n_179),
.B1(n_177),
.B2(n_173),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_165),
.B1(n_170),
.B2(n_169),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_200),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_219),
.A2(n_206),
.B1(n_213),
.B2(n_202),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_215),
.Y(n_252)
);

AO22x2_ASAP7_75t_L g253 ( 
.A1(n_206),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_212),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_206),
.B(n_154),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_202),
.B(n_156),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_160),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_209),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_L g259 ( 
.A1(n_209),
.A2(n_172),
.B1(n_166),
.B2(n_161),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_219),
.B(n_22),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_23),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_219),
.B(n_211),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_201),
.Y(n_263)
);

AO22x2_ASAP7_75t_L g264 ( 
.A1(n_211),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_200),
.Y(n_266)
);

AND2x2_ASAP7_75t_SL g267 ( 
.A(n_230),
.B(n_10),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_209),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g270 ( 
.A1(n_234),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_25),
.Y(n_271)
);

AO22x2_ASAP7_75t_L g272 ( 
.A1(n_221),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_272)
);

AND2x6_ASAP7_75t_L g273 ( 
.A(n_221),
.B(n_28),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_210),
.Y(n_274)
);

AND2x2_ASAP7_75t_SL g275 ( 
.A(n_221),
.B(n_19),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_234),
.A2(n_20),
.B1(n_21),
.B2(n_30),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_221),
.B(n_20),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_201),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_21),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_235),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_218),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_210),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_201),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_218),
.A2(n_39),
.B1(n_40),
.B2(n_45),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_239),
.B(n_222),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_240),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_228),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_222),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_199),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_249),
.B(n_228),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_257),
.B(n_199),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_258),
.Y(n_295)
);

AOI21x1_ASAP7_75t_L g296 ( 
.A1(n_250),
.A2(n_220),
.B(n_231),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_226),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_275),
.B(n_223),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_263),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_263),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_250),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

OR2x6_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_207),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_242),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_256),
.B(n_226),
.Y(n_307)
);

NOR2xp67_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_199),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_242),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_241),
.Y(n_310)
);

AND2x2_ASAP7_75t_SL g311 ( 
.A(n_267),
.B(n_281),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_273),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_273),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_271),
.B(n_198),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_205),
.Y(n_316)
);

XOR2x2_ASAP7_75t_L g317 ( 
.A(n_279),
.B(n_207),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

INVx3_ASAP7_75t_R g319 ( 
.A(n_254),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_272),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_272),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_246),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_246),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_244),
.B(n_228),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_253),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_261),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_253),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_259),
.B(n_228),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_247),
.B(n_220),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_248),
.B(n_220),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_281),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_243),
.B(n_231),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_265),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_276),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_260),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_245),
.B(n_198),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_238),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_252),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_284),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_268),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_238),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_269),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_270),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_274),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_274),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_274),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_255),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_307),
.B(n_231),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_307),
.B(n_205),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_302),
.Y(n_351)
);

AND2x4_ASAP7_75t_L g352 ( 
.A(n_318),
.B(n_46),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_310),
.B(n_348),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_318),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_290),
.B(n_204),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_348),
.B(n_223),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_336),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_326),
.B(n_227),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_312),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_290),
.B(n_204),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_285),
.B(n_227),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_296),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_302),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_326),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_227),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_296),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_313),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_286),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_316),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_285),
.B(n_227),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_311),
.A2(n_229),
.B1(n_232),
.B2(n_225),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_335),
.B(n_229),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_286),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_331),
.B(n_223),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_330),
.A2(n_229),
.B(n_203),
.Y(n_375)
);

AND2x2_ASAP7_75t_SL g376 ( 
.A(n_311),
.B(n_223),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_299),
.B(n_315),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_316),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_299),
.B(n_229),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_288),
.B(n_223),
.Y(n_380)
);

AND2x4_ASAP7_75t_L g381 ( 
.A(n_314),
.B(n_47),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_336),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_292),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_315),
.B(n_298),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_292),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_298),
.B(n_223),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_289),
.B(n_225),
.Y(n_387)
);

AND2x6_ASAP7_75t_L g388 ( 
.A(n_320),
.B(n_201),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_332),
.B(n_225),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_347),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_297),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_345),
.B(n_225),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_346),
.B(n_225),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_303),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_304),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_329),
.B(n_225),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_340),
.B(n_232),
.Y(n_397)
);

AND2x2_ASAP7_75t_SL g398 ( 
.A(n_324),
.B(n_232),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_305),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_305),
.B(n_232),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_300),
.B(n_232),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_301),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_338),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_305),
.B(n_232),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_333),
.B(n_201),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_305),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_338),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_291),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_294),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_321),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_322),
.Y(n_413)
);

AND2x2_ASAP7_75t_SL g414 ( 
.A(n_328),
.B(n_201),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_323),
.Y(n_415)
);

NOR2xp67_ASAP7_75t_L g416 ( 
.A(n_357),
.B(n_295),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_351),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g418 ( 
.A(n_397),
.B(n_295),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_354),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_369),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_368),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_382),
.B(n_306),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_368),
.Y(n_424)
);

BUFx12f_ASAP7_75t_L g425 ( 
.A(n_399),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_384),
.B(n_306),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_344),
.Y(n_427)
);

OR2x6_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_341),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_409),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_396),
.B(n_344),
.Y(n_430)
);

BUFx12f_ASAP7_75t_L g431 ( 
.A(n_412),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_384),
.B(n_343),
.Y(n_432)
);

NOR2x1_ASAP7_75t_L g433 ( 
.A(n_382),
.B(n_308),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_382),
.B(n_334),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_368),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_364),
.B(n_325),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_409),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_376),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_363),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_369),
.B(n_337),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_350),
.Y(n_441)
);

NAND2x1p5_ASAP7_75t_L g442 ( 
.A(n_352),
.B(n_381),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_414),
.B(n_293),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_391),
.B(n_327),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_391),
.B(n_287),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_389),
.B(n_309),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_414),
.B(n_309),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_406),
.Y(n_448)
);

AND2x6_ASAP7_75t_L g449 ( 
.A(n_371),
.B(n_319),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_391),
.B(n_339),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_409),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_350),
.B(n_317),
.Y(n_452)
);

BUFx4f_ASAP7_75t_L g453 ( 
.A(n_409),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_376),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_373),
.Y(n_455)
);

BUFx8_ASAP7_75t_L g456 ( 
.A(n_415),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_409),
.Y(n_457)
);

OR2x6_ASAP7_75t_L g458 ( 
.A(n_400),
.B(n_319),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_414),
.B(n_339),
.Y(n_459)
);

INVx6_ASAP7_75t_L g460 ( 
.A(n_409),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_412),
.B(n_48),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_413),
.B(n_49),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_361),
.B(n_199),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_355),
.B(n_317),
.Y(n_464)
);

CKINVDCx6p67_ASAP7_75t_R g465 ( 
.A(n_378),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_398),
.B(n_199),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_415),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_400),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_349),
.B(n_199),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_373),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_389),
.B(n_377),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_417),
.Y(n_472)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

NAND2x1p5_ASAP7_75t_L g474 ( 
.A(n_453),
.B(n_352),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_422),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_425),
.Y(n_476)
);

OR2x6_ASAP7_75t_L g477 ( 
.A(n_442),
.B(n_352),
.Y(n_477)
);

BUFx2_ASAP7_75t_SL g478 ( 
.A(n_429),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_440),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g480 ( 
.A(n_453),
.Y(n_480)
);

CKINVDCx11_ASAP7_75t_R g481 ( 
.A(n_465),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_420),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_421),
.Y(n_483)
);

BUFx2_ASAP7_75t_SL g484 ( 
.A(n_429),
.Y(n_484)
);

BUFx2_ASAP7_75t_SL g485 ( 
.A(n_437),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_431),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_426),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_448),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_424),
.Y(n_489)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_437),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_450),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_460),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_437),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_442),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_468),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_428),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_460),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_451),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_450),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_456),
.Y(n_500)
);

BUFx12f_ASAP7_75t_L g501 ( 
.A(n_456),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_451),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_444),
.Y(n_503)
);

INVx5_ASAP7_75t_SL g504 ( 
.A(n_458),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_443),
.A2(n_376),
.B1(n_398),
.B2(n_361),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_464),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_439),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_451),
.Y(n_508)
);

NAND2x1p5_ASAP7_75t_L g509 ( 
.A(n_457),
.B(n_352),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_457),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_435),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_428),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_444),
.Y(n_513)
);

NAND2x1p5_ASAP7_75t_L g514 ( 
.A(n_457),
.B(n_381),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_455),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_428),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_427),
.B(n_370),
.Y(n_517)
);

CKINVDCx6p67_ASAP7_75t_R g518 ( 
.A(n_458),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_419),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_472),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_493),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_483),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_488),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_472),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_473),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_487),
.A2(n_447),
.B1(n_443),
.B2(n_459),
.Y(n_526)
);

NAND2x1p5_ASAP7_75t_L g527 ( 
.A(n_490),
.B(n_419),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_505),
.A2(n_447),
.B1(n_459),
.B2(n_446),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_506),
.A2(n_446),
.B1(n_423),
.B2(n_432),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_496),
.A2(n_452),
.B(n_441),
.Y(n_530)
);

CKINVDCx11_ASAP7_75t_R g531 ( 
.A(n_481),
.Y(n_531)
);

BUFx8_ASAP7_75t_L g532 ( 
.A(n_501),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_493),
.Y(n_533)
);

NAND2x1p5_ASAP7_75t_L g534 ( 
.A(n_490),
.B(n_467),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_475),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_493),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_496),
.A2(n_512),
.B1(n_516),
.B2(n_449),
.Y(n_537)
);

CKINVDCx11_ASAP7_75t_R g538 ( 
.A(n_501),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_475),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_517),
.B(n_427),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_474),
.A2(n_398),
.B1(n_430),
.B2(n_438),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_479),
.B(n_378),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_490),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_483),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_473),
.Y(n_545)
);

OAI21xp33_ASAP7_75t_SL g546 ( 
.A1(n_477),
.A2(n_371),
.B(n_375),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_474),
.A2(n_438),
.B1(n_454),
.B2(n_430),
.Y(n_547)
);

BUFx12f_ASAP7_75t_L g548 ( 
.A(n_500),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_488),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_474),
.A2(n_454),
.B1(n_436),
.B2(n_433),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_512),
.A2(n_445),
.B1(n_449),
.B2(n_434),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_507),
.B(n_370),
.Y(n_552)
);

BUFx12f_ASAP7_75t_L g553 ( 
.A(n_500),
.Y(n_553)
);

BUFx2_ASAP7_75t_SL g554 ( 
.A(n_486),
.Y(n_554)
);

BUFx4f_ASAP7_75t_L g555 ( 
.A(n_518),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_507),
.A2(n_436),
.B1(n_462),
.B2(n_471),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_495),
.Y(n_557)
);

BUFx12f_ASAP7_75t_L g558 ( 
.A(n_486),
.Y(n_558)
);

BUFx12f_ASAP7_75t_L g559 ( 
.A(n_476),
.Y(n_559)
);

NAND2x1p5_ASAP7_75t_L g560 ( 
.A(n_490),
.B(n_462),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_528),
.A2(n_526),
.B1(n_529),
.B2(n_540),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_529),
.B(n_495),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_531),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_552),
.B(n_482),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_520),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_525),
.Y(n_566)
);

AOI21xp33_ASAP7_75t_SL g567 ( 
.A1(n_542),
.A2(n_458),
.B(n_353),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_522),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_521),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_528),
.A2(n_416),
.B1(n_418),
.B2(n_477),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_556),
.A2(n_445),
.B1(n_491),
.B2(n_499),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_551),
.A2(n_477),
.B1(n_516),
.B2(n_509),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_556),
.A2(n_499),
.B1(n_491),
.B2(n_449),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_544),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_546),
.A2(n_449),
.B1(n_390),
.B2(n_471),
.Y(n_575)
);

INVx5_ASAP7_75t_SL g576 ( 
.A(n_521),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_521),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_557),
.B(n_503),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_524),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_557),
.B(n_349),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_546),
.A2(n_390),
.B1(n_374),
.B2(n_539),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_535),
.A2(n_355),
.B1(n_360),
.B2(n_466),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_525),
.Y(n_583)
);

OAI222xp33_ASAP7_75t_L g584 ( 
.A1(n_537),
.A2(n_477),
.B1(n_494),
.B2(n_405),
.C1(n_515),
.C2(n_509),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_541),
.A2(n_360),
.B1(n_466),
.B2(n_375),
.Y(n_585)
);

AOI222xp33_ASAP7_75t_L g586 ( 
.A1(n_530),
.A2(n_513),
.B1(n_503),
.B2(n_504),
.C1(n_413),
.C2(n_404),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_533),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_533),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_533),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_550),
.A2(n_461),
.B1(n_513),
.B2(n_477),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_530),
.B(n_537),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_560),
.A2(n_509),
.B1(n_555),
.B2(n_518),
.Y(n_592)
);

AOI222xp33_ASAP7_75t_L g593 ( 
.A1(n_532),
.A2(n_504),
.B1(n_413),
.B2(n_404),
.C1(n_407),
.C2(n_403),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_538),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_541),
.A2(n_363),
.B1(n_405),
.B2(n_515),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_555),
.A2(n_514),
.B1(n_504),
.B2(n_547),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_536),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_548),
.A2(n_410),
.B1(n_489),
.B2(n_511),
.Y(n_598)
);

BUFx12f_ASAP7_75t_L g599 ( 
.A(n_532),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_553),
.A2(n_410),
.B1(n_489),
.B2(n_511),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_534),
.A2(n_381),
.B(n_480),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_523),
.B(n_411),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_SL g603 ( 
.A1(n_545),
.A2(n_381),
.B(n_480),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_549),
.B(n_504),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_554),
.A2(n_410),
.B1(n_395),
.B2(n_408),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_545),
.A2(n_407),
.B(n_403),
.Y(n_606)
);

OAI22xp33_ASAP7_75t_L g607 ( 
.A1(n_558),
.A2(n_514),
.B1(n_559),
.B2(n_379),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_543),
.B(n_476),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_586),
.A2(n_395),
.B1(n_408),
.B2(n_386),
.Y(n_609)
);

OAI21xp5_ASAP7_75t_SL g610 ( 
.A1(n_561),
.A2(n_356),
.B(n_514),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_561),
.A2(n_408),
.B1(n_402),
.B2(n_358),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_591),
.A2(n_386),
.B1(n_402),
.B2(n_469),
.Y(n_612)
);

OAI22xp33_ASAP7_75t_L g613 ( 
.A1(n_564),
.A2(n_519),
.B1(n_543),
.B2(n_527),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_570),
.A2(n_394),
.B1(n_393),
.B2(n_392),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_571),
.A2(n_497),
.B1(n_492),
.B2(n_519),
.Y(n_615)
);

AOI221xp5_ASAP7_75t_L g616 ( 
.A1(n_567),
.A2(n_581),
.B1(n_575),
.B2(n_562),
.C(n_580),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_573),
.A2(n_394),
.B1(n_393),
.B2(n_392),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_585),
.A2(n_497),
.B1(n_492),
.B2(n_519),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_578),
.B(n_411),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_604),
.Y(n_620)
);

OA21x2_ASAP7_75t_L g621 ( 
.A1(n_581),
.A2(n_358),
.B(n_372),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_568),
.B(n_536),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_574),
.B(n_411),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_585),
.A2(n_590),
.B1(n_605),
.B2(n_598),
.Y(n_624)
);

AOI222xp33_ASAP7_75t_L g625 ( 
.A1(n_582),
.A2(n_380),
.B1(n_372),
.B2(n_365),
.C1(n_394),
.C2(n_385),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_565),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_579),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_593),
.A2(n_359),
.B1(n_380),
.B2(n_365),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_605),
.A2(n_359),
.B1(n_508),
.B2(n_484),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_572),
.A2(n_359),
.B1(n_388),
.B2(n_463),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_596),
.A2(n_359),
.B1(n_388),
.B2(n_385),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_598),
.A2(n_359),
.B1(n_508),
.B2(n_485),
.Y(n_632)
);

OAI221xp5_ASAP7_75t_L g633 ( 
.A1(n_603),
.A2(n_387),
.B1(n_373),
.B2(n_383),
.C(n_385),
.Y(n_633)
);

AOI222xp33_ASAP7_75t_L g634 ( 
.A1(n_582),
.A2(n_383),
.B1(n_470),
.B2(n_388),
.C1(n_359),
.C2(n_367),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_575),
.A2(n_388),
.B1(n_383),
.B2(n_367),
.Y(n_635)
);

NAND4xp25_ASAP7_75t_L g636 ( 
.A(n_595),
.B(n_498),
.C(n_473),
.D(n_401),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_607),
.A2(n_600),
.B1(n_595),
.B2(n_599),
.Y(n_637)
);

NAND3xp33_ASAP7_75t_SL g638 ( 
.A(n_594),
.B(n_498),
.C(n_485),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_600),
.B(n_493),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_607),
.A2(n_388),
.B1(n_367),
.B2(n_354),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_592),
.A2(n_388),
.B1(n_367),
.B2(n_354),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_608),
.A2(n_388),
.B1(n_498),
.B2(n_510),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_608),
.A2(n_597),
.B1(n_602),
.B2(n_587),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_601),
.A2(n_478),
.B1(n_484),
.B2(n_502),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_563),
.A2(n_388),
.B1(n_510),
.B2(n_493),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_616),
.B(n_588),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_626),
.B(n_589),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_627),
.B(n_566),
.Y(n_648)
);

NAND4xp25_ASAP7_75t_L g649 ( 
.A(n_637),
.B(n_606),
.C(n_583),
.D(n_566),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_620),
.B(n_583),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_613),
.B(n_569),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_619),
.B(n_569),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_613),
.B(n_643),
.Y(n_653)
);

NAND3xp33_ASAP7_75t_L g654 ( 
.A(n_636),
.B(n_577),
.C(n_569),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_622),
.B(n_569),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_624),
.A2(n_577),
.B1(n_510),
.B2(n_478),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_609),
.A2(n_577),
.B1(n_510),
.B2(n_576),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_611),
.B(n_577),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_611),
.B(n_584),
.Y(n_659)
);

NAND3xp33_ASAP7_75t_L g660 ( 
.A(n_612),
.B(n_510),
.C(n_502),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_639),
.B(n_576),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_621),
.B(n_576),
.Y(n_662)
);

NAND3xp33_ASAP7_75t_L g663 ( 
.A(n_610),
.B(n_502),
.C(n_490),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_621),
.B(n_51),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_638),
.B(n_52),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_SL g666 ( 
.A1(n_645),
.A2(n_53),
.B(n_55),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_621),
.B(n_56),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_630),
.B(n_60),
.Y(n_668)
);

AOI21xp33_ASAP7_75t_L g669 ( 
.A1(n_615),
.A2(n_502),
.B(n_490),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_644),
.B(n_502),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_623),
.B(n_61),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_618),
.B(n_64),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_631),
.B(n_65),
.Y(n_673)
);

OAI221xp5_ASAP7_75t_L g674 ( 
.A1(n_645),
.A2(n_502),
.B1(n_366),
.B2(n_362),
.C(n_69),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_614),
.B(n_66),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_646),
.B(n_67),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_655),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_647),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_661),
.B(n_640),
.Y(n_679)
);

NOR3xp33_ASAP7_75t_L g680 ( 
.A(n_653),
.B(n_632),
.C(n_633),
.Y(n_680)
);

NAND3xp33_ASAP7_75t_L g681 ( 
.A(n_653),
.B(n_628),
.C(n_641),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_650),
.B(n_68),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_659),
.A2(n_617),
.B1(n_634),
.B2(n_625),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_662),
.B(n_642),
.Y(n_684)
);

NAND3xp33_ASAP7_75t_L g685 ( 
.A(n_665),
.B(n_635),
.C(n_629),
.Y(n_685)
);

AOI211xp5_ASAP7_75t_L g686 ( 
.A1(n_659),
.A2(n_71),
.B(n_73),
.C(n_74),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_675),
.A2(n_366),
.B1(n_362),
.B2(n_81),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_648),
.Y(n_688)
);

OAI21xp33_ASAP7_75t_L g689 ( 
.A1(n_649),
.A2(n_366),
.B(n_362),
.Y(n_689)
);

AND4x1_ASAP7_75t_L g690 ( 
.A(n_663),
.B(n_75),
.C(n_79),
.D(n_82),
.Y(n_690)
);

NAND3xp33_ASAP7_75t_L g691 ( 
.A(n_654),
.B(n_203),
.C(n_85),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_678),
.Y(n_692)
);

NAND4xp75_ASAP7_75t_SL g693 ( 
.A(n_676),
.B(n_662),
.C(n_675),
.D(n_668),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_688),
.B(n_652),
.Y(n_694)
);

NOR4xp25_ASAP7_75t_L g695 ( 
.A(n_681),
.B(n_651),
.C(n_666),
.D(n_660),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_677),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_684),
.Y(n_697)
);

NAND4xp75_ASAP7_75t_L g698 ( 
.A(n_682),
.B(n_651),
.C(n_670),
.D(n_672),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_684),
.B(n_667),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_679),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_680),
.B(n_664),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_697),
.B(n_680),
.Y(n_702)
);

XOR2x2_ASAP7_75t_L g703 ( 
.A(n_693),
.B(n_686),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_692),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_701),
.B(n_689),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_700),
.B(n_683),
.Y(n_706)
);

OA22x2_ASAP7_75t_L g707 ( 
.A1(n_706),
.A2(n_700),
.B1(n_697),
.B2(n_696),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_704),
.Y(n_708)
);

OA22x2_ASAP7_75t_L g709 ( 
.A1(n_706),
.A2(n_700),
.B1(n_699),
.B2(n_694),
.Y(n_709)
);

AOI22x1_ASAP7_75t_L g710 ( 
.A1(n_702),
.A2(n_701),
.B1(n_703),
.B2(n_695),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_705),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_702),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_708),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_711),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_712),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_707),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_709),
.Y(n_717)
);

OAI322xp33_ASAP7_75t_L g718 ( 
.A1(n_716),
.A2(n_710),
.A3(n_685),
.B1(n_691),
.B2(n_674),
.C1(n_670),
.C2(n_658),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_715),
.A2(n_710),
.B1(n_698),
.B2(n_687),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_713),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_719),
.A2(n_717),
.B1(n_715),
.B2(n_714),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_SL g722 ( 
.A1(n_720),
.A2(n_687),
.B(n_671),
.C(n_673),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_718),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_719),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_721),
.Y(n_725)
);

NOR4xp25_ASAP7_75t_L g726 ( 
.A(n_723),
.B(n_656),
.C(n_669),
.D(n_657),
.Y(n_726)
);

NOR4xp25_ASAP7_75t_L g727 ( 
.A(n_724),
.B(n_690),
.C(n_86),
.D(n_89),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_722),
.Y(n_728)
);

AOI221xp5_ASAP7_75t_L g729 ( 
.A1(n_723),
.A2(n_84),
.B1(n_90),
.B2(n_91),
.C(n_94),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_721),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_725),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_730),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_728),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_727),
.B(n_203),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_726),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_729),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_732),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_735),
.A2(n_203),
.B1(n_97),
.B2(n_98),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_731),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_733),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_733),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_736),
.Y(n_742)
);

NOR2x1_ASAP7_75t_L g743 ( 
.A(n_734),
.B(n_96),
.Y(n_743)
);

NAND4xp25_ASAP7_75t_L g744 ( 
.A(n_731),
.B(n_99),
.C(n_101),
.D(n_104),
.Y(n_744)
);

AOI22xp5_ASAP7_75t_L g745 ( 
.A1(n_735),
.A2(n_203),
.B1(n_106),
.B2(n_107),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_741),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_739),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_742),
.A2(n_203),
.B1(n_110),
.B2(n_111),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_737),
.B(n_105),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_740),
.B(n_743),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_745),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_744),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_738),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_746),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_754)
);

OAI22x1_ASAP7_75t_L g755 ( 
.A1(n_747),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_750),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_753),
.A2(n_752),
.B1(n_751),
.B2(n_748),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_749),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_756),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_757),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_760),
.A2(n_753),
.B1(n_758),
.B2(n_755),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_759),
.A2(n_754),
.B1(n_123),
.B2(n_124),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_761),
.Y(n_763)
);

AO22x1_ASAP7_75t_L g764 ( 
.A1(n_763),
.A2(n_762),
.B1(n_125),
.B2(n_126),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_764),
.Y(n_765)
);

AOI221xp5_ASAP7_75t_L g766 ( 
.A1(n_765),
.A2(n_121),
.B1(n_130),
.B2(n_131),
.C(n_132),
.Y(n_766)
);

AOI211xp5_ASAP7_75t_L g767 ( 
.A1(n_766),
.A2(n_134),
.B(n_135),
.C(n_136),
.Y(n_767)
);


endmodule