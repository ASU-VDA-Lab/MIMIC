module fake_jpeg_4729_n_317 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_16),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_29),
.B1(n_33),
.B2(n_25),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_27),
.Y(n_46)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_34),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_46),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_47),
.Y(n_84)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_60),
.B1(n_32),
.B2(n_22),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_52),
.Y(n_94)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_32),
.C(n_27),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_35),
.A2(n_29),
.B1(n_33),
.B2(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_34),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_18),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_26),
.Y(n_90)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_67),
.Y(n_88)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_58),
.A2(n_33),
.B1(n_29),
.B2(n_19),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_85),
.B1(n_92),
.B2(n_56),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_32),
.C(n_19),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_26),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_86),
.B1(n_96),
.B2(n_51),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_31),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_83),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_32),
.B1(n_20),
.B2(n_23),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_81),
.B1(n_51),
.B2(n_56),
.Y(n_108)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_49),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_18),
.B1(n_21),
.B2(n_30),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_31),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_32),
.B1(n_21),
.B2(n_30),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_22),
.B(n_31),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_83),
.B(n_90),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_12),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_23),
.B1(n_20),
.B2(n_31),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_55),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_97),
.A2(n_98),
.B1(n_108),
.B2(n_88),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_69),
.B1(n_68),
.B2(n_67),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_101),
.B(n_106),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_74),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_104),
.Y(n_131)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_47),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_107),
.B(n_112),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_69),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_76),
.B1(n_71),
.B2(n_92),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_94),
.B1(n_80),
.B2(n_73),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_70),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_54),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_116),
.A2(n_93),
.B(n_91),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_120),
.Y(n_151)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_119),
.A2(n_121),
.B1(n_123),
.B2(n_72),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_49),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_89),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_31),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_88),
.Y(n_147)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_125),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_90),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_130),
.Y(n_162)
);

AO21x2_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_84),
.B(n_23),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_128),
.A2(n_144),
.B1(n_150),
.B2(n_107),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_129),
.B(n_97),
.Y(n_183)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_84),
.B(n_49),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_135),
.Y(n_163)
);

NAND2x1p5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_26),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_133),
.A2(n_116),
.B(n_114),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_139),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_94),
.C(n_93),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_97),
.C(n_26),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_73),
.B1(n_91),
.B2(n_23),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_143),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_104),
.A2(n_88),
.B1(n_65),
.B2(n_11),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_102),
.Y(n_153)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_148),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_65),
.B1(n_20),
.B2(n_26),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_65),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_157),
.C(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_131),
.B(n_111),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_156),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_109),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_102),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_158),
.B(n_161),
.Y(n_189)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_167),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_112),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_170),
.Y(n_190)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_125),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_183),
.Y(n_203)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_176),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_173),
.B1(n_170),
.B2(n_161),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_134),
.A2(n_110),
.B1(n_105),
.B2(n_151),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_122),
.B(n_120),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_179),
.B(n_142),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_152),
.B(n_101),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_132),
.B(n_98),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_130),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_155),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_158),
.B(n_142),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_185),
.B(n_193),
.Y(n_221)
);

FAx1_ASAP7_75t_SL g214 ( 
.A(n_186),
.B(n_183),
.CI(n_174),
.CON(n_214),
.SN(n_214)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_163),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_194),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_166),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_157),
.C(n_168),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_198),
.C(n_210),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_147),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_154),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_202),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_210),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_176),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_162),
.B1(n_182),
.B2(n_178),
.Y(n_204)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_97),
.B1(n_128),
.B2(n_145),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_159),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_138),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_156),
.B(n_128),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_211),
.A2(n_197),
.B(n_1),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_216),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_197),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_155),
.B(n_160),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_218),
.A2(n_227),
.B(n_233),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_181),
.C(n_179),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_228),
.C(n_235),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_177),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_232),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_195),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_230),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_213),
.Y(n_236)
);

AO21x1_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_165),
.B(n_145),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_137),
.C(n_135),
.Y(n_228)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_199),
.B(n_164),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_124),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_208),
.B(n_159),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_99),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_193),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_138),
.C(n_99),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_243),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_205),
.B1(n_190),
.B2(n_194),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_239),
.Y(n_259)
);

OAI221xp5_ASAP7_75t_SL g240 ( 
.A1(n_226),
.A2(n_188),
.B1(n_190),
.B2(n_200),
.C(n_201),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_240),
.B(n_223),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_186),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_201),
.B(n_184),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_244),
.A2(n_255),
.B(n_227),
.Y(n_263)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_220),
.A2(n_204),
.B1(n_206),
.B2(n_189),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_253),
.B1(n_8),
.B2(n_15),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_188),
.C(n_208),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_219),
.C(n_228),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_211),
.A2(n_225),
.B1(n_214),
.B2(n_232),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_0),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_254),
.C(n_253),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_260),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_235),
.C(n_218),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_262),
.C(n_264),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_221),
.C(n_215),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_263),
.A2(n_265),
.B(n_267),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_231),
.C(n_212),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_249),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_244),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_99),
.C(n_20),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_242),
.C(n_248),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_246),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_271),
.B(n_241),
.Y(n_280)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_274),
.C(n_281),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_256),
.A2(n_245),
.B1(n_238),
.B2(n_252),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_276),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_280),
.Y(n_288)
);

A2O1A1O1Ixp25_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_255),
.B(n_243),
.C(n_236),
.D(n_252),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_279),
.B(n_284),
.Y(n_285)
);

AOI21x1_ASAP7_75t_SL g282 ( 
.A1(n_263),
.A2(n_270),
.B(n_262),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_261),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_0),
.C(n_1),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_11),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_7),
.C(n_14),
.Y(n_284)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_282),
.A2(n_268),
.B1(n_258),
.B2(n_259),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_14),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_257),
.B1(n_269),
.B2(n_10),
.Y(n_291)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_287),
.A3(n_285),
.B1(n_294),
.B2(n_273),
.C1(n_283),
.C2(n_286),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_16),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_292),
.A2(n_293),
.B(n_294),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

NOR2x1_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_0),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_295),
.A2(n_278),
.B(n_10),
.Y(n_298)
);

OAI31xp33_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_301),
.A3(n_302),
.B(n_2),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_300),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_272),
.A3(n_278),
.B1(n_16),
.B2(n_14),
.C1(n_13),
.C2(n_12),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_304),
.C(n_303),
.Y(n_305)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_13),
.B(n_1),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_289),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_292),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_310),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_2),
.B(n_4),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_306),
.A2(n_308),
.B(n_309),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_296),
.A2(n_2),
.B(n_4),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_6),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_307),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_311),
.B(n_307),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_312),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_313),
.B(n_5),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_4),
.Y(n_317)
);


endmodule