module fake_jpeg_20542_n_289 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_289);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_14;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_10),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx24_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_10),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_20),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_32),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_20),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_33),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_23),
.B1(n_13),
.B2(n_16),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_26),
.B1(n_13),
.B2(n_32),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_26),
.B(n_13),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_31),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_49),
.B(n_55),
.C(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_47),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_43),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_25),
.B1(n_30),
.B2(n_32),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_40),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_40),
.B1(n_32),
.B2(n_25),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_32),
.B1(n_30),
.B2(n_25),
.Y(n_55)
);

AND2x4_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_40),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_27),
.B(n_29),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_40),
.B(n_43),
.Y(n_78)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_68),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_69),
.B(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_70),
.B(n_43),
.Y(n_87)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_43),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_78),
.Y(n_80)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_47),
.B1(n_56),
.B2(n_49),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_86),
.B1(n_88),
.B2(n_73),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_93),
.Y(n_115)
);

AND2x4_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_59),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_89),
.B(n_37),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_56),
.B1(n_54),
.B2(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_87),
.B(n_94),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_45),
.B1(n_77),
.B2(n_71),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_44),
.B(n_54),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_69),
.B(n_33),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_76),
.B(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_37),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_19),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_98),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_40),
.Y(n_98)
);

AOI22x1_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_72),
.B1(n_78),
.B2(n_68),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_31),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_100),
.B(n_107),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_83),
.A2(n_72),
.B1(n_66),
.B2(n_62),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_101),
.A2(n_102),
.B1(n_120),
.B2(n_24),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_37),
.B1(n_65),
.B2(n_67),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_111),
.B1(n_84),
.B2(n_80),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_61),
.B(n_65),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_104),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_110),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_63),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_67),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_113),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_19),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_30),
.B1(n_36),
.B2(n_24),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_53),
.Y(n_113)
);

INVxp33_ASAP7_75t_SL g114 ( 
.A(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_85),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_91),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_13),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_42),
.B1(n_24),
.B2(n_28),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_96),
.B(n_20),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_31),
.Y(n_144)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_112),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_130),
.B(n_136),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_99),
.A2(n_84),
.B1(n_96),
.B2(n_95),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_109),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_42),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_147),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_110),
.B(n_16),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_140),
.B(n_16),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_23),
.B1(n_42),
.B2(n_22),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_150),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_142),
.B(n_144),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_143),
.A2(n_116),
.B1(n_51),
.B2(n_46),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_31),
.Y(n_166)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_149),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_42),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_24),
.C(n_28),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_39),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_21),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_23),
.B1(n_22),
.B2(n_11),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_11),
.Y(n_156)
);

AO22x1_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_117),
.B1(n_45),
.B2(n_100),
.Y(n_152)
);

AO22x1_ASAP7_75t_L g196 ( 
.A1(n_152),
.A2(n_178),
.B1(n_158),
.B2(n_166),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_22),
.C(n_28),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_144),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_156),
.B(n_174),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_158),
.A2(n_51),
.B1(n_46),
.B2(n_45),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_159),
.B(n_173),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_53),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_169),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_53),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_172),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_166),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_146),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_53),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_53),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_15),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_175),
.B(n_177),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_15),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_179),
.Y(n_213)
);

XOR2x2_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_131),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_183),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_SL g183 ( 
.A1(n_171),
.A2(n_145),
.B(n_143),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_148),
.C(n_123),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_185),
.B(n_191),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_161),
.B(n_143),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_192),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_128),
.B(n_127),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_200),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_139),
.B(n_1),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_139),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_28),
.C(n_38),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_199),
.C(n_34),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_174),
.B(n_15),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_197),
.Y(n_215)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_15),
.Y(n_197)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_15),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_178),
.A2(n_34),
.B1(n_15),
.B2(n_18),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_180),
.C(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_208),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_182),
.A2(n_176),
.B1(n_166),
.B2(n_167),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_211),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_152),
.C(n_168),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_152),
.C(n_168),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_210),
.B(n_219),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_187),
.A2(n_167),
.B1(n_164),
.B2(n_170),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_193),
.A2(n_164),
.B1(n_170),
.B2(n_153),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_218),
.B1(n_184),
.B2(n_188),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_197),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_184),
.A2(n_34),
.B1(n_18),
.B2(n_14),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_34),
.C(n_18),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_34),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_39),
.Y(n_237)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_225),
.Y(n_246)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_228),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_189),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_233),
.Y(n_239)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_229),
.B(n_234),
.Y(n_240)
);

AO221x1_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_201),
.B1(n_190),
.B2(n_39),
.C(n_18),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_235),
.B(n_206),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_190),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_39),
.B1(n_14),
.B2(n_12),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_203),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_203),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_230),
.C(n_227),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_243),
.C(n_244),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_17),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_213),
.C(n_204),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_222),
.C(n_235),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_220),
.C(n_215),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_247),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_215),
.C(n_219),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_17),
.B(n_39),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_249),
.A2(n_246),
.B(n_1),
.Y(n_254)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_250),
.A2(n_14),
.B1(n_12),
.B2(n_2),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_4),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_248),
.A2(n_17),
.B(n_14),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_255),
.A2(n_260),
.B(n_3),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_0),
.B(n_2),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_259),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_240),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_12),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_261),
.B(n_5),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_0),
.B(n_2),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_262),
.A2(n_3),
.B(n_4),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_264),
.B(n_265),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_12),
.C(n_4),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_269),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_3),
.B(n_4),
.Y(n_268)
);

NAND2x1p5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_271),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_6),
.B(n_7),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_251),
.B1(n_257),
.B2(n_7),
.Y(n_273)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_273),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_5),
.C(n_6),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_275),
.A2(n_278),
.B(n_263),
.Y(n_282)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_277),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_6),
.B(n_7),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_282),
.B(n_279),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_283),
.A2(n_284),
.B(n_263),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_280),
.Y(n_284)
);

AO21x1_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_276),
.B(n_274),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_281),
.B(n_9),
.Y(n_287)
);

A2O1A1O1Ixp25_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_8),
.B(n_9),
.C(n_10),
.D(n_276),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_8),
.C(n_9),
.Y(n_289)
);


endmodule