module fake_jpeg_18908_n_66 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_66);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_66;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx16f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx5_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_20),
.Y(n_28)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_13),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_22),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_15),
.B(n_13),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_16),
.B1(n_10),
.B2(n_15),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_10),
.B1(n_17),
.B2(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_18),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_21),
.B(n_17),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_34),
.B(n_35),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_29),
.B1(n_26),
.B2(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_9),
.B(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_26),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_9),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_39),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_42),
.B1(n_43),
.B2(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_25),
.B1(n_14),
.B2(n_9),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_47),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_SL g49 ( 
.A(n_45),
.B(n_38),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_5),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_38),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_52),
.Y(n_57)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_42),
.C(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_58),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_47),
.C(n_39),
.Y(n_59)
);

AOI31xp67_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_56),
.A3(n_55),
.B(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_55),
.Y(n_62)
);

XOR2x2_ASAP7_75t_SL g64 ( 
.A(n_62),
.B(n_63),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_6),
.C(n_4),
.Y(n_63)
);

AOI321xp33_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_1),
.A3(n_6),
.B1(n_36),
.B2(n_44),
.C(n_60),
.Y(n_65)
);

BUFx24_ASAP7_75t_SL g66 ( 
.A(n_65),
.Y(n_66)
);


endmodule