module real_jpeg_28381_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_344, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_344;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_0),
.A2(n_27),
.B1(n_31),
.B2(n_37),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_0),
.A2(n_37),
.B1(n_58),
.B2(n_60),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_0),
.A2(n_37),
.B1(n_53),
.B2(n_54),
.Y(n_120)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_1),
.Y(n_94)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_1),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_1),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_2),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_2),
.A2(n_27),
.B1(n_31),
.B2(n_46),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_2),
.A2(n_46),
.B1(n_58),
.B2(n_60),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_3),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_3),
.A2(n_27),
.B1(n_31),
.B2(n_139),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_3),
.A2(n_53),
.B1(n_54),
.B2(n_139),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_3),
.A2(n_58),
.B1(n_60),
.B2(n_139),
.Y(n_251)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_5),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_5),
.A2(n_48),
.B1(n_58),
.B2(n_60),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_5),
.A2(n_27),
.B1(n_31),
.B2(n_48),
.Y(n_148)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_6),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_6),
.B(n_26),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_6),
.B(n_31),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g215 ( 
.A1(n_6),
.A2(n_31),
.B(n_211),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_6),
.A2(n_53),
.B1(n_54),
.B2(n_172),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_6),
.A2(n_55),
.B(n_58),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_6),
.B(n_77),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_6),
.A2(n_94),
.B1(n_115),
.B2(n_259),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_8),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_8),
.A2(n_27),
.B1(n_31),
.B2(n_111),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_111),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_8),
.A2(n_58),
.B1(n_60),
.B2(n_111),
.Y(n_246)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_10),
.A2(n_25),
.B1(n_53),
.B2(n_54),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_10),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_10),
.A2(n_25),
.B1(n_58),
.B2(n_60),
.Y(n_100)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_12),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_12),
.A2(n_27),
.B1(n_31),
.B2(n_174),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_174),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_12),
.A2(n_58),
.B1(n_60),
.B2(n_174),
.Y(n_259)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

INVx11_ASAP7_75t_SL g59 ( 
.A(n_15),
.Y(n_59)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_342),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_82),
.B(n_340),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_38),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_20),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_21),
.A2(n_44),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_22),
.A2(n_33),
.B(n_81),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_22),
.A2(n_26),
.B(n_33),
.Y(n_342)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_26),
.B(n_29),
.C(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_29),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g171 ( 
.A(n_23),
.B(n_172),
.CON(n_171),
.SN(n_171)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_26),
.A2(n_33),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_27),
.A2(n_31),
.B1(n_66),
.B2(n_68),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_27),
.A2(n_34),
.B1(n_171),
.B2(n_185),
.Y(n_184)
);

AOI32xp33_ASAP7_75t_L g209 ( 
.A1(n_27),
.A2(n_53),
.A3(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_209)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_29),
.B(n_31),
.Y(n_185)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_32),
.A2(n_45),
.B(n_49),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_33),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_36),
.B(n_49),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_39),
.B(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_74),
.C(n_79),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_40),
.A2(n_41),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_50),
.C(n_63),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_42),
.A2(n_43),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_44),
.A2(n_49),
.B1(n_110),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_44),
.A2(n_49),
.B1(n_138),
.B2(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_50),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_50),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_50),
.A2(n_63),
.B1(n_308),
.B2(n_322),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_57),
.B(n_61),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_51),
.A2(n_57),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_51),
.A2(n_103),
.B(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_51),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_51),
.A2(n_61),
.B(n_119),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_51),
.A2(n_57),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_51),
.A2(n_145),
.B(n_219),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_51),
.A2(n_57),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_51),
.A2(n_57),
.B1(n_218),
.B2(n_236),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_54),
.B1(n_66),
.B2(n_68),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_54),
.B(n_66),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_54),
.A2(n_56),
.B(n_172),
.C(n_238),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_57),
.A2(n_102),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_57),
.B(n_172),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_58),
.Y(n_60)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_60),
.B(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_62),
.B(n_121),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_63),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_70),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_64),
.A2(n_76),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_65),
.B(n_71),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_65),
.A2(n_72),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_65),
.A2(n_72),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_65),
.A2(n_72),
.B1(n_168),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_65),
.A2(n_72),
.B1(n_197),
.B2(n_215),
.Y(n_214)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_66),
.Y(n_210)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_70),
.A2(n_77),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_74),
.A2(n_75),
.B1(n_79),
.B2(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_78),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_76),
.A2(n_78),
.B(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_76),
.A2(n_135),
.B(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_79),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_333),
.B(n_339),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_303),
.A3(n_325),
.B1(n_331),
.B2(n_332),
.C(n_344),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_157),
.B(n_302),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_140),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_86),
.B(n_140),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_112),
.C(n_123),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_87),
.A2(n_88),
.B1(n_112),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_104),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_89),
.B(n_106),
.C(n_108),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_101),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_90),
.B(n_101),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_91),
.A2(n_187),
.B(n_188),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_92),
.A2(n_100),
.B(n_128),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_92),
.A2(n_98),
.B1(n_250),
.B2(n_252),
.Y(n_249)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_94),
.A2(n_115),
.B1(n_251),
.B2(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_94),
.B(n_172),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_97),
.A2(n_115),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

INVx5_ASAP7_75t_SL g116 ( 
.A(n_98),
.Y(n_116)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_98),
.Y(n_188)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_100),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_107),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_112),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_122),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_114),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_118),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g316 ( 
.A1(n_114),
.A2(n_151),
.B(n_154),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B(n_117),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_115),
.A2(n_126),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_118),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_120),
.B(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_123),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_134),
.C(n_136),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_124),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_131),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_131),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_134),
.A2(n_136),
.B1(n_137),
.B2(n_292),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_134),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_155),
.B2(n_156),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_150),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_143),
.B(n_150),
.C(n_156),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B(n_149),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_146),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_148),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_149),
.B(n_305),
.C(n_315),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_149),
.A2(n_305),
.B1(n_306),
.B2(n_330),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_149),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_155),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_296),
.B(n_301),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_201),
.B(n_282),
.C(n_295),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_189),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_160),
.B(n_189),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_175),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_162),
.B(n_163),
.C(n_175),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_170),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_170),
.B(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_173),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_183),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_177),
.B(n_181),
.C(n_183),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_186),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.C(n_195),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_190),
.A2(n_191),
.B1(n_277),
.B2(n_279),
.Y(n_276)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_195),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.C(n_200),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_200),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_281),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_274),
.B(n_280),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_229),
.B(n_273),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_220),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_205),
.B(n_220),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_213),
.C(n_216),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_206),
.A2(n_207),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_209),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_217),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_221),
.B(n_227),
.C(n_228),
.Y(n_275)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_267),
.B(n_272),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_247),
.B(n_266),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_239),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_232),
.B(n_239),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_237),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_245),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_244),
.C(n_245),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_246),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_255),
.B(n_265),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_253),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_260),
.B(n_264),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_257),
.B(n_258),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_275),
.B(n_276),
.Y(n_280)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_277),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_283),
.B(n_284),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_293),
.B2(n_294),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_290),
.C(n_294),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_317),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_317),
.Y(n_332)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.Y(n_306)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_307),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_310),
.C(n_312),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_312),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_312),
.A2(n_314),
.B1(n_319),
.B2(n_323),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_323),
.C(n_324),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_315),
.A2(n_316),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_324),
.Y(n_317)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_326),
.B(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_335),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_336),
.Y(n_338)
);


endmodule