module real_aes_6539_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_719;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g167 ( .A1(n_0), .A2(n_168), .B(n_169), .C(n_173), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_1), .B(n_162), .Y(n_175) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_3), .B(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_4), .A2(n_156), .B(n_470), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_5), .A2(n_136), .B(n_153), .C(n_514), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_6), .A2(n_156), .B(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_7), .B(n_162), .Y(n_476) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_8), .A2(n_128), .B(n_250), .Y(n_249) );
AND2x6_ASAP7_75t_L g153 ( .A(n_9), .B(n_154), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_10), .A2(n_136), .B(n_153), .C(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g567 ( .A(n_11), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_12), .B(n_40), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_13), .B(n_172), .Y(n_516) );
INVx1_ASAP7_75t_L g133 ( .A(n_14), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_15), .B(n_147), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_16), .A2(n_148), .B(n_525), .C(n_527), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_17), .B(n_162), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_18), .B(n_190), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_19), .A2(n_136), .B(n_182), .C(n_189), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_20), .A2(n_171), .B(n_224), .C(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_21), .B(n_172), .Y(n_498) );
AOI222xp33_ASAP7_75t_L g445 ( .A1(n_22), .A2(n_446), .B1(n_716), .B2(n_717), .C1(n_726), .C2(n_730), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_23), .B(n_172), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_24), .Y(n_494) );
INVx1_ASAP7_75t_L g464 ( .A(n_25), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_26), .A2(n_136), .B(n_189), .C(n_253), .Y(n_252) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_27), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_28), .Y(n_512) );
INVx1_ASAP7_75t_L g488 ( .A(n_29), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_30), .A2(n_156), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_31), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g138 ( .A(n_32), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_33), .A2(n_151), .B(n_205), .C(n_206), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_34), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_35), .A2(n_171), .B(n_473), .C(n_475), .Y(n_472) );
INVxp67_ASAP7_75t_L g489 ( .A(n_36), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_37), .B(n_255), .Y(n_254) );
CKINVDCx14_ASAP7_75t_R g471 ( .A(n_38), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_39), .A2(n_136), .B(n_189), .C(n_463), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g564 ( .A1(n_41), .A2(n_173), .B(n_565), .C(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_42), .B(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_43), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_44), .B(n_147), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_45), .B(n_156), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_46), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_47), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_48), .A2(n_151), .B(n_205), .C(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g170 ( .A(n_49), .Y(n_170) );
OAI22xp5_ASAP7_75t_SL g114 ( .A1(n_50), .A2(n_66), .B1(n_115), .B2(n_116), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_50), .Y(n_116) );
INVx1_ASAP7_75t_L g234 ( .A(n_51), .Y(n_234) );
INVx1_ASAP7_75t_L g532 ( .A(n_52), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_53), .B(n_156), .Y(n_231) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_54), .A2(n_71), .B1(n_119), .B2(n_120), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_54), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_55), .Y(n_194) );
CKINVDCx14_ASAP7_75t_R g563 ( .A(n_56), .Y(n_563) );
INVx1_ASAP7_75t_L g154 ( .A(n_57), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_58), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_59), .B(n_162), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_60), .A2(n_143), .B(n_188), .C(n_245), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_61), .A2(n_70), .B1(n_723), .B2(n_724), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_61), .Y(n_723) );
INVx1_ASAP7_75t_L g132 ( .A(n_62), .Y(n_132) );
INVx1_ASAP7_75t_SL g474 ( .A(n_63), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_64), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_65), .B(n_147), .Y(n_208) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_66), .A2(n_104), .B1(n_436), .B2(n_444), .C1(n_733), .C2(n_736), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_66), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_66), .B(n_162), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_67), .B(n_148), .Y(n_221) );
INVx1_ASAP7_75t_L g497 ( .A(n_68), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_69), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_70), .Y(n_724) );
INVx1_ASAP7_75t_L g120 ( .A(n_71), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_72), .B(n_184), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g135 ( .A1(n_73), .A2(n_136), .B(n_141), .C(n_151), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g243 ( .A(n_74), .Y(n_243) );
INVx1_ASAP7_75t_L g443 ( .A(n_75), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_76), .A2(n_156), .B(n_562), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_77), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_78), .A2(n_156), .B(n_522), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_79), .A2(n_180), .B(n_484), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_80), .Y(n_461) );
INVx1_ASAP7_75t_L g523 ( .A(n_81), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_82), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_82), .Y(n_720) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_83), .B(n_186), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_84), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_85), .A2(n_156), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g526 ( .A(n_86), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_87), .A2(n_718), .B1(n_719), .B2(n_725), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_87), .Y(n_718) );
INVx2_ASAP7_75t_L g130 ( .A(n_88), .Y(n_130) );
INVx1_ASAP7_75t_L g515 ( .A(n_89), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_90), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_91), .B(n_172), .Y(n_222) );
OR2x2_ASAP7_75t_L g108 ( .A(n_92), .B(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g450 ( .A(n_92), .B(n_110), .Y(n_450) );
INVx2_ASAP7_75t_L g715 ( .A(n_92), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_93), .A2(n_136), .B(n_151), .C(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_94), .B(n_156), .Y(n_203) );
INVx1_ASAP7_75t_L g207 ( .A(n_95), .Y(n_207) );
INVxp67_ASAP7_75t_L g246 ( .A(n_96), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_97), .B(n_128), .Y(n_568) );
INVx1_ASAP7_75t_L g142 ( .A(n_98), .Y(n_142) );
INVx1_ASAP7_75t_L g217 ( .A(n_99), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_100), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g535 ( .A(n_101), .Y(n_535) );
AND2x2_ASAP7_75t_L g236 ( .A(n_102), .B(n_192), .Y(n_236) );
OAI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_113), .B(n_433), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NAND2xp33_ASAP7_75t_L g734 ( .A(n_106), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_108), .Y(n_435) );
BUFx2_ASAP7_75t_L g738 ( .A(n_108), .Y(n_738) );
NOR2x2_ASAP7_75t_L g732 ( .A(n_109), .B(n_715), .Y(n_732) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g714 ( .A(n_110), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AOI22xp33_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_117), .B1(n_431), .B2(n_432), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_114), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_117), .Y(n_432) );
XNOR2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_121), .Y(n_117) );
INVx1_ASAP7_75t_L g447 ( .A(n_121), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_121), .A2(n_452), .B1(n_727), .B2(n_728), .Y(n_726) );
OR3x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_339), .C(n_388), .Y(n_121) );
NAND5xp2_ASAP7_75t_L g122 ( .A(n_123), .B(n_273), .C(n_302), .D(n_310), .E(n_325), .Y(n_122) );
O2A1O1Ixp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_196), .B(n_212), .C(n_257), .Y(n_123) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_176), .Y(n_124) );
AND2x2_ASAP7_75t_L g268 ( .A(n_125), .B(n_265), .Y(n_268) );
AND2x2_ASAP7_75t_L g301 ( .A(n_125), .B(n_177), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_125), .B(n_200), .Y(n_394) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_161), .Y(n_125) );
INVx2_ASAP7_75t_L g199 ( .A(n_126), .Y(n_199) );
BUFx2_ASAP7_75t_L g368 ( .A(n_126), .Y(n_368) );
AO21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_134), .B(n_159), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_127), .B(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g162 ( .A(n_127), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_127), .B(n_211), .Y(n_210) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_127), .A2(n_216), .B(n_226), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_127), .B(n_467), .Y(n_466) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_127), .A2(n_493), .B(n_500), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_127), .B(n_518), .Y(n_517) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_128), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_128), .A2(n_251), .B(n_252), .Y(n_250) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g228 ( .A(n_129), .Y(n_228) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g192 ( .A(n_130), .B(n_131), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_155), .Y(n_134) );
INVx5_ASAP7_75t_L g166 ( .A(n_136), .Y(n_166) );
AND2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
BUFx3_ASAP7_75t_L g174 ( .A(n_137), .Y(n_174) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g158 ( .A(n_138), .Y(n_158) );
INVx1_ASAP7_75t_L g225 ( .A(n_138), .Y(n_225) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_140), .Y(n_145) );
INVx3_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
AND2x2_ASAP7_75t_L g157 ( .A(n_140), .B(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_140), .Y(n_172) );
INVx1_ASAP7_75t_L g255 ( .A(n_140), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_146), .C(n_149), .Y(n_141) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_144), .A2(n_147), .B1(n_488), .B2(n_489), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_144), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_144), .B(n_535), .Y(n_534) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g184 ( .A(n_145), .Y(n_184) );
INVx2_ASAP7_75t_L g168 ( .A(n_147), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_147), .B(n_246), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_147), .A2(n_187), .B(n_464), .C(n_465), .Y(n_463) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_148), .B(n_567), .Y(n_566) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g475 ( .A(n_150), .Y(n_475) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_SL g164 ( .A1(n_152), .A2(n_165), .B(n_166), .C(n_167), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_152), .A2(n_166), .B(n_243), .C(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_152), .A2(n_166), .B(n_471), .C(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_152), .A2(n_166), .B(n_485), .C(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_152), .A2(n_166), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_SL g531 ( .A1(n_152), .A2(n_166), .B(n_532), .C(n_533), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_SL g562 ( .A1(n_152), .A2(n_166), .B(n_563), .C(n_564), .Y(n_562) );
INVx4_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g156 ( .A(n_153), .B(n_157), .Y(n_156) );
BUFx3_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
NAND2x1p5_ASAP7_75t_L g218 ( .A(n_153), .B(n_157), .Y(n_218) );
BUFx2_ASAP7_75t_L g180 ( .A(n_156), .Y(n_180) );
INVx1_ASAP7_75t_L g188 ( .A(n_158), .Y(n_188) );
AND2x2_ASAP7_75t_L g176 ( .A(n_161), .B(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g266 ( .A(n_161), .Y(n_266) );
AND2x2_ASAP7_75t_L g352 ( .A(n_161), .B(n_265), .Y(n_352) );
AND2x2_ASAP7_75t_L g407 ( .A(n_161), .B(n_199), .Y(n_407) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_175), .Y(n_161) );
INVx2_ASAP7_75t_L g205 ( .A(n_166), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_171), .B(n_474), .Y(n_473) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g565 ( .A(n_172), .Y(n_565) );
INVx2_ASAP7_75t_L g499 ( .A(n_173), .Y(n_499) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_174), .Y(n_209) );
INVx1_ASAP7_75t_L g527 ( .A(n_174), .Y(n_527) );
INVx1_ASAP7_75t_L g324 ( .A(n_176), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_176), .B(n_200), .Y(n_371) );
INVx5_ASAP7_75t_L g265 ( .A(n_177), .Y(n_265) );
AND2x4_ASAP7_75t_L g286 ( .A(n_177), .B(n_266), .Y(n_286) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_177), .Y(n_308) );
AND2x2_ASAP7_75t_L g383 ( .A(n_177), .B(n_368), .Y(n_383) );
AND2x2_ASAP7_75t_L g386 ( .A(n_177), .B(n_201), .Y(n_386) );
OR2x6_ASAP7_75t_L g177 ( .A(n_178), .B(n_193), .Y(n_177) );
AOI21xp5_ASAP7_75t_SL g178 ( .A1(n_179), .A2(n_181), .B(n_190), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_185), .B(n_187), .Y(n_182) );
INVx2_ASAP7_75t_L g186 ( .A(n_184), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_186), .A2(n_207), .B(n_208), .C(n_209), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_186), .A2(n_209), .B(n_234), .C(n_235), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_186), .A2(n_497), .B(n_498), .C(n_499), .Y(n_496) );
O2A1O1Ixp5_ASAP7_75t_L g514 ( .A1(n_186), .A2(n_499), .B(n_515), .C(n_516), .Y(n_514) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_188), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_191), .B(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g195 ( .A(n_192), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_192), .A2(n_203), .B(n_204), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_192), .A2(n_231), .B(n_232), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_192), .A2(n_218), .B(n_461), .C(n_462), .Y(n_460) );
OA21x2_ASAP7_75t_L g560 ( .A1(n_192), .A2(n_561), .B(n_568), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_195), .A2(n_511), .B(n_517), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_196), .B(n_266), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_196), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_200), .Y(n_197) );
AND2x2_ASAP7_75t_L g291 ( .A(n_198), .B(n_266), .Y(n_291) );
AND2x2_ASAP7_75t_L g309 ( .A(n_198), .B(n_201), .Y(n_309) );
INVx1_ASAP7_75t_L g329 ( .A(n_198), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_198), .B(n_265), .Y(n_374) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_198), .Y(n_416) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_199), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_200), .B(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_200), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_200), .A2(n_261), .B(n_322), .C(n_324), .Y(n_321) );
AND2x2_ASAP7_75t_L g328 ( .A(n_200), .B(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g337 ( .A(n_200), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g341 ( .A(n_200), .B(n_265), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_200), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g356 ( .A(n_200), .B(n_266), .Y(n_356) );
AND2x2_ASAP7_75t_L g406 ( .A(n_200), .B(n_407), .Y(n_406) );
INVx5_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
BUFx2_ASAP7_75t_L g270 ( .A(n_201), .Y(n_270) );
AND2x2_ASAP7_75t_L g311 ( .A(n_201), .B(n_264), .Y(n_311) );
AND2x2_ASAP7_75t_L g323 ( .A(n_201), .B(n_298), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_201), .B(n_352), .Y(n_370) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_210), .Y(n_201) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_237), .Y(n_212) );
INVx1_ASAP7_75t_L g259 ( .A(n_213), .Y(n_259) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_229), .Y(n_213) );
OR2x2_ASAP7_75t_L g261 ( .A(n_214), .B(n_229), .Y(n_261) );
NAND3xp33_ASAP7_75t_L g267 ( .A(n_214), .B(n_268), .C(n_269), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_214), .B(n_239), .Y(n_278) );
OR2x2_ASAP7_75t_L g293 ( .A(n_214), .B(n_281), .Y(n_293) );
AND2x2_ASAP7_75t_L g299 ( .A(n_214), .B(n_248), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_214), .B(n_430), .Y(n_429) );
INVx5_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_215), .B(n_239), .Y(n_296) );
AND2x2_ASAP7_75t_L g335 ( .A(n_215), .B(n_249), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_215), .B(n_248), .Y(n_363) );
OR2x2_ASAP7_75t_L g366 ( .A(n_215), .B(n_248), .Y(n_366) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_219), .Y(n_216) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_218), .A2(n_494), .B(n_495), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_218), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_223), .A2(n_254), .B(n_256), .Y(n_253) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g482 ( .A(n_228), .Y(n_482) );
INVx5_ASAP7_75t_SL g281 ( .A(n_229), .Y(n_281) );
OR2x2_ASAP7_75t_L g287 ( .A(n_229), .B(n_238), .Y(n_287) );
AND2x2_ASAP7_75t_L g303 ( .A(n_229), .B(n_304), .Y(n_303) );
AOI321xp33_ASAP7_75t_L g310 ( .A1(n_229), .A2(n_311), .A3(n_312), .B1(n_313), .B2(n_319), .C(n_321), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_229), .B(n_237), .Y(n_320) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_229), .Y(n_333) );
OR2x2_ASAP7_75t_L g380 ( .A(n_229), .B(n_278), .Y(n_380) );
AND2x2_ASAP7_75t_L g402 ( .A(n_229), .B(n_299), .Y(n_402) );
AND2x2_ASAP7_75t_L g421 ( .A(n_229), .B(n_239), .Y(n_421) );
OR2x6_ASAP7_75t_L g229 ( .A(n_230), .B(n_236), .Y(n_229) );
INVx1_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_248), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_239), .B(n_248), .Y(n_262) );
AND2x2_ASAP7_75t_L g271 ( .A(n_239), .B(n_272), .Y(n_271) );
INVx3_ASAP7_75t_L g298 ( .A(n_239), .Y(n_298) );
AND2x2_ASAP7_75t_L g304 ( .A(n_239), .B(n_299), .Y(n_304) );
INVxp67_ASAP7_75t_L g334 ( .A(n_239), .Y(n_334) );
OR2x2_ASAP7_75t_L g376 ( .A(n_239), .B(n_281), .Y(n_376) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_247), .Y(n_239) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_240), .A2(n_469), .B(n_476), .Y(n_468) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_240), .A2(n_521), .B(n_528), .Y(n_520) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_240), .A2(n_530), .B(n_536), .Y(n_529) );
OR2x2_ASAP7_75t_L g258 ( .A(n_248), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_SL g272 ( .A(n_248), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_248), .B(n_261), .Y(n_305) );
AND2x2_ASAP7_75t_L g354 ( .A(n_248), .B(n_298), .Y(n_354) );
AND2x2_ASAP7_75t_L g392 ( .A(n_248), .B(n_281), .Y(n_392) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_249), .B(n_281), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_260), .B(n_263), .C(n_267), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_258), .A2(n_260), .B1(n_385), .B2(n_387), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_260), .A2(n_283), .B1(n_338), .B2(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx1_ASAP7_75t_SL g412 ( .A(n_261), .Y(n_412) );
INVx1_ASAP7_75t_SL g312 ( .A(n_262), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_264), .B(n_284), .Y(n_314) );
AOI222xp33_ASAP7_75t_L g325 ( .A1(n_264), .A2(n_305), .B1(n_312), .B2(n_326), .C1(n_330), .C2(n_336), .Y(n_325) );
AND2x2_ASAP7_75t_L g415 ( .A(n_264), .B(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g290 ( .A(n_265), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_265), .B(n_285), .Y(n_360) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_265), .Y(n_397) );
AND2x2_ASAP7_75t_L g400 ( .A(n_265), .B(n_309), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_265), .B(n_416), .Y(n_426) );
INVx1_ASAP7_75t_L g317 ( .A(n_266), .Y(n_317) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_266), .Y(n_345) );
O2A1O1Ixp33_ASAP7_75t_L g408 ( .A1(n_268), .A2(n_409), .B(n_410), .C(n_413), .Y(n_408) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND3xp33_ASAP7_75t_L g331 ( .A(n_270), .B(n_332), .C(n_335), .Y(n_331) );
OR2x2_ASAP7_75t_L g359 ( .A(n_270), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_270), .B(n_286), .Y(n_387) );
OR2x2_ASAP7_75t_L g292 ( .A(n_272), .B(n_293), .Y(n_292) );
AOI211xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_276), .B(n_282), .C(n_294), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_275), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g381 ( .A(n_276), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_279), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_277), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g295 ( .A(n_280), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_281), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g349 ( .A(n_281), .B(n_299), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_281), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_281), .B(n_298), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_287), .B1(n_288), .B2(n_292), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_284), .B(n_356), .Y(n_355) );
BUFx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_286), .B(n_328), .Y(n_327) );
OAI221xp5_ASAP7_75t_SL g350 ( .A1(n_287), .A2(n_351), .B1(n_353), .B2(n_355), .C(n_357), .Y(n_350) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AND2x2_ASAP7_75t_L g405 ( .A(n_290), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g418 ( .A(n_290), .B(n_407), .Y(n_418) );
INVx1_ASAP7_75t_L g338 ( .A(n_291), .Y(n_338) );
INVx1_ASAP7_75t_L g409 ( .A(n_292), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_293), .A2(n_376), .B(n_399), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_297), .B(n_300), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OAI21xp5_ASAP7_75t_SL g302 ( .A1(n_303), .A2(n_305), .B(n_306), .Y(n_302) );
INVx1_ASAP7_75t_L g342 ( .A(n_303), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_304), .A2(n_390), .B1(n_393), .B2(n_395), .C(n_398), .Y(n_389) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_312), .A2(n_402), .B1(n_403), .B2(n_405), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g378 ( .A(n_314), .Y(n_378) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2xp67_ASAP7_75t_SL g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g382 ( .A(n_318), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g347 ( .A(n_323), .Y(n_347) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_328), .B(n_352), .Y(n_404) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_334), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g420 ( .A(n_335), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g427 ( .A(n_335), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI211xp5_ASAP7_75t_SL g339 ( .A1(n_340), .A2(n_342), .B(n_343), .C(n_377), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI211xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_346), .B(n_350), .C(n_369), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_SL g430 ( .A(n_354), .Y(n_430) );
AND2x2_ASAP7_75t_L g367 ( .A(n_356), .B(n_368), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_361), .B1(n_365), .B2(n_367), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
OR2x2_ASAP7_75t_L g375 ( .A(n_363), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g428 ( .A(n_364), .Y(n_428) );
INVxp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI31xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .A3(n_372), .B(n_375), .Y(n_369) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI211xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B(n_381), .C(n_384), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
CKINVDCx16_ASAP7_75t_R g385 ( .A(n_386), .Y(n_385) );
NAND5xp2_ASAP7_75t_L g388 ( .A(n_389), .B(n_401), .C(n_408), .D(n_422), .E(n_425), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_400), .A2(n_426), .B1(n_427), .B2(n_429), .Y(n_425) );
INVx1_ASAP7_75t_SL g424 ( .A(n_402), .Y(n_424) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI21xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_417), .B(n_419), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_SL g735 ( .A(n_440), .B(n_442), .Y(n_735) );
OA21x2_ASAP7_75t_L g737 ( .A1(n_440), .A2(n_441), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVxp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_447), .A2(n_448), .B1(n_451), .B2(n_714), .Y(n_446) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g727 ( .A(n_449), .Y(n_727) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR3x1_ASAP7_75t_L g452 ( .A(n_453), .B(n_625), .C(n_672), .Y(n_452) );
NAND3xp33_ASAP7_75t_SL g453 ( .A(n_454), .B(n_571), .C(n_596), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_509), .B1(n_537), .B2(n_540), .C(n_548), .Y(n_454) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_477), .B(n_502), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_457), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_457), .B(n_553), .Y(n_669) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_468), .Y(n_457) );
AND2x2_ASAP7_75t_L g539 ( .A(n_458), .B(n_508), .Y(n_539) );
AND2x2_ASAP7_75t_L g589 ( .A(n_458), .B(n_507), .Y(n_589) );
AND2x2_ASAP7_75t_L g610 ( .A(n_458), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g615 ( .A(n_458), .B(n_582), .Y(n_615) );
OR2x2_ASAP7_75t_L g623 ( .A(n_458), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g695 ( .A(n_458), .B(n_491), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_458), .B(n_644), .Y(n_709) );
INVx3_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g554 ( .A(n_459), .B(n_468), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_459), .B(n_491), .Y(n_555) );
AND2x4_ASAP7_75t_L g577 ( .A(n_459), .B(n_508), .Y(n_577) );
AND2x2_ASAP7_75t_L g607 ( .A(n_459), .B(n_479), .Y(n_607) );
AND2x2_ASAP7_75t_L g616 ( .A(n_459), .B(n_606), .Y(n_616) );
AND2x2_ASAP7_75t_L g632 ( .A(n_459), .B(n_492), .Y(n_632) );
OR2x2_ASAP7_75t_L g641 ( .A(n_459), .B(n_624), .Y(n_641) );
AND2x2_ASAP7_75t_L g647 ( .A(n_459), .B(n_582), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_459), .B(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g661 ( .A(n_459), .B(n_504), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_459), .B(n_550), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_459), .B(n_611), .Y(n_700) );
OR2x6_ASAP7_75t_L g459 ( .A(n_460), .B(n_466), .Y(n_459) );
INVx2_ASAP7_75t_L g508 ( .A(n_468), .Y(n_508) );
AND2x2_ASAP7_75t_L g606 ( .A(n_468), .B(n_491), .Y(n_606) );
AND2x2_ASAP7_75t_L g611 ( .A(n_468), .B(n_492), .Y(n_611) );
INVx1_ASAP7_75t_L g667 ( .A(n_468), .Y(n_667) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g576 ( .A(n_478), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_491), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_479), .B(n_539), .Y(n_538) );
BUFx3_ASAP7_75t_L g553 ( .A(n_479), .Y(n_553) );
OR2x2_ASAP7_75t_L g624 ( .A(n_479), .B(n_491), .Y(n_624) );
OR2x2_ASAP7_75t_L g685 ( .A(n_479), .B(n_592), .Y(n_685) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_483), .B(n_490), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_481), .A2(n_505), .B(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g505 ( .A(n_483), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_490), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_491), .B(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g644 ( .A(n_491), .B(n_504), .Y(n_644) );
INVx2_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
BUFx2_ASAP7_75t_L g583 ( .A(n_492), .Y(n_583) );
INVx1_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_503), .A2(n_689), .B1(n_693), .B2(n_696), .C(n_697), .Y(n_688) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .Y(n_503) );
INVx1_ASAP7_75t_SL g551 ( .A(n_504), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_504), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g683 ( .A(n_504), .B(n_539), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_507), .B(n_553), .Y(n_675) );
AND2x2_ASAP7_75t_L g582 ( .A(n_508), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_SL g586 ( .A(n_509), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_509), .B(n_592), .Y(n_622) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_519), .Y(n_509) );
AND2x2_ASAP7_75t_L g547 ( .A(n_510), .B(n_520), .Y(n_547) );
INVx4_ASAP7_75t_L g559 ( .A(n_510), .Y(n_559) );
BUFx3_ASAP7_75t_L g602 ( .A(n_510), .Y(n_602) );
AND3x2_ASAP7_75t_L g617 ( .A(n_510), .B(n_618), .C(n_619), .Y(n_617) );
AND2x2_ASAP7_75t_L g699 ( .A(n_519), .B(n_613), .Y(n_699) );
AND2x2_ASAP7_75t_L g707 ( .A(n_519), .B(n_592), .Y(n_707) );
INVx1_ASAP7_75t_SL g712 ( .A(n_519), .Y(n_712) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_529), .Y(n_519) );
INVx1_ASAP7_75t_SL g570 ( .A(n_520), .Y(n_570) );
AND2x2_ASAP7_75t_L g593 ( .A(n_520), .B(n_559), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_520), .B(n_543), .Y(n_595) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_520), .Y(n_635) );
OR2x2_ASAP7_75t_L g640 ( .A(n_520), .B(n_559), .Y(n_640) );
INVx2_ASAP7_75t_L g545 ( .A(n_529), .Y(n_545) );
AND2x2_ASAP7_75t_L g580 ( .A(n_529), .B(n_560), .Y(n_580) );
OR2x2_ASAP7_75t_L g600 ( .A(n_529), .B(n_560), .Y(n_600) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_529), .Y(n_620) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g670 ( .A1(n_538), .A2(n_579), .B(n_671), .Y(n_670) );
AOI322xp5_ASAP7_75t_L g706 ( .A1(n_540), .A2(n_550), .A3(n_577), .B1(n_707), .B2(n_708), .C1(n_710), .C2(n_713), .Y(n_706) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_542), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_543), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g569 ( .A(n_544), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g637 ( .A(n_545), .B(n_559), .Y(n_637) );
AND2x2_ASAP7_75t_L g704 ( .A(n_545), .B(n_560), .Y(n_704) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g645 ( .A(n_547), .B(n_599), .Y(n_645) );
AOI31xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_552), .A3(n_555), .B(n_556), .Y(n_548) );
AND2x2_ASAP7_75t_L g604 ( .A(n_550), .B(n_582), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_550), .B(n_574), .Y(n_686) );
AND2x2_ASAP7_75t_L g705 ( .A(n_550), .B(n_610), .Y(n_705) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_553), .B(n_582), .Y(n_594) );
NAND2x1p5_ASAP7_75t_L g628 ( .A(n_553), .B(n_611), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_553), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_553), .B(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_554), .B(n_611), .Y(n_643) );
INVx1_ASAP7_75t_L g687 ( .A(n_554), .Y(n_687) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_569), .Y(n_557) );
INVxp67_ASAP7_75t_L g639 ( .A(n_558), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_559), .B(n_570), .Y(n_575) );
INVx1_ASAP7_75t_L g681 ( .A(n_559), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_559), .B(n_658), .Y(n_692) );
BUFx3_ASAP7_75t_L g592 ( .A(n_560), .Y(n_592) );
AND2x2_ASAP7_75t_L g618 ( .A(n_560), .B(n_570), .Y(n_618) );
INVx2_ASAP7_75t_L g658 ( .A(n_560), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_569), .B(n_691), .Y(n_690) );
AOI211xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_576), .B(n_578), .C(n_587), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AOI21xp33_ASAP7_75t_L g621 ( .A1(n_573), .A2(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_574), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_574), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g654 ( .A(n_575), .B(n_600), .Y(n_654) );
INVx3_ASAP7_75t_L g585 ( .A(n_577), .Y(n_585) );
OAI22xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_581), .B1(n_584), .B2(n_586), .Y(n_578) );
OAI21xp5_ASAP7_75t_SL g603 ( .A1(n_580), .A2(n_604), .B(n_605), .Y(n_603) );
AND2x2_ASAP7_75t_L g629 ( .A(n_580), .B(n_593), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_580), .B(n_681), .Y(n_680) );
INVxp67_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g584 ( .A(n_583), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g653 ( .A(n_583), .Y(n_653) );
OAI21xp5_ASAP7_75t_SL g597 ( .A1(n_584), .A2(n_598), .B(n_603), .Y(n_597) );
OAI22xp33_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_590), .B1(n_594), .B2(n_595), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_589), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g613 ( .A(n_592), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_592), .B(n_635), .Y(n_634) );
NOR3xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_608), .C(n_621), .Y(n_596) );
OAI22xp5_ASAP7_75t_SL g663 ( .A1(n_598), .A2(n_664), .B1(n_668), .B2(n_669), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_599), .B(n_601), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g668 ( .A(n_600), .B(n_601), .Y(n_668) );
AND2x2_ASAP7_75t_L g676 ( .A(n_601), .B(n_657), .Y(n_676) );
CKINVDCx16_ASAP7_75t_R g601 ( .A(n_602), .Y(n_601) );
O2A1O1Ixp33_ASAP7_75t_SL g684 ( .A1(n_602), .A2(n_685), .B(n_686), .C(n_687), .Y(n_684) );
OR2x2_ASAP7_75t_L g711 ( .A(n_602), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
OAI21xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_612), .B(n_614), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g646 ( .A1(n_610), .A2(n_647), .B(n_648), .C(n_651), .Y(n_646) );
OAI21xp33_ASAP7_75t_SL g614 ( .A1(n_615), .A2(n_616), .B(n_617), .Y(n_614) );
AND2x2_ASAP7_75t_L g679 ( .A(n_618), .B(n_637), .Y(n_679) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g657 ( .A(n_620), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g662 ( .A(n_622), .Y(n_662) );
NAND3xp33_ASAP7_75t_SL g625 ( .A(n_626), .B(n_646), .C(n_659), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B(n_630), .C(n_638), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g696 ( .A(n_633), .Y(n_696) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g656 ( .A(n_635), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_635), .B(n_704), .Y(n_703) );
INVxp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B(n_641), .C(n_642), .Y(n_638) );
INVx2_ASAP7_75t_SL g650 ( .A(n_640), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_641), .A2(n_652), .B1(n_654), .B2(n_655), .Y(n_651) );
OAI21xp33_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_644), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
AOI211xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_662), .B(n_663), .C(n_670), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVxp33_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g713 ( .A(n_667), .Y(n_713) );
NAND4xp25_ASAP7_75t_L g672 ( .A(n_673), .B(n_688), .C(n_701), .D(n_706), .Y(n_672) );
AOI211xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_676), .B(n_677), .C(n_684), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .B(n_682), .Y(n_677) );
AOI21xp33_ASAP7_75t_L g697 ( .A1(n_678), .A2(n_698), .B(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_685), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_705), .Y(n_701) );
INVxp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g729 ( .A(n_714), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_717), .Y(n_716) );
CKINVDCx16_ASAP7_75t_R g725 ( .A(n_719), .Y(n_725) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx3_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
endmodule