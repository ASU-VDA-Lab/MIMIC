module real_jpeg_23130_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_249;
wire n_83;
wire n_215;
wire n_166;
wire n_221;
wire n_292;
wire n_286;
wire n_288;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_197;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_200;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_258;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_1),
.A2(n_32),
.B1(n_61),
.B2(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_1),
.A2(n_32),
.B1(n_68),
.B2(n_69),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_1),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx8_ASAP7_75t_SL g67 ( 
.A(n_4),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_5),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_5),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_5),
.A2(n_60),
.B1(n_68),
.B2(n_69),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_60),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_60),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_6),
.A2(n_46),
.B1(n_68),
.B2(n_69),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_46),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_7),
.A2(n_62),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_7),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_7),
.A2(n_68),
.B1(n_69),
.B2(n_119),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_119),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_119),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_8),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_8),
.B(n_77),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_8),
.B(n_31),
.C(n_50),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_163),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_8),
.B(n_125),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_8),
.A2(n_93),
.B1(n_233),
.B2(n_236),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_10),
.A2(n_61),
.B1(n_73),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_10),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_10),
.A2(n_68),
.B1(n_69),
.B2(n_167),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_167),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_167),
.Y(n_233)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_55),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_12),
.A2(n_55),
.B1(n_68),
.B2(n_69),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_14),
.A2(n_35),
.B1(n_68),
.B2(n_69),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_14),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_14),
.A2(n_35),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_15),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_150),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_148),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_120),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_19),
.B(n_120),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_90),
.C(n_101),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_20),
.A2(n_21),
.B1(n_90),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_56),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_22),
.B(n_78),
.C(n_89),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_23),
.A2(n_24),
.B1(n_39),
.B2(n_40),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_25),
.A2(n_93),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_26),
.A2(n_36),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_27),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_29),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_29),
.A2(n_93),
.B(n_106),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_37),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_31),
.B1(n_50),
.B2(n_51),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_30),
.B(n_238),
.Y(n_237)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_33),
.A2(n_181),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_34),
.B(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_36),
.A2(n_105),
.B1(n_107),
.B2(n_180),
.Y(n_179)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_37),
.Y(n_236)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_38),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_38),
.B(n_163),
.Y(n_238)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_53),
.B2(n_54),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_42),
.A2(n_52),
.B(n_111),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_44),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_44),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_43),
.A2(n_82),
.B(n_247),
.C(n_249),
.Y(n_246)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_44),
.B(n_208),
.Y(n_207)
);

NOR3xp33_ASAP7_75t_L g249 ( 
.A(n_44),
.B(n_68),
.C(n_81),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_47),
.B(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_47),
.A2(n_98),
.B(n_129),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_47),
.A2(n_53),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_47),
.A2(n_53),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_48),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_48),
.A2(n_52),
.B1(n_212),
.B2(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_48),
.A2(n_128),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_52),
.B(n_163),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_53),
.B(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_54),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_78),
.B1(n_79),
.B2(n_89),
.Y(n_56)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_63),
.B(n_75),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_59),
.A2(n_64),
.B1(n_77),
.B2(n_117),
.Y(n_116)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_61),
.B(n_163),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_61),
.B(n_68),
.C(n_71),
.Y(n_183)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_63),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_63),
.A2(n_65),
.B1(n_166),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_64),
.A2(n_77),
.B1(n_162),
.B2(n_165),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_72),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_66),
.A2(n_69),
.B(n_164),
.C(n_183),
.Y(n_182)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_69),
.B1(n_81),
.B2(n_82),
.Y(n_86)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

HAxp5_ASAP7_75t_SL g248 ( 
.A(n_69),
.B(n_163),
.CON(n_248),
.SN(n_248)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_74),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_76),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_77),
.B(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B(n_84),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_80),
.A2(n_175),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_83),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_85),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_85),
.A2(n_125),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_85),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_85),
.A2(n_125),
.B1(n_198),
.B2(n_248),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_90),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_100),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_91),
.A2(n_92),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_95),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_104),
.B(n_106),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_93),
.A2(n_108),
.B1(n_226),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_101),
.B(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_113),
.C(n_116),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_102),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_110),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_110),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_113),
.B(n_116),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_114),
.B(n_125),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_117),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_120)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_131),
.B1(n_143),
.B2(n_144),
.Y(n_121)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_127),
.B(n_130),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_127),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_142),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_145),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_289),
.B(n_294),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_200),
.B(n_280),
.C(n_288),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_185),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_153),
.B(n_185),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_168),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_155),
.B(n_156),
.C(n_168),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.C(n_161),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_160),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_187),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_177),
.B2(n_184),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_171),
.B(n_173),
.C(n_184),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B(n_176),
.Y(n_173)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_179),
.B1(n_182),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_182),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.C(n_190),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_186),
.B(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_188),
.B(n_190),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.C(n_196),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_191),
.A2(n_194),
.B1(n_195),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_191),
.Y(n_265)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_196),
.B(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_279),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_274),
.B(n_278),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_259),
.B(n_273),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_242),
.B(n_258),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_222),
.B(n_241),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_213),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_213),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_209),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_217),
.C(n_220),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_215),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_221),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_229),
.B(n_240),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_228),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_234),
.B(n_239),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_232),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_257),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_257),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_252),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_253),
.C(n_254),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_250),
.B2(n_251),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_251),
.Y(n_268)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_256),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_261),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_266),
.B2(n_267),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_269),
.C(n_271),
.Y(n_277)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_269),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_277),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_285),
.C(n_287),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);


endmodule