module fake_netlist_6_2985_n_1780 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1780);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1780;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_11),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_46),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_138),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_16),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_82),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_41),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_4),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_87),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_40),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_74),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_9),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_17),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_39),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_68),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_16),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_18),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_79),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_71),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_129),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_14),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_8),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_35),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_113),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_107),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_26),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_34),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_61),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_157),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_76),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_38),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_86),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_53),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_150),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_125),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_54),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_112),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_88),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_127),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_110),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_141),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_52),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_152),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_42),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_80),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_13),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_70),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_17),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_156),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_2),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_111),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_4),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_134),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_42),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_62),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_7),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_149),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_97),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_154),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_13),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_2),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_105),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_90),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_35),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_14),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_143),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_15),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_57),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_5),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_7),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_99),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_58),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_46),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_26),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_48),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_44),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_135),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_72),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_6),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_159),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_48),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_19),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_75),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_54),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_148),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_83),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_12),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_78),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_43),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_158),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_155),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_92),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_18),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_6),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_20),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_38),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g267 ( 
.A(n_63),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_60),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_102),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_50),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_77),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_118),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_109),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_47),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_22),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_162),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_9),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_44),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_30),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_11),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_49),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_93),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_23),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_15),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_100),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_123),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_57),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_98),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_3),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_29),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_115),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_8),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_94),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_5),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_116),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_65),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_85),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_126),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_73),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_101),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_104),
.Y(n_301)
);

BUFx8_ASAP7_75t_SL g302 ( 
.A(n_103),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_69),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_30),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_37),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_120),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_32),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_52),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_50),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_39),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_132),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_53),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_19),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_24),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_106),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_49),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_95),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_55),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_25),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_1),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_32),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g322 ( 
.A(n_59),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_1),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_165),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_192),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_302),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_165),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_166),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_322),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_322),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_184),
.B(n_160),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_200),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_173),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_322),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_181),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_203),
.Y(n_337)
);

NAND2xp33_ASAP7_75t_R g338 ( 
.A(n_277),
.B(n_0),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_322),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_322),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_322),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_297),
.B(n_0),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_190),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_231),
.B(n_3),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_190),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_186),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_280),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_268),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_271),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_272),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_295),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_214),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_187),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_280),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_174),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_310),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_174),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_182),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_182),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_252),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_283),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_193),
.Y(n_363)
);

INVxp33_ASAP7_75t_SL g364 ( 
.A(n_171),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_184),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_197),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_207),
.B(n_10),
.Y(n_367)
);

BUFx6f_ASAP7_75t_SL g368 ( 
.A(n_273),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_263),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_185),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_202),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_170),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_206),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_185),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_212),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_213),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_221),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_170),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_212),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_223),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_237),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_237),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_225),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_L g384 ( 
.A(n_224),
.B(n_12),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_176),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_164),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_240),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_240),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_227),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_242),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_222),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_164),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_242),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_283),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_207),
.B(n_20),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_243),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_228),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_361),
.Y(n_398)
);

OA21x2_ASAP7_75t_L g399 ( 
.A1(n_325),
.A2(n_249),
.B(n_243),
.Y(n_399)
);

NAND2xp33_ASAP7_75t_L g400 ( 
.A(n_332),
.B(n_188),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_372),
.B(n_222),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_325),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_348),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_330),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_369),
.B(n_283),
.Y(n_406)
);

OR2x6_ASAP7_75t_L g407 ( 
.A(n_332),
.B(n_241),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_330),
.Y(n_408)
);

BUFx8_ASAP7_75t_L g409 ( 
.A(n_368),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_356),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_331),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_332),
.B(n_241),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_363),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_378),
.B(n_168),
.Y(n_414)
);

AND2x2_ASAP7_75t_SL g415 ( 
.A(n_332),
.B(n_172),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_335),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_335),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_386),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_365),
.B(n_168),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_391),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_339),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_339),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_340),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_371),
.Y(n_426)
);

INVx6_ASAP7_75t_L g427 ( 
.A(n_340),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_391),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_341),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_324),
.A2(n_199),
.B1(n_321),
.B2(n_320),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_356),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_341),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_342),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_367),
.B(n_232),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_342),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_358),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_392),
.B(n_172),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_358),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_392),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_344),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_359),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_328),
.A2(n_163),
.B1(n_167),
.B2(n_308),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_359),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_344),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_346),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_346),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_329),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_355),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_360),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_360),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_355),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_395),
.B(n_196),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_370),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_370),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_373),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_374),
.Y(n_456)
);

OA21x2_ASAP7_75t_L g457 ( 
.A1(n_374),
.A2(n_251),
.B(n_249),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_375),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_375),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_379),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_379),
.B(n_169),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_381),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_381),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_382),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_382),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_326),
.Y(n_466)
);

NOR2x1_ASAP7_75t_L g467 ( 
.A(n_376),
.B(n_175),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_387),
.B(n_233),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_387),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_388),
.B(n_169),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_338),
.A2(n_266),
.B1(n_234),
.B2(n_265),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_415),
.B(n_452),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_405),
.Y(n_473)
);

NOR2x1p5_ASAP7_75t_L g474 ( 
.A(n_447),
.B(n_327),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_408),
.Y(n_475)
);

OAI22xp33_ASAP7_75t_L g476 ( 
.A1(n_406),
.A2(n_357),
.B1(n_284),
.B2(n_369),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_399),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_408),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_417),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_417),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_452),
.B(n_343),
.C(n_385),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_417),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_421),
.B(n_388),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_399),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_405),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_415),
.B(n_334),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_SL g487 ( 
.A1(n_406),
.A2(n_368),
.B1(n_353),
.B2(n_352),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_408),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_408),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_405),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_415),
.A2(n_384),
.B1(n_251),
.B2(n_257),
.Y(n_491)
);

OAI22xp33_ASAP7_75t_L g492 ( 
.A1(n_422),
.A2(n_345),
.B1(n_189),
.B2(n_180),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_419),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_412),
.B(n_177),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_423),
.Y(n_495)
);

INVxp33_ASAP7_75t_L g496 ( 
.A(n_430),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_419),
.Y(n_497)
);

INVx5_ASAP7_75t_L g498 ( 
.A(n_405),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_413),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_423),
.Y(n_500)
);

BUFx4f_ASAP7_75t_L g501 ( 
.A(n_399),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_423),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_434),
.B(n_336),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_467),
.A2(n_380),
.B1(n_389),
.B2(n_383),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_447),
.B(n_347),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_412),
.B(n_177),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_421),
.B(n_390),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_405),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_424),
.Y(n_509)
);

OR2x6_ASAP7_75t_L g510 ( 
.A(n_467),
.B(n_257),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_413),
.Y(n_511)
);

AND2x6_ASAP7_75t_L g512 ( 
.A(n_412),
.B(n_175),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_447),
.B(n_364),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_419),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_419),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_412),
.A2(n_270),
.B1(n_274),
.B2(n_275),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_421),
.B(n_390),
.Y(n_517)
);

AND3x2_ASAP7_75t_L g518 ( 
.A(n_412),
.B(n_296),
.C(n_247),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_429),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_405),
.Y(n_520)
);

AND3x2_ASAP7_75t_L g521 ( 
.A(n_428),
.B(n_296),
.C(n_247),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_424),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_428),
.B(n_362),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_414),
.B(n_393),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_461),
.B(n_178),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_414),
.B(n_354),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_426),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_429),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_429),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_401),
.B(n_393),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_399),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_447),
.B(n_366),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_424),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_405),
.Y(n_534)
);

OR2x6_ASAP7_75t_L g535 ( 
.A(n_447),
.B(n_270),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_422),
.B(n_377),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_399),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_399),
.Y(n_538)
);

BUFx10_ASAP7_75t_L g539 ( 
.A(n_426),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_455),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_429),
.Y(n_541)
);

BUFx4f_ASAP7_75t_L g542 ( 
.A(n_457),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_405),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_409),
.B(n_397),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_428),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_411),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_425),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_457),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_409),
.B(n_394),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_432),
.Y(n_550)
);

INVx4_ASAP7_75t_L g551 ( 
.A(n_411),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_401),
.B(n_274),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_425),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_468),
.B(n_396),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_468),
.B(n_396),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_407),
.B(n_248),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_402),
.Y(n_557)
);

BUFx10_ASAP7_75t_L g558 ( 
.A(n_455),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_402),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_402),
.Y(n_560)
);

INVxp33_ASAP7_75t_L g561 ( 
.A(n_430),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_407),
.B(n_402),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_466),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_402),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_409),
.B(n_273),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_432),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_R g567 ( 
.A(n_401),
.B(n_179),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_411),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_466),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_407),
.A2(n_275),
.B1(n_319),
.B2(n_278),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_409),
.B(n_273),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_411),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_432),
.Y(n_573)
);

INVxp67_ASAP7_75t_SL g574 ( 
.A(n_418),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_432),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_433),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_411),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_418),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_398),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_L g580 ( 
.A(n_411),
.B(n_188),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_407),
.B(n_253),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_411),
.Y(n_582)
);

INVx5_ASAP7_75t_L g583 ( 
.A(n_411),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_398),
.B(n_368),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_418),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_433),
.Y(n_586)
);

NAND3xp33_ASAP7_75t_L g587 ( 
.A(n_471),
.B(n_246),
.C(n_323),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_433),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_418),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_409),
.B(n_286),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_418),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_416),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_435),
.Y(n_593)
);

XNOR2x2_ASAP7_75t_L g594 ( 
.A(n_471),
.B(n_278),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_SL g595 ( 
.A(n_409),
.B(n_333),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_435),
.Y(n_596)
);

BUFx4f_ASAP7_75t_L g597 ( 
.A(n_457),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_407),
.B(n_351),
.Y(n_598)
);

NAND2xp33_ASAP7_75t_SL g599 ( 
.A(n_461),
.B(n_191),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_435),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_407),
.A2(n_350),
.B1(n_349),
.B2(n_337),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_433),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_435),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_407),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_461),
.B(n_470),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_427),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_427),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_458),
.B(n_459),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_457),
.Y(n_609)
);

AND2x6_ASAP7_75t_L g610 ( 
.A(n_470),
.B(n_178),
.Y(n_610)
);

AO22x2_ASAP7_75t_L g611 ( 
.A1(n_442),
.A2(n_319),
.B1(n_281),
.B2(n_289),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_427),
.Y(n_612)
);

BUFx10_ASAP7_75t_L g613 ( 
.A(n_437),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_453),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_400),
.A2(n_281),
.B1(n_289),
.B2(n_294),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_435),
.B(n_255),
.Y(n_616)
);

INVxp33_ASAP7_75t_L g617 ( 
.A(n_442),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_457),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_472),
.B(n_400),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_499),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_605),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_605),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_548),
.A2(n_457),
.B1(n_470),
.B2(n_305),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_548),
.A2(n_609),
.B1(n_618),
.B2(n_484),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_605),
.B(n_458),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_503),
.B(n_458),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_479),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_530),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_526),
.B(n_194),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_530),
.B(n_410),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_545),
.Y(n_631)
);

BUFx5_ASAP7_75t_L g632 ( 
.A(n_477),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_491),
.B(n_416),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_609),
.A2(n_618),
.B1(n_484),
.B2(n_531),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_542),
.B(n_188),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_486),
.A2(n_267),
.B1(n_256),
.B2(n_258),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_542),
.B(n_597),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_542),
.B(n_188),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_545),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_477),
.A2(n_309),
.B1(n_305),
.B2(n_294),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_554),
.B(n_416),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_613),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_531),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_579),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_510),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_579),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_L g647 ( 
.A(n_512),
.B(n_276),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_R g648 ( 
.A(n_499),
.B(n_288),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_554),
.B(n_416),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_555),
.B(n_416),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_479),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_563),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_537),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_537),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_538),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_567),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_555),
.B(n_420),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_595),
.B(n_286),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_597),
.B(n_188),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_480),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_563),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_538),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_481),
.B(n_195),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_480),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_597),
.A2(n_437),
.B(n_198),
.Y(n_665)
);

BUFx8_ASAP7_75t_L g666 ( 
.A(n_523),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_536),
.B(n_201),
.Y(n_667)
);

A2O1A1Ixp33_ASAP7_75t_L g668 ( 
.A1(n_501),
.A2(n_309),
.B(n_459),
.C(n_204),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_482),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_510),
.A2(n_291),
.B1(n_293),
.B2(n_298),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_482),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_513),
.B(n_205),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_523),
.B(n_216),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_584),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_475),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_495),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_552),
.B(n_431),
.Y(n_677)
);

AO221x1_ASAP7_75t_L g678 ( 
.A1(n_611),
.A2(n_183),
.B1(n_198),
.B2(n_217),
.C(n_219),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_475),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_495),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_SL g681 ( 
.A(n_569),
.B(n_286),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_483),
.B(n_436),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_613),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_507),
.B(n_420),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_507),
.B(n_420),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_587),
.B(n_218),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_535),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_510),
.A2(n_306),
.B1(n_299),
.B2(n_300),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_478),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_501),
.B(n_437),
.Y(n_690)
);

BUFx12f_ASAP7_75t_L g691 ( 
.A(n_511),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_510),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_501),
.B(n_437),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_599),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_562),
.B(n_437),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_610),
.A2(n_183),
.B1(n_204),
.B2(n_211),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_500),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_525),
.B(n_436),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_511),
.Y(n_699)
);

BUFx12f_ASAP7_75t_SL g700 ( 
.A(n_552),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_511),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_604),
.A2(n_236),
.B1(n_311),
.B2(n_285),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_500),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_604),
.B(n_437),
.Y(n_704)
);

AND2x4_ASAP7_75t_SL g705 ( 
.A(n_527),
.B(n_317),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_517),
.B(n_427),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_532),
.B(n_220),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_535),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_502),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_517),
.B(n_438),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_502),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_524),
.B(n_427),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_527),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_524),
.B(n_427),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_509),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_552),
.B(n_226),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_574),
.B(n_578),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_608),
.B(n_427),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_599),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_613),
.B(n_453),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_535),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_610),
.A2(n_598),
.B1(n_552),
.B2(n_581),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_509),
.B(n_453),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_478),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_522),
.B(n_453),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_522),
.B(n_453),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_496),
.B(n_438),
.Y(n_727)
);

INVxp67_ASAP7_75t_SL g728 ( 
.A(n_473),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_533),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_492),
.B(n_230),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_547),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_488),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_547),
.B(n_453),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_553),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_553),
.B(n_453),
.Y(n_735)
);

BUFx8_ASAP7_75t_L g736 ( 
.A(n_594),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_557),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_594),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_504),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_610),
.A2(n_301),
.B1(n_303),
.B2(n_210),
.Y(n_740)
);

INVxp67_ASAP7_75t_SL g741 ( 
.A(n_473),
.Y(n_741)
);

NOR2xp67_ASAP7_75t_L g742 ( 
.A(n_601),
.B(n_544),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_557),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_559),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_592),
.B(n_453),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_592),
.B(n_445),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_559),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_494),
.B(n_506),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_488),
.Y(n_749)
);

NOR3xp33_ASAP7_75t_L g750 ( 
.A(n_476),
.B(n_290),
.C(n_279),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_L g751 ( 
.A(n_505),
.B(n_441),
.Y(n_751)
);

BUFx5_ASAP7_75t_L g752 ( 
.A(n_560),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_561),
.A2(n_459),
.B(n_315),
.C(n_311),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_535),
.B(n_235),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_494),
.B(n_208),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_560),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_564),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_489),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_489),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_525),
.B(n_454),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_525),
.B(n_454),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_617),
.B(n_238),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_585),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_585),
.B(n_454),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_589),
.B(n_209),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_589),
.B(n_440),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_591),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_593),
.B(n_454),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_527),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_556),
.A2(n_211),
.B1(n_315),
.B2(n_285),
.Y(n_770)
);

BUFx4f_ASAP7_75t_L g771 ( 
.A(n_610),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_596),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_565),
.B(n_239),
.Y(n_773)
);

NOR2x1p5_ASAP7_75t_L g774 ( 
.A(n_487),
.B(n_244),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_516),
.B(n_259),
.C(n_264),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_521),
.B(n_518),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_596),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_L g778 ( 
.A(n_512),
.B(n_215),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_665),
.A2(n_534),
.B(n_490),
.Y(n_779)
);

O2A1O1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_753),
.A2(n_738),
.B(n_668),
.C(n_719),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_634),
.A2(n_570),
.B1(n_615),
.B2(n_549),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_619),
.A2(n_534),
.B(n_490),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_657),
.B(n_610),
.Y(n_783)
);

AOI21x1_ASAP7_75t_L g784 ( 
.A1(n_635),
.A2(n_616),
.B(n_603),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_703),
.Y(n_785)
);

AOI21x1_ASAP7_75t_L g786 ( 
.A1(n_635),
.A2(n_603),
.B(n_600),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_628),
.B(n_539),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_707),
.B(n_610),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_690),
.A2(n_534),
.B(n_490),
.Y(n_789)
);

AOI21x1_ASAP7_75t_L g790 ( 
.A1(n_638),
.A2(n_600),
.B(n_614),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_690),
.A2(n_577),
.B(n_551),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_638),
.A2(n_519),
.B(n_493),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_727),
.Y(n_793)
);

NOR2x1_ASAP7_75t_L g794 ( 
.A(n_742),
.B(n_474),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_628),
.B(n_539),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_L g796 ( 
.A(n_667),
.B(n_571),
.C(n_590),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_762),
.B(n_539),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_656),
.B(n_762),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_703),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_693),
.A2(n_551),
.B(n_577),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_672),
.A2(n_229),
.B(n_219),
.C(n_217),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_707),
.B(n_512),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_641),
.B(n_512),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_649),
.B(n_512),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_693),
.A2(n_551),
.B(n_577),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_637),
.A2(n_543),
.B(n_546),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_644),
.B(n_540),
.Y(n_807)
);

AOI21x1_ASAP7_75t_L g808 ( 
.A1(n_659),
.A2(n_614),
.B(n_493),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_650),
.B(n_508),
.Y(n_809)
);

O2A1O1Ixp33_ASAP7_75t_SL g810 ( 
.A1(n_668),
.A2(n_659),
.B(n_753),
.C(n_626),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_653),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_637),
.A2(n_546),
.B(n_543),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_672),
.A2(n_215),
.B(n_229),
.C(n_236),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_745),
.A2(n_546),
.B(n_543),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_711),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_667),
.B(n_508),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_663),
.A2(n_250),
.B(n_269),
.C(n_282),
.Y(n_817)
);

NAND2x1p5_ASAP7_75t_L g818 ( 
.A(n_653),
.B(n_606),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_632),
.B(n_540),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_745),
.A2(n_720),
.B(n_746),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_621),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_682),
.B(n_710),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_630),
.B(n_508),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_629),
.B(n_520),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_646),
.B(n_540),
.Y(n_825)
);

AOI21xp33_ASAP7_75t_L g826 ( 
.A1(n_663),
.A2(n_611),
.B(n_250),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_739),
.B(n_558),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_711),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_694),
.B(n_558),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_629),
.B(n_558),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_625),
.A2(n_514),
.B(n_497),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_653),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_643),
.B(n_520),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_720),
.A2(n_572),
.B(n_473),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_701),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_SL g836 ( 
.A(n_620),
.B(n_317),
.Y(n_836)
);

NAND2x1_ASAP7_75t_L g837 ( 
.A(n_653),
.B(n_520),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_632),
.B(n_473),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_623),
.B(n_568),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_623),
.B(n_568),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_773),
.A2(n_686),
.B(n_622),
.C(n_730),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_684),
.B(n_685),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_718),
.A2(n_485),
.B(n_572),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_748),
.A2(n_485),
.B(n_572),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_706),
.A2(n_485),
.B(n_572),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_712),
.A2(n_485),
.B(n_582),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_714),
.A2(n_485),
.B(n_582),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_652),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_715),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_654),
.B(n_582),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_673),
.B(n_611),
.Y(n_851)
);

BUFx4f_ASAP7_75t_L g852 ( 
.A(n_691),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_674),
.B(n_673),
.Y(n_853)
);

AOI21x1_ASAP7_75t_L g854 ( 
.A1(n_766),
.A2(n_519),
.B(n_497),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_631),
.B(n_514),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_640),
.A2(n_611),
.B1(n_282),
.B2(n_269),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_715),
.Y(n_857)
);

O2A1O1Ixp33_ASAP7_75t_L g858 ( 
.A1(n_702),
.A2(n_580),
.B(n_528),
.C(n_529),
.Y(n_858)
);

AOI21x1_ASAP7_75t_L g859 ( 
.A1(n_766),
.A2(n_573),
.B(n_515),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_654),
.A2(n_576),
.B(n_529),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_655),
.B(n_515),
.Y(n_861)
);

AOI21x1_ASAP7_75t_L g862 ( 
.A1(n_695),
.A2(n_541),
.B(n_566),
.Y(n_862)
);

OAI22xp33_ASAP7_75t_L g863 ( 
.A1(n_658),
.A2(n_449),
.B1(n_441),
.B2(n_443),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_695),
.A2(n_761),
.B(n_760),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_737),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_773),
.A2(n_586),
.B(n_573),
.C(n_575),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_743),
.Y(n_867)
);

AO22x1_ASAP7_75t_L g868 ( 
.A1(n_736),
.A2(n_245),
.B1(n_254),
.B2(n_287),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_662),
.A2(n_633),
.B(n_634),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_704),
.A2(n_583),
.B(n_498),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_722),
.A2(n_612),
.B1(n_607),
.B2(n_606),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_639),
.B(n_550),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_624),
.B(n_550),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_677),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_698),
.B(n_576),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_728),
.A2(n_583),
.B(n_498),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_661),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_627),
.B(n_588),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_744),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_686),
.A2(n_602),
.B(n_588),
.C(n_606),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_632),
.B(n_317),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_771),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_776),
.B(n_443),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_640),
.A2(n_602),
.B1(n_612),
.B2(n_607),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_771),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_730),
.A2(n_612),
.B(n_607),
.C(n_449),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_692),
.B(n_292),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_651),
.B(n_456),
.Y(n_888)
);

BUFx2_ASAP7_75t_L g889 ( 
.A(n_700),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_747),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_741),
.A2(n_439),
.B(n_465),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_716),
.B(n_304),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_756),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_660),
.B(n_456),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_664),
.B(n_456),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_632),
.B(n_450),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_666),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_754),
.A2(n_716),
.B(n_751),
.C(n_721),
.Y(n_898)
);

O2A1O1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_770),
.A2(n_464),
.B(n_463),
.C(n_462),
.Y(n_899)
);

O2A1O1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_765),
.A2(n_464),
.B(n_463),
.C(n_462),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_708),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_669),
.B(n_469),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_636),
.A2(n_469),
.B1(n_456),
.B2(n_460),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_754),
.B(n_687),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_632),
.A2(n_460),
.B1(n_450),
.B2(n_439),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_671),
.B(n_403),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_642),
.A2(n_448),
.B(n_403),
.Y(n_907)
);

AOI21x1_ASAP7_75t_L g908 ( 
.A1(n_723),
.A2(n_404),
.B(n_448),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_676),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_642),
.A2(n_448),
.B(n_404),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_681),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_680),
.B(n_307),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_666),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_683),
.A2(n_446),
.B(n_444),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_757),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_697),
.B(n_444),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_709),
.B(n_312),
.Y(n_917)
);

AO21x1_ASAP7_75t_L g918 ( 
.A1(n_765),
.A2(n_444),
.B(n_22),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_729),
.B(n_451),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_705),
.B(n_318),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_717),
.A2(n_451),
.B(n_440),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_763),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_767),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_778),
.A2(n_451),
.B(n_440),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_647),
.A2(n_451),
.B(n_440),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_750),
.B(n_313),
.Y(n_926)
);

NAND2x1p5_ASAP7_75t_L g927 ( 
.A(n_731),
.B(n_451),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_734),
.B(n_451),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_772),
.Y(n_929)
);

OAI21xp33_ASAP7_75t_L g930 ( 
.A1(n_648),
.A2(n_316),
.B(n_314),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_777),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_752),
.B(n_451),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_755),
.A2(n_440),
.B(n_23),
.C(n_24),
.Y(n_933)
);

O2A1O1Ixp5_ASAP7_75t_L g934 ( 
.A1(n_755),
.A2(n_440),
.B(n_66),
.C(n_67),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_696),
.A2(n_440),
.B(n_25),
.C(n_27),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_699),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_675),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_764),
.A2(n_21),
.B(n_27),
.C(n_28),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_679),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_752),
.B(n_440),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_689),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_725),
.A2(n_81),
.B(n_151),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_726),
.A2(n_64),
.B(n_145),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_752),
.B(n_153),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_733),
.A2(n_735),
.B(n_768),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_R g946 ( 
.A(n_713),
.B(n_140),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_645),
.B(n_139),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_670),
.B(n_21),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_696),
.A2(n_136),
.B1(n_133),
.B2(n_131),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_705),
.B(n_28),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_724),
.A2(n_128),
.B(n_124),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_732),
.A2(n_122),
.B(n_121),
.Y(n_952)
);

INVx4_ASAP7_75t_L g953 ( 
.A(n_752),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_SL g954 ( 
.A1(n_848),
.A2(n_835),
.B1(n_830),
.B2(n_911),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_883),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_877),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_798),
.B(n_793),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_953),
.A2(n_749),
.B(n_759),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_953),
.A2(n_779),
.B(n_842),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_864),
.A2(n_758),
.B(n_740),
.Y(n_960)
);

OAI21xp33_ASAP7_75t_SL g961 ( 
.A1(n_869),
.A2(n_678),
.B(n_688),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_856),
.A2(n_774),
.B1(n_775),
.B2(n_769),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_798),
.A2(n_736),
.B1(n_776),
.B2(n_752),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_811),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_803),
.A2(n_752),
.B(n_114),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_856),
.A2(n_648),
.B1(n_31),
.B2(n_33),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_804),
.A2(n_119),
.B(n_117),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_797),
.B(n_108),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_841),
.A2(n_29),
.B(n_31),
.C(n_33),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_802),
.A2(n_91),
.B(n_84),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_853),
.B(n_34),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_826),
.A2(n_36),
.B(n_37),
.C(n_40),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_882),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_892),
.A2(n_36),
.B1(n_41),
.B2(n_43),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_948),
.A2(n_45),
.B1(n_47),
.B2(n_51),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_811),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_892),
.A2(n_45),
.B(n_51),
.C(n_55),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_887),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_788),
.A2(n_56),
.B(n_58),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_874),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_853),
.A2(n_56),
.B(n_59),
.C(n_948),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_854),
.A2(n_859),
.B(n_862),
.Y(n_982)
);

AOI21x1_ASAP7_75t_L g983 ( 
.A1(n_808),
.A2(n_790),
.B(n_786),
.Y(n_983)
);

BUFx8_ASAP7_75t_L g984 ( 
.A(n_889),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_822),
.B(n_793),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_830),
.B(n_827),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_780),
.A2(n_945),
.B(n_783),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_909),
.B(n_851),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_827),
.B(n_904),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_SL g990 ( 
.A(n_852),
.B(n_936),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_785),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_796),
.A2(n_904),
.B(n_898),
.C(n_781),
.Y(n_992)
);

OAI22x1_ASAP7_75t_L g993 ( 
.A1(n_911),
.A2(n_874),
.B1(n_829),
.B2(n_807),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_817),
.A2(n_813),
.B(n_801),
.C(n_863),
.Y(n_994)
);

AND2x6_ASAP7_75t_L g995 ( 
.A(n_882),
.B(n_885),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_R g996 ( 
.A(n_829),
.B(n_807),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_883),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_824),
.A2(n_809),
.B(n_816),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_855),
.B(n_872),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_815),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_794),
.B(n_901),
.Y(n_1001)
);

O2A1O1Ixp5_ASAP7_75t_L g1002 ( 
.A1(n_881),
.A2(n_947),
.B(n_886),
.C(n_820),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_887),
.B(n_912),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_901),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_855),
.B(n_872),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_857),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_882),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_789),
.A2(n_800),
.B(n_805),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_917),
.A2(n_923),
.B(n_929),
.C(n_893),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_825),
.B(n_930),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_863),
.B(n_825),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_926),
.B(n_821),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_791),
.A2(n_782),
.B(n_838),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_810),
.A2(n_873),
.B(n_806),
.Y(n_1014)
);

NOR3xp33_ASAP7_75t_SL g1015 ( 
.A(n_787),
.B(n_795),
.C(n_933),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_843),
.A2(n_812),
.B(n_846),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_857),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_865),
.B(n_867),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_901),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_897),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_879),
.B(n_890),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_915),
.B(n_922),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_814),
.A2(n_932),
.B(n_940),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_SL g1024 ( 
.A1(n_913),
.A2(n_901),
.B1(n_949),
.B2(n_821),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_931),
.B(n_882),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_950),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_885),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_823),
.B(n_799),
.Y(n_1028)
);

INVxp67_ASAP7_75t_L g1029 ( 
.A(n_920),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_836),
.B(n_868),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_839),
.A2(n_840),
.B(n_833),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_946),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_935),
.A2(n_885),
.B1(n_828),
.B2(n_849),
.Y(n_1033)
);

OAI21xp33_ASAP7_75t_L g1034 ( 
.A1(n_946),
.A2(n_875),
.B(n_906),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_941),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_916),
.B(n_832),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_R g1037 ( 
.A(n_852),
.B(n_832),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_939),
.B(n_918),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_885),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_888),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_937),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_878),
.B(n_902),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_894),
.B(n_895),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_880),
.A2(n_866),
.B(n_831),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_847),
.A2(n_845),
.B(n_860),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_937),
.B(n_819),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_938),
.A2(n_899),
.B(n_900),
.C(n_944),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_905),
.A2(n_952),
.B1(n_944),
.B2(n_871),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_861),
.B(n_850),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_937),
.A2(n_896),
.B1(n_903),
.B2(n_884),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_919),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_844),
.A2(n_834),
.B(n_837),
.Y(n_1052)
);

AOI21x1_ASAP7_75t_L g1053 ( 
.A1(n_784),
.A2(n_908),
.B(n_928),
.Y(n_1053)
);

BUFx4f_ASAP7_75t_SL g1054 ( 
.A(n_937),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_818),
.Y(n_1055)
);

NOR2x1_ASAP7_75t_L g1056 ( 
.A(n_914),
.B(n_943),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_927),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_927),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_792),
.B(n_907),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_818),
.A2(n_925),
.B(n_921),
.Y(n_1060)
);

O2A1O1Ixp5_ASAP7_75t_L g1061 ( 
.A1(n_934),
.A2(n_910),
.B(n_891),
.C(n_942),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_858),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_951),
.A2(n_870),
.B1(n_924),
.B2(n_876),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_953),
.A2(n_665),
.B(n_637),
.Y(n_1064)
);

NOR3xp33_ASAP7_75t_SL g1065 ( 
.A(n_948),
.B(n_661),
.C(n_652),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_909),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_856),
.A2(n_634),
.B1(n_624),
.B2(n_623),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_953),
.A2(n_665),
.B(n_637),
.Y(n_1068)
);

OR2x6_ASAP7_75t_L g1069 ( 
.A(n_877),
.B(n_889),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_848),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_953),
.A2(n_665),
.B(n_637),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_883),
.B(n_628),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_841),
.A2(n_826),
.B(n_892),
.C(n_853),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_841),
.A2(n_826),
.B(n_892),
.C(n_853),
.Y(n_1074)
);

INVx2_ASAP7_75t_SL g1075 ( 
.A(n_883),
.Y(n_1075)
);

NAND3xp33_ASAP7_75t_SL g1076 ( 
.A(n_892),
.B(n_499),
.C(n_652),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_841),
.A2(n_892),
.B(n_798),
.C(n_667),
.Y(n_1077)
);

BUFx12f_ASAP7_75t_L g1078 ( 
.A(n_889),
.Y(n_1078)
);

NAND2x1p5_ASAP7_75t_L g1079 ( 
.A(n_882),
.B(n_653),
.Y(n_1079)
);

HB1xp67_ASAP7_75t_L g1080 ( 
.A(n_874),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_856),
.A2(n_634),
.B1(n_624),
.B2(n_623),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_848),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_793),
.B(n_634),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_798),
.B(n_853),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_953),
.A2(n_665),
.B(n_637),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_901),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_811),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_SL g1088 ( 
.A1(n_848),
.A2(n_661),
.B1(n_652),
.B2(n_561),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_848),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_848),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_793),
.B(n_634),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_841),
.A2(n_892),
.B(n_798),
.C(n_667),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_909),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_798),
.B(n_853),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_811),
.Y(n_1095)
);

NAND2xp33_ASAP7_75t_R g1096 ( 
.A(n_797),
.B(n_652),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_854),
.A2(n_859),
.B(n_862),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_798),
.B(n_853),
.Y(n_1098)
);

NAND3xp33_ASAP7_75t_SL g1099 ( 
.A(n_892),
.B(n_499),
.C(n_652),
.Y(n_1099)
);

OR2x6_ASAP7_75t_SL g1100 ( 
.A(n_796),
.B(n_413),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_798),
.B(n_853),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_856),
.A2(n_634),
.B1(n_624),
.B2(n_623),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1003),
.B(n_1084),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_991),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_992),
.A2(n_1077),
.A3(n_1092),
.B(n_1048),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1018),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1094),
.A2(n_966),
.B1(n_1012),
.B2(n_971),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_SL g1108 ( 
.A(n_1067),
.B(n_1081),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_959),
.A2(n_998),
.B(n_1064),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_1069),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1010),
.A2(n_994),
.B(n_961),
.C(n_1047),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1000),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1021),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1068),
.A2(n_1085),
.B(n_1071),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_1078),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_966),
.A2(n_978),
.B1(n_1101),
.B2(n_1098),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_985),
.B(n_988),
.Y(n_1117)
);

AOI221x1_ASAP7_75t_L g1118 ( 
.A1(n_969),
.A2(n_993),
.B1(n_979),
.B2(n_1048),
.C(n_1014),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_987),
.A2(n_1008),
.B(n_1060),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1001),
.B(n_1072),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1022),
.Y(n_1121)
);

INVxp67_ASAP7_75t_SL g1122 ( 
.A(n_1067),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_987),
.A2(n_1031),
.B(n_1002),
.Y(n_1123)
);

AO21x1_ASAP7_75t_L g1124 ( 
.A1(n_986),
.A2(n_1102),
.B(n_1081),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1013),
.A2(n_1023),
.B(n_960),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_957),
.B(n_989),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_1001),
.B(n_1072),
.Y(n_1127)
);

OAI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1096),
.A2(n_1102),
.B1(n_963),
.B2(n_990),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_980),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_981),
.A2(n_1009),
.B(n_1034),
.C(n_1015),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_955),
.B(n_1075),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_995),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1052),
.A2(n_1016),
.B(n_1045),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_SL g1134 ( 
.A1(n_1079),
.A2(n_1042),
.B(n_968),
.Y(n_1134)
);

BUFx2_ASAP7_75t_R g1135 ( 
.A(n_1070),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1061),
.A2(n_1044),
.B(n_965),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_960),
.A2(n_1044),
.B(n_1042),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1066),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1076),
.B(n_1099),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_SL g1140 ( 
.A1(n_1025),
.A2(n_1091),
.B(n_1083),
.C(n_999),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_975),
.A2(n_974),
.B1(n_1024),
.B2(n_962),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_SL g1142 ( 
.A1(n_1079),
.A2(n_1043),
.B(n_1005),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1093),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1083),
.B(n_1091),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1062),
.A2(n_1043),
.B(n_1059),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1019),
.B(n_1026),
.Y(n_1146)
);

NAND3xp33_ASAP7_75t_L g1147 ( 
.A(n_977),
.B(n_972),
.C(n_1030),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1006),
.Y(n_1148)
);

OA22x2_ASAP7_75t_L g1149 ( 
.A1(n_1080),
.A2(n_1088),
.B1(n_997),
.B2(n_954),
.Y(n_1149)
);

INVx1_ASAP7_75t_SL g1150 ( 
.A(n_956),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1040),
.B(n_996),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_1069),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1032),
.B(n_1029),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_995),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1035),
.B(n_1028),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_962),
.A2(n_1062),
.B(n_1038),
.C(n_970),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1059),
.A2(n_1049),
.B(n_1033),
.Y(n_1157)
);

AOI221xp5_ASAP7_75t_SL g1158 ( 
.A1(n_1051),
.A2(n_1036),
.B1(n_1050),
.B2(n_1057),
.C(n_967),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1036),
.B(n_1017),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1004),
.Y(n_1160)
);

AO31x2_ASAP7_75t_L g1161 ( 
.A1(n_958),
.A2(n_1056),
.A3(n_973),
.B(n_1027),
.Y(n_1161)
);

OA21x2_ASAP7_75t_L g1162 ( 
.A1(n_1063),
.A2(n_1058),
.B(n_1065),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1055),
.A2(n_1041),
.B(n_1095),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1039),
.B(n_1100),
.Y(n_1164)
);

NOR2xp67_ASAP7_75t_L g1165 ( 
.A(n_973),
.B(n_1027),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1039),
.B(n_1007),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_964),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_995),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1054),
.A2(n_1007),
.B1(n_1041),
.B2(n_1086),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1055),
.A2(n_1041),
.B(n_976),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_964),
.A2(n_976),
.B(n_1087),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1089),
.Y(n_1172)
);

AO21x2_ASAP7_75t_L g1173 ( 
.A1(n_1037),
.A2(n_1095),
.B(n_1087),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_1082),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_995),
.A2(n_1004),
.B(n_1086),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_SL g1176 ( 
.A1(n_1020),
.A2(n_1069),
.B1(n_1090),
.B2(n_1004),
.Y(n_1176)
);

INVxp67_ASAP7_75t_L g1177 ( 
.A(n_984),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1086),
.Y(n_1178)
);

AO21x2_ASAP7_75t_L g1179 ( 
.A1(n_995),
.A2(n_1044),
.B(n_992),
.Y(n_1179)
);

AO21x1_ASAP7_75t_L g1180 ( 
.A1(n_984),
.A2(n_1074),
.B(n_1073),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_959),
.A2(n_953),
.B(n_998),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1073),
.A2(n_1074),
.B(n_1092),
.C(n_1077),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_959),
.A2(n_953),
.B(n_998),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1018),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1084),
.B(n_1094),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1077),
.A2(n_1092),
.B(n_1074),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1003),
.B(n_797),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1084),
.B(n_1094),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_SL g1189 ( 
.A1(n_994),
.A2(n_918),
.B(n_780),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1003),
.B(n_797),
.Y(n_1190)
);

AOI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1053),
.A2(n_1060),
.B(n_1014),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1004),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_956),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_1003),
.B(n_797),
.Y(n_1194)
);

AO22x2_ASAP7_75t_L g1195 ( 
.A1(n_966),
.A2(n_1011),
.B1(n_986),
.B2(n_1067),
.Y(n_1195)
);

OR2x6_ASAP7_75t_L g1196 ( 
.A(n_1069),
.B(n_1067),
.Y(n_1196)
);

NAND2x1_ASAP7_75t_L g1197 ( 
.A(n_995),
.B(n_973),
.Y(n_1197)
);

CKINVDCx11_ASAP7_75t_R g1198 ( 
.A(n_1089),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_995),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1084),
.B(n_1094),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_959),
.A2(n_953),
.B(n_998),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1078),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_959),
.A2(n_953),
.B(n_998),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_956),
.Y(n_1204)
);

AO32x2_ASAP7_75t_L g1205 ( 
.A1(n_966),
.A2(n_1024),
.A3(n_1048),
.B1(n_1081),
.B2(n_1067),
.Y(n_1205)
);

O2A1O1Ixp5_ASAP7_75t_SL g1206 ( 
.A1(n_986),
.A2(n_989),
.B(n_1011),
.C(n_826),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_991),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_959),
.A2(n_953),
.B(n_998),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1073),
.A2(n_1074),
.B(n_1092),
.C(n_1077),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1084),
.A2(n_948),
.B1(n_798),
.B2(n_1094),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_995),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1084),
.B(n_1094),
.Y(n_1212)
);

NAND3xp33_ASAP7_75t_L g1213 ( 
.A(n_1077),
.B(n_1092),
.C(n_1074),
.Y(n_1213)
);

AOI31xp67_ASAP7_75t_L g1214 ( 
.A1(n_986),
.A2(n_1046),
.A3(n_1011),
.B(n_788),
.Y(n_1214)
);

BUFx2_ASAP7_75t_L g1215 ( 
.A(n_956),
.Y(n_1215)
);

AO21x1_ASAP7_75t_L g1216 ( 
.A1(n_1073),
.A2(n_1074),
.B(n_1011),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_959),
.A2(n_953),
.B(n_998),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_959),
.A2(n_953),
.B(n_998),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_1089),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_SL g1220 ( 
.A1(n_994),
.A2(n_918),
.B(n_780),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1004),
.Y(n_1221)
);

AOI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1053),
.A2(n_1060),
.B(n_1014),
.Y(n_1222)
);

NAND2x1p5_ASAP7_75t_L g1223 ( 
.A(n_973),
.B(n_1007),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_992),
.A2(n_1092),
.A3(n_1077),
.B(n_1048),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_982),
.A2(n_1097),
.B(n_983),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_992),
.A2(n_1092),
.A3(n_1077),
.B(n_1048),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1077),
.A2(n_1092),
.B(n_1074),
.Y(n_1227)
);

NOR2xp67_ASAP7_75t_L g1228 ( 
.A(n_973),
.B(n_796),
.Y(n_1228)
);

INVx5_ASAP7_75t_L g1229 ( 
.A(n_995),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_992),
.A2(n_1092),
.A3(n_1077),
.B(n_1048),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_959),
.A2(n_953),
.B(n_998),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_959),
.A2(n_953),
.B(n_998),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1084),
.B(n_1094),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_982),
.A2(n_1097),
.B(n_983),
.Y(n_1234)
);

AOI221x1_ASAP7_75t_L g1235 ( 
.A1(n_1077),
.A2(n_1092),
.B1(n_992),
.B2(n_969),
.C(n_841),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_992),
.A2(n_1092),
.A3(n_1077),
.B(n_1048),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1018),
.Y(n_1237)
);

AOI221xp5_ASAP7_75t_SL g1238 ( 
.A1(n_966),
.A2(n_981),
.B1(n_1073),
.B2(n_1074),
.C(n_826),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1004),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_959),
.A2(n_953),
.B(n_998),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_959),
.A2(n_953),
.B(n_998),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1078),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_959),
.A2(n_953),
.B(n_998),
.Y(n_1243)
);

INVxp67_ASAP7_75t_SL g1244 ( 
.A(n_1067),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1084),
.B(n_1094),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_959),
.A2(n_953),
.B(n_998),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1073),
.A2(n_1074),
.B(n_1092),
.C(n_1077),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1084),
.B(n_1094),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_982),
.A2(n_1097),
.B(n_983),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1084),
.B(n_1094),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_992),
.A2(n_1092),
.A3(n_1077),
.B(n_1048),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_982),
.A2(n_1097),
.B(n_983),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_959),
.A2(n_953),
.B(n_998),
.Y(n_1253)
);

BUFx8_ASAP7_75t_SL g1254 ( 
.A(n_1219),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1198),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_1172),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1135),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1185),
.A2(n_1212),
.B1(n_1245),
.B2(n_1210),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1210),
.A2(n_1108),
.B1(n_1141),
.B2(n_1107),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1112),
.Y(n_1260)
);

BUFx8_ASAP7_75t_L g1261 ( 
.A(n_1193),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1204),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1207),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1141),
.A2(n_1128),
.B1(n_1250),
.B2(n_1248),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_SL g1265 ( 
.A1(n_1188),
.A2(n_1233),
.B1(n_1200),
.B2(n_1176),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1187),
.A2(n_1190),
.B1(n_1194),
.B2(n_1139),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1115),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1151),
.A2(n_1116),
.B1(n_1111),
.B2(n_1147),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1138),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_1215),
.Y(n_1270)
);

INVx6_ASAP7_75t_L g1271 ( 
.A(n_1229),
.Y(n_1271)
);

INVx4_ASAP7_75t_L g1272 ( 
.A(n_1229),
.Y(n_1272)
);

INVx4_ASAP7_75t_L g1273 ( 
.A(n_1229),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1120),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1143),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1106),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1108),
.A2(n_1195),
.B1(n_1216),
.B2(n_1147),
.Y(n_1277)
);

CKINVDCx11_ASAP7_75t_R g1278 ( 
.A(n_1202),
.Y(n_1278)
);

INVx3_ASAP7_75t_SL g1279 ( 
.A(n_1150),
.Y(n_1279)
);

BUFx12f_ASAP7_75t_L g1280 ( 
.A(n_1110),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1113),
.Y(n_1281)
);

BUFx2_ASAP7_75t_SL g1282 ( 
.A(n_1242),
.Y(n_1282)
);

INVx8_ASAP7_75t_L g1283 ( 
.A(n_1160),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1127),
.Y(n_1284)
);

CKINVDCx11_ASAP7_75t_R g1285 ( 
.A(n_1150),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1121),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1103),
.A2(n_1116),
.B1(n_1174),
.B2(n_1238),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_1129),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_1153),
.Y(n_1289)
);

BUFx10_ASAP7_75t_L g1290 ( 
.A(n_1131),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1184),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1237),
.A2(n_1117),
.B1(n_1126),
.B2(n_1130),
.Y(n_1292)
);

OAI21xp33_ASAP7_75t_L g1293 ( 
.A1(n_1186),
.A2(n_1182),
.B(n_1209),
.Y(n_1293)
);

CKINVDCx11_ASAP7_75t_R g1294 ( 
.A(n_1174),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1195),
.A2(n_1213),
.B1(n_1124),
.B2(n_1227),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1146),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1149),
.A2(n_1213),
.B1(n_1227),
.B2(n_1176),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1180),
.A2(n_1196),
.B1(n_1244),
.B2(n_1122),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1196),
.A2(n_1155),
.B1(n_1247),
.B2(n_1164),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1148),
.Y(n_1300)
);

INVx4_ASAP7_75t_L g1301 ( 
.A(n_1160),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1196),
.A2(n_1220),
.B1(n_1189),
.B2(n_1179),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_SL g1303 ( 
.A(n_1146),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1159),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1144),
.B(n_1238),
.Y(n_1305)
);

INVx1_ASAP7_75t_SL g1306 ( 
.A(n_1131),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_SL g1307 ( 
.A1(n_1152),
.A2(n_1177),
.B1(n_1162),
.B2(n_1166),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1167),
.Y(n_1308)
);

CKINVDCx11_ASAP7_75t_R g1309 ( 
.A(n_1160),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1179),
.A2(n_1137),
.B1(n_1157),
.B2(n_1145),
.Y(n_1310)
);

CKINVDCx11_ASAP7_75t_R g1311 ( 
.A(n_1192),
.Y(n_1311)
);

INVx8_ASAP7_75t_L g1312 ( 
.A(n_1192),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1169),
.Y(n_1313)
);

BUFx12f_ASAP7_75t_L g1314 ( 
.A(n_1192),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1178),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1157),
.A2(n_1145),
.B1(n_1123),
.B2(n_1205),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1173),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1205),
.B(n_1221),
.Y(n_1318)
);

INVx11_ASAP7_75t_L g1319 ( 
.A(n_1221),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1221),
.Y(n_1320)
);

CKINVDCx11_ASAP7_75t_R g1321 ( 
.A(n_1239),
.Y(n_1321)
);

BUFx12f_ASAP7_75t_L g1322 ( 
.A(n_1239),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1173),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1171),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1239),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1142),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1156),
.A2(n_1228),
.B1(n_1134),
.B2(n_1165),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1123),
.A2(n_1205),
.B1(n_1228),
.B2(n_1162),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1197),
.Y(n_1329)
);

INVx6_ASAP7_75t_L g1330 ( 
.A(n_1223),
.Y(n_1330)
);

BUFx12f_ASAP7_75t_L g1331 ( 
.A(n_1140),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1132),
.A2(n_1211),
.B1(n_1199),
.B2(n_1168),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1132),
.A2(n_1168),
.B1(n_1211),
.B2(n_1199),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1175),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1154),
.Y(n_1335)
);

INVx1_ASAP7_75t_SL g1336 ( 
.A(n_1163),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1154),
.A2(n_1119),
.B1(n_1253),
.B2(n_1218),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_SL g1338 ( 
.A(n_1170),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1114),
.Y(n_1339)
);

BUFx4_ASAP7_75t_SL g1340 ( 
.A(n_1118),
.Y(n_1340)
);

INVx6_ASAP7_75t_L g1341 ( 
.A(n_1214),
.Y(n_1341)
);

BUFx12f_ASAP7_75t_L g1342 ( 
.A(n_1206),
.Y(n_1342)
);

INVx6_ASAP7_75t_L g1343 ( 
.A(n_1161),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1235),
.A2(n_1136),
.B1(n_1125),
.B2(n_1236),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1105),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1158),
.A2(n_1109),
.B1(n_1246),
.B2(n_1203),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1224),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1224),
.A2(n_1226),
.B1(n_1230),
.B2(n_1236),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1224),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1226),
.B(n_1251),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1226),
.A2(n_1251),
.B1(n_1230),
.B2(n_1236),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_1181),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1230),
.A2(n_1251),
.B1(n_1243),
.B2(n_1241),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1161),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_SL g1355 ( 
.A1(n_1183),
.A2(n_1240),
.B(n_1232),
.Y(n_1355)
);

CKINVDCx11_ASAP7_75t_R g1356 ( 
.A(n_1158),
.Y(n_1356)
);

CKINVDCx11_ASAP7_75t_R g1357 ( 
.A(n_1161),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1225),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1201),
.A2(n_1208),
.B1(n_1217),
.B2(n_1231),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1234),
.A2(n_1249),
.B1(n_1252),
.B2(n_1133),
.Y(n_1360)
);

CKINVDCx11_ASAP7_75t_R g1361 ( 
.A(n_1191),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1222),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1129),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1210),
.A2(n_426),
.B1(n_455),
.B2(n_413),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1104),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_1198),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1129),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1103),
.B(n_1185),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1229),
.Y(n_1369)
);

CKINVDCx6p67_ASAP7_75t_R g1370 ( 
.A(n_1198),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1104),
.Y(n_1371)
);

CKINVDCx11_ASAP7_75t_R g1372 ( 
.A(n_1198),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1210),
.A2(n_1141),
.B1(n_1108),
.B2(n_966),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1193),
.Y(n_1374)
);

INVx6_ASAP7_75t_L g1375 ( 
.A(n_1229),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1185),
.A2(n_1212),
.B1(n_1245),
.B2(n_1210),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1104),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1185),
.B(n_1212),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1185),
.A2(n_1212),
.B1(n_1245),
.B2(n_1210),
.Y(n_1379)
);

CKINVDCx11_ASAP7_75t_R g1380 ( 
.A(n_1198),
.Y(n_1380)
);

OAI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1210),
.A2(n_1141),
.B1(n_1108),
.B2(n_966),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_1198),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1185),
.A2(n_1212),
.B1(n_1245),
.B2(n_1210),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1185),
.A2(n_1212),
.B1(n_1245),
.B2(n_1210),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1104),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1104),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1104),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1345),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1254),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1350),
.B(n_1334),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1347),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1373),
.A2(n_1381),
.B1(n_1259),
.B2(n_1293),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1349),
.B(n_1316),
.Y(n_1393)
);

NAND2x1_ASAP7_75t_L g1394 ( 
.A(n_1343),
.B(n_1327),
.Y(n_1394)
);

BUFx4f_ASAP7_75t_L g1395 ( 
.A(n_1369),
.Y(n_1395)
);

INVx4_ASAP7_75t_L g1396 ( 
.A(n_1369),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1363),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1354),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1326),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1367),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1317),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1323),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1330),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1318),
.B(n_1316),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1351),
.B(n_1348),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1337),
.A2(n_1359),
.B(n_1360),
.Y(n_1406)
);

AOI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1268),
.A2(n_1362),
.B(n_1358),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1324),
.B(n_1339),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1288),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1330),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1279),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1329),
.B(n_1351),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1279),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1359),
.A2(n_1360),
.B(n_1355),
.Y(n_1414)
);

NAND2x1_ASAP7_75t_L g1415 ( 
.A(n_1341),
.B(n_1271),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1346),
.A2(n_1353),
.B(n_1310),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1260),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1373),
.A2(n_1381),
.B1(n_1259),
.B2(n_1297),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1365),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1371),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1387),
.Y(n_1421)
);

AO21x2_ASAP7_75t_L g1422 ( 
.A1(n_1305),
.A2(n_1299),
.B(n_1266),
.Y(n_1422)
);

AND2x4_ASAP7_75t_L g1423 ( 
.A(n_1302),
.B(n_1352),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1271),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1269),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1275),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1276),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1281),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1286),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1291),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1340),
.Y(n_1431)
);

OAI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1258),
.A2(n_1376),
.B(n_1383),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1328),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1328),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1295),
.B(n_1277),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1295),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1263),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1289),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1377),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1258),
.B(n_1376),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1277),
.B(n_1302),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1315),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_SL g1443 ( 
.A1(n_1265),
.A2(n_1307),
.B1(n_1331),
.B2(n_1378),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1331),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1385),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1386),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1310),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1357),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1353),
.A2(n_1333),
.B(n_1332),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1344),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1368),
.B(n_1298),
.Y(n_1451)
);

NAND2x1p5_ASAP7_75t_L g1452 ( 
.A(n_1272),
.B(n_1273),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1287),
.B(n_1298),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1335),
.A2(n_1292),
.B(n_1308),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1300),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1304),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1379),
.B(n_1384),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1342),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1296),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1342),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1264),
.B(n_1384),
.Y(n_1461)
);

AO21x2_ASAP7_75t_L g1462 ( 
.A1(n_1361),
.A2(n_1356),
.B(n_1325),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1320),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1379),
.A2(n_1383),
.B(n_1364),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1336),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1338),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1338),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1271),
.A2(n_1375),
.B(n_1273),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1375),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1330),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1262),
.B(n_1374),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1306),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1375),
.Y(n_1473)
);

O2A1O1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1464),
.A2(n_1267),
.B(n_1313),
.C(n_1284),
.Y(n_1474)
);

A2O1A1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1432),
.A2(n_1284),
.B(n_1274),
.C(n_1282),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1447),
.B(n_1370),
.Y(n_1476)
);

NAND2xp33_ASAP7_75t_R g1477 ( 
.A(n_1389),
.B(n_1255),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1418),
.A2(n_1270),
.B1(n_1303),
.B2(n_1256),
.Y(n_1478)
);

A2O1A1Ixp33_ASAP7_75t_L g1479 ( 
.A1(n_1392),
.A2(n_1257),
.B(n_1312),
.C(n_1283),
.Y(n_1479)
);

NOR2xp67_ASAP7_75t_L g1480 ( 
.A(n_1466),
.B(n_1280),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1456),
.B(n_1294),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1461),
.A2(n_1303),
.B1(n_1366),
.B2(n_1382),
.Y(n_1482)
);

OAI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1461),
.A2(n_1301),
.B(n_1280),
.Y(n_1483)
);

A2O1A1Ixp33_ASAP7_75t_L g1484 ( 
.A1(n_1443),
.A2(n_1312),
.B(n_1283),
.C(n_1290),
.Y(n_1484)
);

NOR2x1_ASAP7_75t_SL g1485 ( 
.A(n_1422),
.B(n_1314),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1408),
.B(n_1285),
.Y(n_1486)
);

INVx2_ASAP7_75t_SL g1487 ( 
.A(n_1471),
.Y(n_1487)
);

AOI221xp5_ASAP7_75t_L g1488 ( 
.A1(n_1440),
.A2(n_1301),
.B1(n_1312),
.B2(n_1283),
.C(n_1261),
.Y(n_1488)
);

OAI221xp5_ASAP7_75t_SL g1489 ( 
.A1(n_1457),
.A2(n_1380),
.B1(n_1372),
.B2(n_1261),
.C(n_1278),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1411),
.B(n_1309),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1451),
.B(n_1311),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1471),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1447),
.B(n_1321),
.Y(n_1493)
);

OA21x2_ASAP7_75t_L g1494 ( 
.A1(n_1414),
.A2(n_1314),
.B(n_1322),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1423),
.B(n_1322),
.Y(n_1495)
);

OA21x2_ASAP7_75t_L g1496 ( 
.A1(n_1414),
.A2(n_1319),
.B(n_1406),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_SL g1497 ( 
.A(n_1399),
.B(n_1467),
.Y(n_1497)
);

O2A1O1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1453),
.A2(n_1466),
.B(n_1458),
.C(n_1422),
.Y(n_1498)
);

NOR2x1_ASAP7_75t_SL g1499 ( 
.A(n_1422),
.B(n_1462),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1394),
.A2(n_1465),
.B(n_1416),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1431),
.A2(n_1423),
.B(n_1435),
.C(n_1394),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1413),
.B(n_1399),
.Y(n_1502)
);

AND2x6_ASAP7_75t_L g1503 ( 
.A(n_1444),
.B(n_1412),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1390),
.B(n_1428),
.Y(n_1504)
);

BUFx8_ASAP7_75t_SL g1505 ( 
.A(n_1399),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1404),
.B(n_1393),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1409),
.B(n_1472),
.Y(n_1507)
);

AOI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1435),
.A2(n_1436),
.B1(n_1441),
.B2(n_1450),
.C(n_1438),
.Y(n_1508)
);

OAI211xp5_ASAP7_75t_SL g1509 ( 
.A1(n_1458),
.A2(n_1448),
.B(n_1431),
.C(n_1436),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1441),
.A2(n_1423),
.B1(n_1462),
.B2(n_1448),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1406),
.A2(n_1454),
.B(n_1449),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1423),
.A2(n_1462),
.B1(n_1465),
.B2(n_1450),
.Y(n_1512)
);

AOI221xp5_ASAP7_75t_L g1513 ( 
.A1(n_1433),
.A2(n_1434),
.B1(n_1405),
.B2(n_1397),
.C(n_1400),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1454),
.A2(n_1468),
.B(n_1449),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1468),
.A2(n_1460),
.B(n_1452),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1442),
.B(n_1425),
.Y(n_1516)
);

AO32x2_ASAP7_75t_L g1517 ( 
.A1(n_1403),
.A2(n_1470),
.A3(n_1410),
.B1(n_1396),
.B2(n_1390),
.Y(n_1517)
);

O2A1O1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1459),
.A2(n_1460),
.B(n_1463),
.C(n_1403),
.Y(n_1518)
);

OA21x2_ASAP7_75t_L g1519 ( 
.A1(n_1407),
.A2(n_1398),
.B(n_1401),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1425),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1426),
.B(n_1427),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1437),
.B(n_1455),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1439),
.B(n_1445),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1427),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1395),
.A2(n_1410),
.B1(n_1470),
.B2(n_1424),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1439),
.B(n_1445),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1395),
.A2(n_1424),
.B1(n_1469),
.B2(n_1433),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1519),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1511),
.B(n_1391),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1524),
.Y(n_1530)
);

OAI222xp33_ASAP7_75t_L g1531 ( 
.A1(n_1510),
.A2(n_1429),
.B1(n_1430),
.B2(n_1446),
.C1(n_1460),
.C2(n_1415),
.Y(n_1531)
);

NOR2xp67_ASAP7_75t_L g1532 ( 
.A(n_1500),
.B(n_1515),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1506),
.B(n_1402),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1517),
.B(n_1504),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1517),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1520),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1514),
.B(n_1391),
.Y(n_1537)
);

NAND4xp25_ASAP7_75t_L g1538 ( 
.A(n_1508),
.B(n_1446),
.C(n_1460),
.D(n_1420),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1515),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1496),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1478),
.A2(n_1412),
.B1(n_1473),
.B2(n_1421),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1516),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1503),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_L g1544 ( 
.A(n_1498),
.B(n_1419),
.C(n_1417),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1521),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1522),
.Y(n_1546)
);

NOR2xp67_ASAP7_75t_L g1547 ( 
.A(n_1523),
.B(n_1401),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1526),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1512),
.B(n_1388),
.Y(n_1549)
);

INVx5_ASAP7_75t_L g1550 ( 
.A(n_1503),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1494),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1499),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1550),
.B(n_1503),
.Y(n_1553)
);

INVx2_ASAP7_75t_SL g1554 ( 
.A(n_1550),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1548),
.B(n_1485),
.Y(n_1555)
);

AO21x2_ASAP7_75t_L g1556 ( 
.A1(n_1528),
.A2(n_1512),
.B(n_1407),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1529),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1529),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1537),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1529),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1529),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1536),
.Y(n_1562)
);

NOR2x1_ASAP7_75t_SL g1563 ( 
.A(n_1550),
.B(n_1527),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1530),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1535),
.B(n_1412),
.Y(n_1565)
);

OAI31xp33_ASAP7_75t_L g1566 ( 
.A1(n_1538),
.A2(n_1501),
.A3(n_1475),
.B(n_1479),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1546),
.B(n_1513),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1547),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1535),
.B(n_1487),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1535),
.B(n_1492),
.Y(n_1570)
);

AOI211xp5_ASAP7_75t_SL g1571 ( 
.A1(n_1531),
.A2(n_1484),
.B(n_1489),
.C(n_1482),
.Y(n_1571)
);

NAND4xp25_ASAP7_75t_L g1572 ( 
.A(n_1538),
.B(n_1482),
.C(n_1474),
.D(n_1481),
.Y(n_1572)
);

OAI33xp33_ASAP7_75t_L g1573 ( 
.A1(n_1549),
.A2(n_1509),
.A3(n_1493),
.B1(n_1476),
.B2(n_1518),
.B3(n_1525),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1541),
.A2(n_1497),
.B1(n_1488),
.B2(n_1491),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1541),
.A2(n_1507),
.B1(n_1486),
.B2(n_1495),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1553),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1562),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1568),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1568),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1554),
.Y(n_1580)
);

NOR2x1_ASAP7_75t_L g1581 ( 
.A(n_1556),
.B(n_1544),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1562),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1557),
.B(n_1534),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1557),
.B(n_1540),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1564),
.Y(n_1585)
);

NOR4xp25_ASAP7_75t_SL g1586 ( 
.A(n_1571),
.B(n_1543),
.C(n_1539),
.D(n_1477),
.Y(n_1586)
);

NOR2x1_ASAP7_75t_L g1587 ( 
.A(n_1556),
.B(n_1544),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1558),
.B(n_1539),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1567),
.B(n_1545),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1562),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1567),
.B(n_1545),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1558),
.B(n_1532),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1559),
.B(n_1532),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1558),
.B(n_1532),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1560),
.B(n_1549),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1555),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1553),
.Y(n_1597)
);

NOR4xp25_ASAP7_75t_SL g1598 ( 
.A(n_1571),
.B(n_1543),
.C(n_1551),
.D(n_1552),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1560),
.B(n_1533),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1561),
.B(n_1533),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1567),
.B(n_1545),
.Y(n_1601)
);

AND2x2_ASAP7_75t_SL g1602 ( 
.A(n_1553),
.B(n_1543),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1553),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1585),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1589),
.B(n_1570),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1602),
.B(n_1565),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1585),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1589),
.B(n_1573),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1602),
.B(n_1565),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1584),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1577),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1577),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1577),
.Y(n_1613)
);

INVx2_ASAP7_75t_SL g1614 ( 
.A(n_1602),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1602),
.B(n_1565),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1591),
.B(n_1542),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1582),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1591),
.B(n_1542),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1582),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1576),
.B(n_1565),
.Y(n_1620)
);

NAND2x1p5_ASAP7_75t_L g1621 ( 
.A(n_1581),
.B(n_1550),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1601),
.B(n_1564),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1576),
.B(n_1563),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1576),
.B(n_1554),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1601),
.B(n_1570),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1578),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1578),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1579),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1579),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1596),
.B(n_1555),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1576),
.B(n_1563),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1596),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1582),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1597),
.A2(n_1573),
.B1(n_1572),
.B2(n_1566),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1590),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1592),
.B(n_1555),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1597),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1590),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1590),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1592),
.B(n_1569),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1599),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1597),
.B(n_1563),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1597),
.B(n_1572),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1592),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1584),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1599),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1606),
.B(n_1603),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1608),
.B(n_1595),
.Y(n_1648)
);

XNOR2xp5_ASAP7_75t_L g1649 ( 
.A(n_1634),
.B(n_1572),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1606),
.B(n_1603),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1607),
.B(n_1595),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1610),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1609),
.B(n_1603),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1609),
.B(n_1603),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1615),
.B(n_1593),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1607),
.B(n_1595),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_1626),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1615),
.B(n_1593),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1611),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1604),
.B(n_1599),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1643),
.B(n_1505),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1632),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1614),
.B(n_1593),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1627),
.B(n_1583),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1612),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1622),
.B(n_1592),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1628),
.Y(n_1668)
);

NOR3xp33_ASAP7_75t_L g1669 ( 
.A(n_1614),
.B(n_1587),
.C(n_1581),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1612),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1616),
.B(n_1490),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1610),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1620),
.B(n_1594),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1629),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1620),
.B(n_1594),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1605),
.B(n_1600),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1644),
.A2(n_1574),
.B1(n_1497),
.B2(n_1575),
.Y(n_1677)
);

AOI211xp5_ASAP7_75t_L g1678 ( 
.A1(n_1630),
.A2(n_1566),
.B(n_1586),
.C(n_1574),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1645),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1637),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1605),
.B(n_1600),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1613),
.Y(n_1682)
);

AOI31xp33_ASAP7_75t_L g1683 ( 
.A1(n_1649),
.A2(n_1571),
.A3(n_1621),
.B(n_1502),
.Y(n_1683)
);

AOI222xp33_ASAP7_75t_L g1684 ( 
.A1(n_1649),
.A2(n_1587),
.B1(n_1581),
.B2(n_1575),
.C1(n_1588),
.C2(n_1636),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1647),
.B(n_1637),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1647),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1651),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1663),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1662),
.B(n_1671),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1650),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1651),
.Y(n_1691)
);

AOI222xp33_ASAP7_75t_L g1692 ( 
.A1(n_1648),
.A2(n_1587),
.B1(n_1588),
.B2(n_1594),
.C1(n_1618),
.C2(n_1640),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1648),
.B(n_1625),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1650),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1674),
.B(n_1625),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1678),
.A2(n_1574),
.B1(n_1623),
.B2(n_1642),
.Y(n_1696)
);

OAI21xp33_ASAP7_75t_L g1697 ( 
.A1(n_1677),
.A2(n_1594),
.B(n_1641),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1679),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_1654),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1658),
.B(n_1645),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1660),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1660),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1666),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1666),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1678),
.A2(n_1598),
.B(n_1586),
.Y(n_1705)
);

AOI21xp33_ASAP7_75t_R g1706 ( 
.A1(n_1653),
.A2(n_1637),
.B(n_1641),
.Y(n_1706)
);

AOI32xp33_ASAP7_75t_L g1707 ( 
.A1(n_1669),
.A2(n_1631),
.A3(n_1642),
.B1(n_1623),
.B2(n_1588),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1654),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1705),
.A2(n_1668),
.B1(n_1658),
.B2(n_1677),
.C(n_1652),
.Y(n_1709)
);

OAI31xp33_ASAP7_75t_L g1710 ( 
.A1(n_1697),
.A2(n_1668),
.A3(n_1621),
.B(n_1655),
.Y(n_1710)
);

OAI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1683),
.A2(n_1621),
.B(n_1680),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1688),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1688),
.B(n_1656),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1685),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1684),
.B(n_1680),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1686),
.B(n_1655),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1696),
.A2(n_1667),
.B1(n_1656),
.B2(n_1659),
.Y(n_1717)
);

A2O1A1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1707),
.A2(n_1566),
.B(n_1659),
.C(n_1631),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1694),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1692),
.B(n_1653),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1689),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1694),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1693),
.A2(n_1598),
.B(n_1652),
.Y(n_1723)
);

A2O1A1Ixp33_ASAP7_75t_L g1724 ( 
.A1(n_1698),
.A2(n_1657),
.B(n_1483),
.C(n_1480),
.Y(n_1724)
);

OAI21xp33_ASAP7_75t_L g1725 ( 
.A1(n_1699),
.A2(n_1664),
.B(n_1665),
.Y(n_1725)
);

AOI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1700),
.A2(n_1657),
.B(n_1653),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1702),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1686),
.B(n_1687),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1716),
.B(n_1687),
.Y(n_1729)
);

INVx2_ASAP7_75t_SL g1730 ( 
.A(n_1714),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1709),
.A2(n_1708),
.B1(n_1691),
.B2(n_1695),
.Y(n_1731)
);

AOI21xp33_ASAP7_75t_SL g1732 ( 
.A1(n_1715),
.A2(n_1708),
.B(n_1691),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1713),
.Y(n_1733)
);

AOI221xp5_ASAP7_75t_L g1734 ( 
.A1(n_1715),
.A2(n_1706),
.B1(n_1701),
.B2(n_1690),
.C(n_1702),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1712),
.Y(n_1735)
);

NAND2x1p5_ASAP7_75t_L g1736 ( 
.A(n_1714),
.B(n_1685),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1720),
.A2(n_1664),
.B1(n_1673),
.B2(n_1675),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1721),
.B(n_1673),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1720),
.A2(n_1672),
.B(n_1703),
.Y(n_1739)
);

NOR3xp33_ASAP7_75t_L g1740 ( 
.A(n_1734),
.B(n_1723),
.C(n_1728),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_L g1741 ( 
.A(n_1732),
.B(n_1717),
.C(n_1711),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1736),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1730),
.Y(n_1743)
);

NAND4xp25_ASAP7_75t_L g1744 ( 
.A(n_1738),
.B(n_1710),
.C(n_1718),
.D(n_1725),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1735),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1729),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1735),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1731),
.A2(n_1726),
.B1(n_1672),
.B2(n_1675),
.Y(n_1748)
);

OAI211xp5_ASAP7_75t_L g1749 ( 
.A1(n_1740),
.A2(n_1739),
.B(n_1733),
.C(n_1737),
.Y(n_1749)
);

O2A1O1Ixp5_ASAP7_75t_L g1750 ( 
.A1(n_1742),
.A2(n_1724),
.B(n_1672),
.C(n_1722),
.Y(n_1750)
);

AOI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1740),
.A2(n_1724),
.B1(n_1727),
.B2(n_1719),
.C(n_1704),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1744),
.B(n_1746),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1743),
.Y(n_1753)
);

OAI221xp5_ASAP7_75t_SL g1754 ( 
.A1(n_1749),
.A2(n_1748),
.B1(n_1741),
.B2(n_1745),
.C(n_1747),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1752),
.B(n_1703),
.Y(n_1755)
);

XOR2xp5_ASAP7_75t_L g1756 ( 
.A(n_1753),
.B(n_1704),
.Y(n_1756)
);

O2A1O1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1750),
.A2(n_1682),
.B(n_1670),
.C(n_1661),
.Y(n_1757)
);

INVx1_ASAP7_75t_SL g1758 ( 
.A(n_1751),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1751),
.B(n_1661),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1756),
.Y(n_1760)
);

INVxp67_ASAP7_75t_L g1761 ( 
.A(n_1759),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1758),
.B(n_1665),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1755),
.B(n_1757),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1754),
.B(n_1682),
.Y(n_1764)
);

NAND2x1p5_ASAP7_75t_L g1765 ( 
.A(n_1760),
.B(n_1480),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1761),
.A2(n_1670),
.B1(n_1624),
.B2(n_1681),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1764),
.A2(n_1681),
.B1(n_1676),
.B2(n_1624),
.Y(n_1767)
);

NOR2xp67_ASAP7_75t_SL g1768 ( 
.A(n_1765),
.B(n_1763),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1768),
.Y(n_1769)
);

XNOR2xp5_ASAP7_75t_L g1770 ( 
.A(n_1769),
.B(n_1762),
.Y(n_1770)
);

XNOR2x1_ASAP7_75t_SL g1771 ( 
.A(n_1769),
.B(n_1766),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1770),
.A2(n_1767),
.B1(n_1676),
.B2(n_1646),
.Y(n_1772)
);

OAI22x1_ASAP7_75t_SL g1773 ( 
.A1(n_1771),
.A2(n_1646),
.B1(n_1580),
.B2(n_1619),
.Y(n_1773)
);

INVxp67_ASAP7_75t_L g1774 ( 
.A(n_1773),
.Y(n_1774)
);

AOI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1772),
.A2(n_1617),
.B(n_1613),
.Y(n_1775)
);

AOI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1774),
.A2(n_1624),
.B1(n_1580),
.B2(n_1619),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1776),
.B(n_1775),
.Y(n_1777)
);

AOI22x1_ASAP7_75t_L g1778 ( 
.A1(n_1777),
.A2(n_1639),
.B1(n_1617),
.B2(n_1633),
.Y(n_1778)
);

OAI221xp5_ASAP7_75t_R g1779 ( 
.A1(n_1778),
.A2(n_1580),
.B1(n_1633),
.B2(n_1639),
.C(n_1638),
.Y(n_1779)
);

AOI211xp5_ASAP7_75t_L g1780 ( 
.A1(n_1779),
.A2(n_1635),
.B(n_1580),
.C(n_1552),
.Y(n_1780)
);


endmodule