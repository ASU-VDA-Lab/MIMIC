module fake_jpeg_12284_n_170 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_170);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_49),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_29),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_24),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_19),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_8),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_6),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_82),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_80),
.Y(n_88)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_77),
.Y(n_91)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_18),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_1),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_55),
.C(n_2),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_59),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_94),
.Y(n_103)
);

NAND2x1p5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_51),
.Y(n_106)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_58),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_60),
.B1(n_64),
.B2(n_62),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_96),
.B1(n_73),
.B2(n_65),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_60),
.B1(n_64),
.B2(n_62),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_73),
.B1(n_56),
.B2(n_65),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_104),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_66),
.B1(n_70),
.B2(n_69),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_111),
.B1(n_114),
.B2(n_118),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_12),
.B(n_13),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_68),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_52),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_58),
.B1(n_72),
.B2(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_54),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_12),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_53),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_22),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_23),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_5),
.C(n_7),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_125),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_25),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_131),
.C(n_21),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_113),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_105),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_37),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_139),
.B1(n_14),
.B2(n_20),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_134),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_32),
.C(n_42),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_103),
.A2(n_115),
.B(n_117),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_35),
.B(n_36),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_142),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_140),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_145),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_140),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_31),
.B(n_33),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_146),
.A2(n_149),
.B(n_154),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_152),
.A2(n_153),
.B1(n_135),
.B2(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_38),
.B(n_39),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_147),
.A2(n_128),
.B1(n_122),
.B2(n_129),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_159),
.A2(n_154),
.B(n_146),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_133),
.C(n_124),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_161),
.B(n_162),
.Y(n_164)
);

AOI21x1_ASAP7_75t_L g162 ( 
.A1(n_160),
.A2(n_143),
.B(n_149),
.Y(n_162)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_158),
.A3(n_156),
.B1(n_157),
.B2(n_135),
.C1(n_155),
.C2(n_150),
.Y(n_165)
);

BUFx24_ASAP7_75t_SL g166 ( 
.A(n_165),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_148),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_120),
.B(n_142),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_164),
.C(n_131),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_169),
.B(n_50),
.Y(n_170)
);


endmodule