module real_aes_4951_n_9 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_1, n_9);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_1;
output n_9;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_23;
wire n_20;
wire n_18;
wire n_21;
wire n_10;
AOI321xp33_ASAP7_75t_L g9 ( .A1(n_0), .A2(n_7), .A3(n_10), .B1(n_12), .B2(n_13), .C(n_24), .Y(n_9) );
OAI321xp33_ASAP7_75t_L g13 ( .A1(n_1), .A2(n_10), .A3(n_14), .B1(n_15), .B2(n_16), .C(n_23), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
BUFx6f_ASAP7_75t_L g20 ( .A(n_3), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_4), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_5), .Y(n_21) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
INVx1_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_10), .Y(n_15) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
CKINVDCx20_ASAP7_75t_R g23 ( .A(n_12), .Y(n_23) );
NOR2xp33_ASAP7_75t_L g25 ( .A(n_12), .B(n_15), .Y(n_25) );
NOR2xp33_ASAP7_75t_L g24 ( .A(n_13), .B(n_25), .Y(n_24) );
AOI22xp5_ASAP7_75t_L g16 ( .A1(n_17), .A2(n_18), .B1(n_21), .B2(n_22), .Y(n_16) );
INVx2_ASAP7_75t_SL g17 ( .A(n_18), .Y(n_17) );
BUFx2_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
endmodule