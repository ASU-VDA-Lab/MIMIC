module fake_jpeg_18705_n_298 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_51),
.B(n_18),
.Y(n_66)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_9),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_44),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

CKINVDCx9p33_ASAP7_75t_R g47 ( 
.A(n_25),
.Y(n_47)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_52),
.B(n_36),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_36),
.C(n_38),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_88),
.Y(n_108)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_54),
.Y(n_109)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_59),
.Y(n_106)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_63),
.Y(n_112)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_26),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_65),
.B(n_67),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_66),
.Y(n_119)
);

OR2x2_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_25),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_17),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_72),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_44),
.A2(n_33),
.B(n_9),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_70),
.Y(n_131)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_17),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_21),
.B1(n_22),
.B2(n_26),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_76),
.A2(n_97),
.B1(n_100),
.B2(n_20),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_19),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_77),
.Y(n_117)
);

CKINVDCx12_ASAP7_75t_R g79 ( 
.A(n_40),
.Y(n_79)
);

NAND2x1_ASAP7_75t_SL g107 ( 
.A(n_79),
.B(n_84),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_22),
.B1(n_21),
.B2(n_38),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_81),
.B1(n_87),
.B2(n_20),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_45),
.A2(n_21),
.B1(n_22),
.B2(n_38),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_83),
.A2(n_85),
.B1(n_91),
.B2(n_101),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_18),
.B1(n_24),
.B2(n_29),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_90),
.Y(n_110)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_45),
.B(n_23),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_41),
.B(n_37),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_41),
.A2(n_37),
.B1(n_35),
.B2(n_32),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_35),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_34),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_41),
.A2(n_32),
.B1(n_23),
.B2(n_28),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_28),
.B1(n_24),
.B2(n_29),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_103),
.B1(n_111),
.B2(n_56),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_29),
.B1(n_24),
.B2(n_27),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_126),
.B1(n_129),
.B2(n_61),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_66),
.A2(n_0),
.B(n_1),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_121),
.Y(n_158)
);

OR2x4_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_132),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_80),
.A2(n_101),
.B1(n_85),
.B2(n_87),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_95),
.A2(n_34),
.B1(n_20),
.B2(n_27),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_70),
.B1(n_64),
.B2(n_84),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_82),
.A2(n_34),
.B1(n_27),
.B2(n_10),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_123),
.B(n_16),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_133),
.B(n_160),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_58),
.B1(n_60),
.B2(n_56),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_142),
.B1(n_146),
.B2(n_150),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_135),
.A2(n_143),
.B1(n_118),
.B2(n_107),
.Y(n_178)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_136),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_113),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_137),
.B(n_147),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_122),
.B(n_61),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_139),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_98),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_70),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_145),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_98),
.B1(n_94),
.B2(n_73),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_144),
.A2(n_109),
.B1(n_131),
.B2(n_120),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_117),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_119),
.A2(n_94),
.B1(n_89),
.B2(n_74),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_122),
.B(n_108),
.Y(n_147)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_148),
.A2(n_136),
.B1(n_109),
.B2(n_114),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_10),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_152),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_119),
.A2(n_89),
.B1(n_74),
.B2(n_2),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_10),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_113),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_105),
.A2(n_74),
.B1(n_1),
.B2(n_3),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_161),
.B1(n_165),
.B2(n_14),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_0),
.B(n_1),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_156),
.A2(n_159),
.B(n_164),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_12),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_12),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_108),
.B(n_5),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_162),
.B(n_14),
.CI(n_15),
.CON(n_196),
.SN(n_196)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_121),
.A2(n_6),
.B(n_9),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_102),
.A2(n_6),
.B1(n_12),
.B2(n_13),
.Y(n_165)
);

AND2x6_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_107),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_167),
.B(n_196),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_139),
.C(n_140),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_176),
.C(n_150),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_151),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_171),
.Y(n_211)
);

CKINVDCx10_ASAP7_75t_R g171 ( 
.A(n_136),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_182),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_132),
.C(n_110),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_SL g177 ( 
.A1(n_158),
.A2(n_129),
.B(n_115),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_177),
.A2(n_184),
.B(n_197),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_185),
.B1(n_191),
.B2(n_142),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_163),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_186),
.A2(n_144),
.B1(n_152),
.B2(n_149),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_110),
.B(n_107),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_188),
.A2(n_193),
.B(n_133),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_138),
.B(n_106),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_192),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_135),
.A2(n_106),
.B1(n_109),
.B2(n_114),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_141),
.B(n_110),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_164),
.B(n_157),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_145),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_104),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_114),
.B(n_16),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_210),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_202),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_159),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_146),
.C(n_134),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_216),
.C(n_190),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_183),
.A2(n_159),
.B(n_153),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_207),
.B(n_188),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_205),
.A2(n_202),
.B1(n_208),
.B2(n_203),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_155),
.B1(n_161),
.B2(n_165),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_206),
.A2(n_186),
.B1(n_166),
.B2(n_193),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_183),
.A2(n_143),
.B(n_137),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_159),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_212),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_159),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_215),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_148),
.C(n_130),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_166),
.A2(n_148),
.B1(n_130),
.B2(n_104),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_219),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_194),
.B(n_15),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_218),
.B(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_187),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_174),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_221),
.A2(n_228),
.B1(n_236),
.B2(n_239),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_235),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_167),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_230),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_205),
.A2(n_187),
.B1(n_182),
.B2(n_185),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_176),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_199),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_206),
.A2(n_170),
.B1(n_190),
.B2(n_195),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_171),
.B(n_180),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_207),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_181),
.Y(n_238)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

BUFx12_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

BUFx12_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_245),
.A2(n_209),
.B(n_234),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_216),
.C(n_201),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_233),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_249),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_198),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_222),
.B(n_218),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_251),
.Y(n_267)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_198),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_212),
.C(n_232),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_254),
.A2(n_221),
.B1(n_228),
.B2(n_236),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_255),
.B(n_257),
.Y(n_270)
);

AOI22x1_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_237),
.B1(n_204),
.B2(n_231),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_247),
.B(n_169),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_264),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_254),
.A2(n_222),
.B1(n_227),
.B2(n_234),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_213),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_253),
.B(n_172),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g269 ( 
.A(n_261),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_216),
.C(n_232),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_266),
.C(n_248),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_265),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_249),
.C(n_252),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_273),
.C(n_262),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_244),
.C(n_241),
.Y(n_273)
);

OAI322xp33_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_210),
.A3(n_201),
.B1(n_244),
.B2(n_196),
.C1(n_209),
.C2(n_235),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_274),
.A2(n_213),
.B(n_268),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_260),
.A2(n_180),
.B1(n_229),
.B2(n_217),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_277),
.B1(n_258),
.B2(n_211),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_278),
.B(n_279),
.Y(n_290)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_277),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_280),
.A2(n_219),
.B1(n_211),
.B2(n_263),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_270),
.A2(n_259),
.B(n_256),
.C(n_255),
.Y(n_281)
);

O2A1O1Ixp33_ASAP7_75t_SL g285 ( 
.A1(n_281),
.A2(n_275),
.B(n_242),
.C(n_240),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_282),
.B(n_284),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_266),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_200),
.C(n_215),
.Y(n_288)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_242),
.C(n_197),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_286),
.B(n_195),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_278),
.C(n_240),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_269),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_282),
.B1(n_214),
.B2(n_283),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_291),
.Y(n_295)
);

AO21x2_ASAP7_75t_L g296 ( 
.A1(n_292),
.A2(n_293),
.B(n_294),
.Y(n_296)
);

OAI21x1_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_287),
.B(n_290),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_295),
.Y(n_298)
);


endmodule