module fake_jpeg_3071_n_179 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_63),
.B(n_50),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

BUFx2_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_66),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_65),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_56),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_75),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_42),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_46),
.B(n_45),
.C(n_60),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_44),
.B1(n_60),
.B2(n_58),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_78),
.Y(n_92)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_56),
.C(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_85),
.Y(n_99)
);

OR2x2_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_83),
.B(n_84),
.Y(n_112)
);

AOI32xp33_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_42),
.A3(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_86),
.Y(n_111)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_64),
.B1(n_65),
.B2(n_47),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_80),
.B1(n_61),
.B2(n_72),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_55),
.C(n_52),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_7),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_51),
.B1(n_18),
.B2(n_20),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_54),
.A3(n_53),
.B1(n_57),
.B2(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_0),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_114),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_72),
.B1(n_67),
.B2(n_58),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_103),
.A2(n_104),
.B1(n_109),
.B2(n_6),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_64),
.B1(n_47),
.B2(n_43),
.Y(n_104)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_51),
.B1(n_1),
.B2(n_2),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_51),
.B1(n_1),
.B2(n_2),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_128),
.B1(n_129),
.B2(n_9),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_106),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_102),
.B(n_3),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_125),
.Y(n_148)
);

A2O1A1O1Ixp25_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_39),
.B(n_38),
.C(n_36),
.D(n_34),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_106),
.B(n_24),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_126),
.C(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_33),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_121),
.B(n_122),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_111),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_32),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_12),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_112),
.B(n_99),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_111),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_31),
.B1(n_30),
.B2(n_26),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_25),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_131),
.B(n_132),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_98),
.B(n_7),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_8),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_12),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_145),
.B1(n_119),
.B2(n_15),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_138),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_9),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_140),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_10),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_115),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_141),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_11),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_143),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_144),
.Y(n_160)
);

OAI321xp33_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_23),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_116),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_148),
.B(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_154),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_141),
.A2(n_13),
.B1(n_16),
.B2(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_157),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_139),
.B(n_144),
.Y(n_157)
);

AOI221xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_136),
.B1(n_148),
.B2(n_139),
.C(n_150),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_147),
.B1(n_153),
.B2(n_160),
.Y(n_164)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_164),
.B(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_151),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_159),
.C(n_152),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_170),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_171),
.A2(n_164),
.B1(n_165),
.B2(n_163),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_168),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_173),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_177),
.B(n_172),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_155),
.Y(n_179)
);


endmodule