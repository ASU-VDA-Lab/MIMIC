module fake_jpeg_15064_n_360 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_360);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_60),
.Y(n_64)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_32),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_66),
.Y(n_117)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_72),
.B(n_86),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_85),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_25),
.B1(n_43),
.B2(n_35),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_80),
.B1(n_91),
.B2(n_35),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_33),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_84),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_25),
.B1(n_43),
.B2(n_35),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_38),
.C(n_23),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_39),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_20),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_59),
.A2(n_25),
.B1(n_43),
.B2(n_30),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_33),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_89),
.B(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_45),
.B(n_20),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_60),
.A2(n_35),
.B1(n_31),
.B2(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_31),
.B1(n_30),
.B2(n_21),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_SL g104 ( 
.A1(n_84),
.A2(n_38),
.B(n_21),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_121),
.B(n_26),
.C(n_29),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_105),
.Y(n_139)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_108),
.A2(n_48),
.B1(n_46),
.B2(n_76),
.Y(n_144)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_111),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_67),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_31),
.B1(n_35),
.B2(n_21),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_69),
.B1(n_81),
.B2(n_72),
.Y(n_142)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_116),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_68),
.A2(n_31),
.B1(n_63),
.B2(n_61),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_34),
.B1(n_56),
.B2(n_62),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_79),
.B(n_22),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_123),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

BUFx24_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_67),
.A2(n_22),
.B(n_34),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_39),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_64),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_62),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_102),
.B1(n_110),
.B2(n_123),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_87),
.B1(n_69),
.B2(n_92),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_144),
.B1(n_156),
.B2(n_109),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_138),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_38),
.B(n_93),
.C(n_73),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_133),
.A2(n_134),
.B(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_95),
.Y(n_140)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_34),
.A3(n_26),
.B1(n_42),
.B2(n_29),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_42),
.A3(n_117),
.B1(n_96),
.B2(n_41),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_117),
.Y(n_161)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_78),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

AO22x1_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_73),
.B1(n_58),
.B2(n_47),
.Y(n_152)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_125),
.B(n_44),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_157),
.A2(n_53),
.B(n_65),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_119),
.B1(n_96),
.B2(n_108),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_158),
.A2(n_179),
.B1(n_129),
.B2(n_156),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_177),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_161),
.B(n_165),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_163),
.B1(n_145),
.B2(n_151),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_114),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_170),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_132),
.B(n_101),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_172),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_133),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_152),
.Y(n_197)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

OAI32xp33_ASAP7_75t_L g177 ( 
.A1(n_131),
.A2(n_47),
.A3(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_113),
.B1(n_107),
.B2(n_54),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_140),
.C(n_138),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_182),
.C(n_187),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_128),
.C(n_137),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_175),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_186),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_178),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_128),
.C(n_137),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_188),
.A2(n_191),
.B1(n_167),
.B2(n_177),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_157),
.C(n_141),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_196),
.C(n_201),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_157),
.B1(n_134),
.B2(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_157),
.C(n_139),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_197),
.A2(n_176),
.B(n_179),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_200),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_139),
.C(n_129),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_185),
.A2(n_166),
.B1(n_180),
.B2(n_164),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_206),
.B1(n_223),
.B2(n_118),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_192),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_207),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_164),
.Y(n_204)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_185),
.A2(n_180),
.B1(n_174),
.B2(n_158),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_160),
.C(n_176),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_168),
.Y(n_211)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_184),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_122),
.Y(n_240)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_222),
.B1(n_76),
.B2(n_71),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_195),
.A2(n_191),
.B(n_188),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_219),
.A2(n_154),
.B(n_120),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_172),
.C(n_162),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_199),
.C(n_154),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_195),
.A2(n_152),
.B1(n_143),
.B2(n_150),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_224),
.B(n_41),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_189),
.A2(n_135),
.B1(n_150),
.B2(n_136),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_135),
.B1(n_146),
.B2(n_136),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_198),
.A2(n_146),
.B(n_172),
.Y(n_224)
);

AOI32xp33_ASAP7_75t_SL g225 ( 
.A1(n_189),
.A2(n_118),
.A3(n_154),
.B1(n_23),
.B2(n_37),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_225),
.A2(n_199),
.B1(n_193),
.B2(n_148),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_227),
.A2(n_230),
.B(n_231),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_182),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_232),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_244),
.C(n_246),
.Y(n_254)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_0),
.B(n_1),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_154),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_235),
.B(n_223),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_238),
.A2(n_249),
.B1(n_220),
.B2(n_213),
.Y(n_266)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_120),
.B(n_16),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_243),
.A2(n_248),
.B(n_227),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_65),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_245),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_65),
.C(n_120),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_211),
.B(n_23),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_247),
.B(n_225),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_209),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_65),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_203),
.C(n_208),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_224),
.Y(n_251)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_257),
.B1(n_248),
.B2(n_249),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_236),
.B(n_204),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_265),
.Y(n_291)
);

AO32x1_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_216),
.A3(n_221),
.B1(n_202),
.B2(n_206),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_238),
.Y(n_265)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_268),
.C(n_244),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_228),
.B(n_217),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_241),
.Y(n_269)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_233),
.B(n_222),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_270),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_229),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_271),
.A2(n_231),
.B(n_250),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_272),
.B(n_66),
.Y(n_289)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_265),
.A2(n_271),
.B1(n_257),
.B2(n_234),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_275),
.A2(n_287),
.B1(n_258),
.B2(n_262),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_37),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_232),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_280),
.C(n_284),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_279),
.B(n_289),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_246),
.C(n_247),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_208),
.C(n_205),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_254),
.A2(n_205),
.B1(n_230),
.B2(n_1),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_258),
.A2(n_263),
.B1(n_266),
.B2(n_254),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_288),
.A2(n_272),
.B1(n_260),
.B2(n_261),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_256),
.A2(n_41),
.B1(n_37),
.B2(n_36),
.Y(n_292)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_292),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_264),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_293),
.B(n_298),
.C(n_299),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_297),
.B(n_289),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_286),
.A2(n_261),
.B1(n_260),
.B2(n_41),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_37),
.C(n_36),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_307),
.C(n_282),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_283),
.A2(n_13),
.B(n_4),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_306),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_305),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_277),
.B(n_13),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_36),
.C(n_32),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_278),
.B(n_12),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_308),
.B(n_12),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_314),
.C(n_317),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_294),
.A2(n_291),
.B1(n_274),
.B2(n_282),
.Y(n_311)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_279),
.B(n_290),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_312),
.A2(n_301),
.B(n_305),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_300),
.A2(n_275),
.B1(n_287),
.B2(n_280),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_321),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_302),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_318),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_281),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_15),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_322),
.C(n_9),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_301),
.B(n_15),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_307),
.A2(n_36),
.B1(n_32),
.B2(n_28),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_304),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_323),
.B(n_326),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_295),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_333),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_309),
.A2(n_296),
.B1(n_32),
.B2(n_28),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_327),
.A2(n_321),
.B1(n_6),
.B2(n_7),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_330),
.B(n_331),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_9),
.C(n_4),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_2),
.C(n_5),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_313),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_340),
.Y(n_346)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_325),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_339),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_324),
.A2(n_316),
.B1(n_327),
.B2(n_329),
.Y(n_338)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_338),
.Y(n_343)
);

NAND3xp33_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_5),
.C(n_6),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_6),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_342),
.B(n_329),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_345),
.A2(n_347),
.B(n_337),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_7),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_335),
.B(n_19),
.C(n_8),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_348),
.B(n_9),
.C(n_11),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_349),
.B(n_350),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_346),
.A2(n_7),
.B(n_8),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_351),
.A2(n_352),
.B(n_344),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_343),
.A2(n_11),
.B(n_15),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_354),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_355),
.Y(n_356)
);

A2O1A1Ixp33_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_353),
.B(n_348),
.C(n_18),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_16),
.C(n_17),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_358),
.B(n_19),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_16),
.C(n_18),
.Y(n_360)
);


endmodule