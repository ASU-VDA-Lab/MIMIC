module fake_ariane_91_n_1099 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_32, n_28, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_1099);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_32;
input n_28;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_1099;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_160;
wire n_64;
wire n_180;
wire n_730;
wire n_119;
wire n_124;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_423;
wire n_347;
wire n_1042;
wire n_961;
wire n_183;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_133;
wire n_610;
wire n_66;
wire n_205;
wire n_752;
wire n_341;
wire n_71;
wire n_1029;
wire n_985;
wire n_109;
wire n_245;
wire n_421;
wire n_96;
wire n_549;
wire n_522;
wire n_319;
wire n_49;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_50;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_103;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_72;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_57;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_117;
wire n_139;
wire n_524;
wire n_85;
wire n_130;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_515;
wire n_379;
wire n_807;
wire n_445;
wire n_138;
wire n_162;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_137;
wire n_885;
wire n_122;
wire n_198;
wire n_232;
wire n_52;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_73;
wire n_327;
wire n_77;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_87;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_41;
wire n_813;
wire n_926;
wire n_140;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_900;
wire n_154;
wire n_883;
wire n_338;
wire n_142;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_145;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_731;
wire n_59;
wire n_336;
wire n_754;
wire n_665;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_54;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_167;
wire n_90;
wire n_38;
wire n_422;
wire n_47;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_75;
wire n_1018;
wire n_855;
wire n_158;
wire n_1047;
wire n_69;
wire n_259;
wire n_835;
wire n_95;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_143;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_115;
wire n_331;
wire n_559;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_721;
wire n_840;
wire n_600;
wire n_1053;
wire n_1084;
wire n_398;
wire n_62;
wire n_210;
wire n_1090;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_839;
wire n_79;
wire n_821;
wire n_928;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_825;
wire n_567;
wire n_732;
wire n_91;
wire n_971;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_44;
wire n_82;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_604;
wire n_677;
wire n_614;
wire n_439;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_48;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_129;
wire n_126;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_93;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_108;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_168;
wire n_81;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_455;
wire n_365;
wire n_654;
wire n_429;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_136;
wire n_334;
wire n_192;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_163;
wire n_88;
wire n_869;
wire n_141;
wire n_846;
wire n_390;
wire n_498;
wire n_104;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_56;
wire n_60;
wire n_728;
wire n_388;
wire n_449;
wire n_612;
wire n_957;
wire n_413;
wire n_977;
wire n_333;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_685;
wire n_911;
wire n_221;
wire n_321;
wire n_459;
wire n_86;
wire n_458;
wire n_361;
wire n_89;
wire n_149;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_74;
wire n_491;
wire n_810;
wire n_40;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_53;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_46;
wire n_772;
wire n_741;
wire n_747;
wire n_84;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_107;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_42;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_1038;
wire n_70;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_680;
wire n_571;
wire n_287;
wire n_302;
wire n_993;
wire n_948;
wire n_380;
wire n_582;
wire n_94;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_58;
wire n_37;
wire n_65;
wire n_123;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_135;
wire n_1033;
wire n_896;
wire n_409;
wire n_171;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_61;
wire n_526;
wire n_742;
wire n_102;
wire n_716;
wire n_182;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_196;
wire n_125;
wire n_798;
wire n_769;
wire n_820;
wire n_43;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_55;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_848;
wire n_574;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_68;
wire n_415;
wire n_794;
wire n_763;
wire n_78;
wire n_63;
wire n_655;
wire n_99;
wire n_540;
wire n_216;
wire n_692;
wire n_544;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_83;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_951;
wire n_1026;
wire n_213;
wire n_938;
wire n_862;
wire n_110;
wire n_304;
wire n_895;
wire n_659;
wire n_67;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_92;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_98;
wire n_946;
wire n_757;
wire n_375;
wire n_113;
wire n_114;
wire n_324;
wire n_1030;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_697;
wire n_437;
wire n_111;
wire n_274;
wire n_622;
wire n_967;
wire n_337;
wire n_999;
wire n_998;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_174;
wire n_275;
wire n_100;
wire n_704;
wire n_1060;
wire n_132;
wire n_1044;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_51;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_76;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_159;
wire n_1002;
wire n_580;
wire n_105;
wire n_358;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_131;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_165;
wire n_1037;
wire n_144;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_101;
wire n_243;
wire n_803;
wire n_134;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_112;
wire n_45;
wire n_548;
wire n_815;
wire n_542;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_650;
wire n_258;
wire n_782;
wire n_856;
wire n_364;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_121;
wire n_118;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_484;
wire n_712;
wire n_411;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_80;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_1011;
wire n_97;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_116;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_39;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_796;
wire n_805;
wire n_127;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_28),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_12),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_34),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_19),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_22),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_0),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_11),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

BUFx8_ASAP7_75t_SL g75 ( 
.A(n_44),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_2),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_2),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_4),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_5),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_56),
.Y(n_88)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_70),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_70),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_57),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_63),
.B(n_60),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_R g97 ( 
.A(n_83),
.B(n_69),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_52),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_83),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_80),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_80),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_R g110 ( 
.A(n_83),
.B(n_66),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_83),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_83),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_80),
.Y(n_114)
);

BUFx6f_ASAP7_75t_SL g115 ( 
.A(n_89),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_95),
.B(n_83),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_82),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_82),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_77),
.Y(n_124)
);

NOR3xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_51),
.C(n_52),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_77),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_77),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_82),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_77),
.Y(n_132)
);

AO221x1_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_60),
.B1(n_55),
.B2(n_63),
.C(n_53),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_77),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_82),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_82),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_77),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_77),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_97),
.B(n_77),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_77),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g151 ( 
.A(n_90),
.B(n_55),
.C(n_53),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_82),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_82),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_82),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_97),
.B(n_81),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_110),
.B(n_81),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_110),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_92),
.Y(n_160)
);

AND2x6_ASAP7_75t_SL g161 ( 
.A(n_93),
.B(n_82),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_95),
.B(n_81),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_90),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_98),
.B(n_82),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_98),
.B(n_81),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_98),
.B(n_81),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_121),
.A2(n_81),
.B1(n_80),
.B2(n_79),
.Y(n_169)
);

OR2x6_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_81),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_81),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_140),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_81),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_140),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_140),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_126),
.B(n_81),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_164),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_126),
.B(n_79),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_47),
.Y(n_184)
);

AO22x1_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_46),
.B1(n_49),
.B2(n_45),
.Y(n_185)
);

OR2x2_ASAP7_75t_SL g186 ( 
.A(n_148),
.B(n_40),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

AND2x4_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_40),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_48),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_121),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_121),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_74),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_140),
.B(n_79),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_146),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_140),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_130),
.B(n_141),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_140),
.B(n_79),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_42),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_140),
.B(n_144),
.Y(n_202)
);

BUFx4f_ASAP7_75t_L g203 ( 
.A(n_144),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_140),
.B(n_79),
.Y(n_204)
);

NOR2xp67_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_86),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_141),
.B(n_74),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_119),
.B(n_74),
.Y(n_207)
);

NOR2x2_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_54),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_120),
.B(n_74),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_118),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_147),
.B(n_150),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_164),
.Y(n_212)
);

AND3x2_ASAP7_75t_SL g213 ( 
.A(n_161),
.B(n_62),
.C(n_64),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_121),
.B(n_79),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_134),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_150),
.B(n_79),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

NAND2x1p5_ASAP7_75t_L g218 ( 
.A(n_131),
.B(n_86),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_SL g219 ( 
.A(n_131),
.B(n_58),
.C(n_59),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_124),
.A2(n_85),
.B(n_87),
.Y(n_220)
);

CKINVDCx11_ASAP7_75t_R g221 ( 
.A(n_160),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_118),
.Y(n_223)
);

NOR2x1p5_ASAP7_75t_L g224 ( 
.A(n_129),
.B(n_38),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_115),
.A2(n_74),
.B1(n_79),
.B2(n_61),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_153),
.B(n_79),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_SL g227 ( 
.A(n_125),
.B(n_37),
.C(n_67),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_132),
.A2(n_72),
.B1(n_71),
.B2(n_68),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_153),
.B(n_79),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_118),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_127),
.B(n_73),
.Y(n_232)
);

NAND2x1_ASAP7_75t_L g233 ( 
.A(n_118),
.B(n_85),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_168),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_115),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_128),
.B(n_79),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_152),
.A2(n_85),
.B(n_87),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_138),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_133),
.A2(n_79),
.B1(n_74),
.B2(n_86),
.Y(n_239)
);

BUFx4f_ASAP7_75t_L g240 ( 
.A(n_118),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_135),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_136),
.Y(n_242)
);

BUFx4f_ASAP7_75t_L g243 ( 
.A(n_128),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_182),
.A2(n_43),
.B1(n_42),
.B2(n_142),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_162),
.Y(n_246)
);

NOR2xp67_ASAP7_75t_SL g247 ( 
.A(n_174),
.B(n_139),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_170),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_195),
.B(n_159),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_158),
.B(n_156),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_182),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_159),
.Y(n_253)
);

AOI21x1_ASAP7_75t_L g254 ( 
.A1(n_216),
.A2(n_230),
.B(n_226),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_219),
.A2(n_198),
.B1(n_232),
.B2(n_241),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

AND2x4_ASAP7_75t_L g257 ( 
.A(n_170),
.B(n_174),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_243),
.A2(n_137),
.B(n_139),
.C(n_138),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_228),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_201),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_R g261 ( 
.A(n_212),
.B(n_115),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_215),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_192),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g264 ( 
.A(n_170),
.B(n_143),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_177),
.B(n_117),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_212),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_215),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_243),
.A2(n_155),
.B(n_154),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_240),
.A2(n_85),
.B(n_87),
.Y(n_269)
);

O2A1O1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_211),
.A2(n_43),
.B(n_133),
.C(n_78),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_229),
.B(n_79),
.Y(n_271)
);

AOI22x1_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_79),
.B1(n_74),
.B2(n_76),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_172),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_240),
.A2(n_87),
.B(n_74),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_SL g275 ( 
.A1(n_184),
.A2(n_78),
.B(n_76),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_223),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_202),
.A2(n_87),
.B(n_74),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_190),
.B(n_79),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_188),
.B(n_79),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_202),
.A2(n_87),
.B(n_74),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_174),
.A2(n_79),
.B1(n_74),
.B2(n_87),
.Y(n_281)
);

NOR3xp33_ASAP7_75t_SL g282 ( 
.A(n_227),
.B(n_213),
.C(n_171),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_223),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_218),
.A2(n_74),
.B1(n_86),
.B2(n_65),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_188),
.B(n_74),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_187),
.B(n_74),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g288 ( 
.A(n_221),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_223),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_188),
.B(n_74),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_187),
.A2(n_74),
.B1(n_87),
.B2(n_78),
.Y(n_291)
);

OAI21x1_ASAP7_75t_L g292 ( 
.A1(n_214),
.A2(n_78),
.B(n_76),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_200),
.B(n_86),
.Y(n_293)
);

OAI21xp33_ASAP7_75t_L g294 ( 
.A1(n_189),
.A2(n_74),
.B(n_76),
.Y(n_294)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_187),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_205),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_186),
.A2(n_86),
.B1(n_8),
.B2(n_10),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_236),
.A2(n_78),
.B(n_76),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_217),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_236),
.A2(n_78),
.B(n_76),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_223),
.A2(n_78),
.B1(n_76),
.B2(n_86),
.Y(n_301)
);

O2A1O1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_206),
.A2(n_78),
.B(n_76),
.C(n_65),
.Y(n_302)
);

A2O1A1Ixp33_ASAP7_75t_L g303 ( 
.A1(n_203),
.A2(n_78),
.B(n_76),
.C(n_86),
.Y(n_303)
);

BUFx4f_ASAP7_75t_L g304 ( 
.A(n_231),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_176),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_224),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_217),
.B(n_65),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_221),
.B(n_6),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_192),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_237),
.A2(n_78),
.B(n_76),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_238),
.B(n_86),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_238),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_231),
.A2(n_78),
.B1(n_76),
.B2(n_86),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_180),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_210),
.B(n_86),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_252),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_262),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_252),
.Y(n_318)
);

OAI21x1_ASAP7_75t_L g319 ( 
.A1(n_254),
.A2(n_191),
.B(n_180),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_245),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_266),
.B(n_185),
.Y(n_321)
);

CKINVDCx8_ASAP7_75t_R g322 ( 
.A(n_257),
.Y(n_322)
);

OA21x2_ASAP7_75t_L g323 ( 
.A1(n_258),
.A2(n_183),
.B(n_193),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_287),
.B(n_169),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_248),
.B(n_191),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_275),
.A2(n_207),
.B(n_209),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_260),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_262),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_288),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_263),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_257),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

OAI21x1_ASAP7_75t_L g333 ( 
.A1(n_254),
.A2(n_214),
.B(n_181),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_263),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_244),
.B(n_192),
.Y(n_335)
);

BUFx12f_ASAP7_75t_L g336 ( 
.A(n_288),
.Y(n_336)
);

AO21x2_ASAP7_75t_L g337 ( 
.A1(n_268),
.A2(n_175),
.B(n_199),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_263),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_257),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_248),
.B(n_192),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_255),
.B(n_264),
.Y(n_341)
);

CKINVDCx6p67_ASAP7_75t_R g342 ( 
.A(n_259),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_267),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_287),
.B(n_210),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_267),
.Y(n_345)
);

BUFx4f_ASAP7_75t_L g346 ( 
.A(n_256),
.Y(n_346)
);

AO21x2_ASAP7_75t_L g347 ( 
.A1(n_278),
.A2(n_194),
.B(n_199),
.Y(n_347)
);

BUFx2_ASAP7_75t_R g348 ( 
.A(n_245),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_299),
.Y(n_349)
);

AO21x2_ASAP7_75t_L g350 ( 
.A1(n_251),
.A2(n_194),
.B(n_204),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_261),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_259),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_304),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_249),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_299),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_312),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_249),
.B(n_210),
.Y(n_357)
);

AOI21x1_ASAP7_75t_L g358 ( 
.A1(n_247),
.A2(n_233),
.B(n_220),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_263),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

INVx4_ASAP7_75t_SL g361 ( 
.A(n_309),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_246),
.B(n_231),
.Y(n_362)
);

BUFx4_ASAP7_75t_SL g363 ( 
.A(n_276),
.Y(n_363)
);

AOI22x1_ASAP7_75t_L g364 ( 
.A1(n_269),
.A2(n_231),
.B1(n_197),
.B2(n_173),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_314),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_255),
.B(n_203),
.Y(n_366)
);

OAI21x1_ASAP7_75t_L g367 ( 
.A1(n_302),
.A2(n_204),
.B(n_239),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_264),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_273),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_273),
.Y(n_370)
);

OAI21x1_ASAP7_75t_L g371 ( 
.A1(n_272),
.A2(n_225),
.B(n_203),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_264),
.A2(n_179),
.B1(n_173),
.B2(n_197),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_293),
.B(n_86),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_314),
.Y(n_375)
);

OAI21x1_ASAP7_75t_L g376 ( 
.A1(n_272),
.A2(n_178),
.B(n_179),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_279),
.Y(n_377)
);

OAI21x1_ASAP7_75t_L g378 ( 
.A1(n_292),
.A2(n_178),
.B(n_213),
.Y(n_378)
);

OAI21x1_ASAP7_75t_L g379 ( 
.A1(n_292),
.A2(n_208),
.B(n_86),
.Y(n_379)
);

INVx6_ASAP7_75t_L g380 ( 
.A(n_309),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_275),
.A2(n_235),
.B(n_86),
.Y(n_381)
);

AOI22x1_ASAP7_75t_L g382 ( 
.A1(n_309),
.A2(n_235),
.B1(n_208),
.B2(n_13),
.Y(n_382)
);

BUFx12f_ASAP7_75t_L g383 ( 
.A(n_309),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_305),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_285),
.Y(n_386)
);

AO21x2_ASAP7_75t_L g387 ( 
.A1(n_315),
.A2(n_86),
.B(n_36),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_290),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_253),
.B(n_86),
.Y(n_389)
);

OAI21x1_ASAP7_75t_L g390 ( 
.A1(n_307),
.A2(n_86),
.B(n_33),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

INVx8_ASAP7_75t_L g392 ( 
.A(n_256),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_304),
.Y(n_393)
);

BUFx4f_ASAP7_75t_SL g394 ( 
.A(n_276),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_382),
.A2(n_297),
.B1(n_308),
.B2(n_293),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_384),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_384),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

OAI22xp33_ASAP7_75t_L g399 ( 
.A1(n_341),
.A2(n_250),
.B1(n_306),
.B2(n_295),
.Y(n_399)
);

CKINVDCx11_ASAP7_75t_R g400 ( 
.A(n_336),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_328),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_328),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g403 ( 
.A(n_318),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_391),
.A2(n_341),
.B1(n_373),
.B2(n_335),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_384),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_326),
.A2(n_271),
.B(n_303),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_383),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g409 ( 
.A1(n_391),
.A2(n_296),
.B1(n_284),
.B2(n_294),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_328),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_345),
.Y(n_411)
);

NOR2x1_ASAP7_75t_L g412 ( 
.A(n_366),
.B(n_289),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_385),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_327),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_345),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_385),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_SL g417 ( 
.A1(n_382),
.A2(n_270),
.B1(n_282),
.B2(n_295),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_320),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_320),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_385),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_336),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_354),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_369),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_324),
.B(n_368),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_369),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_363),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_331),
.B(n_339),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_370),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_383),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_321),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_345),
.Y(n_431)
);

OR2x6_ASAP7_75t_L g432 ( 
.A(n_368),
.B(n_289),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_370),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_317),
.Y(n_435)
);

AO21x1_ASAP7_75t_L g436 ( 
.A1(n_366),
.A2(n_286),
.B(n_301),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_353),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_324),
.A2(n_295),
.B1(n_86),
.B2(n_256),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_353),
.Y(n_439)
);

CKINVDCx11_ASAP7_75t_R g440 ( 
.A(n_336),
.Y(n_440)
);

BUFx12f_ASAP7_75t_L g441 ( 
.A(n_351),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_331),
.B(n_283),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_317),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_343),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_356),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_373),
.A2(n_313),
.B1(n_283),
.B2(n_295),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_383),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_354),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_343),
.Y(n_449)
);

OA21x2_ASAP7_75t_L g450 ( 
.A1(n_319),
.A2(n_274),
.B(n_277),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_349),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_331),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_377),
.A2(n_295),
.B1(n_304),
.B2(n_300),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_316),
.Y(n_454)
);

CKINVDCx11_ASAP7_75t_R g455 ( 
.A(n_342),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_330),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_326),
.A2(n_281),
.B(n_298),
.Y(n_457)
);

BUFx12f_ASAP7_75t_L g458 ( 
.A(n_329),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_356),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_339),
.B(n_280),
.Y(n_460)
);

AOI21x1_ASAP7_75t_L g461 ( 
.A1(n_323),
.A2(n_247),
.B(n_310),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_349),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_377),
.A2(n_291),
.B1(n_8),
.B2(n_13),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_356),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_339),
.B(n_30),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_386),
.A2(n_6),
.B1(n_14),
.B2(n_15),
.Y(n_466)
);

OAI22xp33_ASAP7_75t_R g467 ( 
.A1(n_342),
.A2(n_16),
.B1(n_18),
.B2(n_23),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_355),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_355),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_360),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_394),
.Y(n_471)
);

OAI21x1_ASAP7_75t_SL g472 ( 
.A1(n_381),
.A2(n_340),
.B(n_325),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_322),
.A2(n_325),
.B1(n_340),
.B2(n_357),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_405),
.B(n_344),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_414),
.B(n_342),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_424),
.B(n_423),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_473),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_424),
.B(n_348),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_423),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_419),
.B(n_344),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_418),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_396),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_396),
.Y(n_483)
);

OR2x6_ASAP7_75t_L g484 ( 
.A(n_473),
.B(n_386),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_419),
.B(n_418),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_454),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_471),
.Y(n_487)
);

AND2x6_ASAP7_75t_L g488 ( 
.A(n_465),
.B(n_334),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_422),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_R g491 ( 
.A(n_465),
.B(n_323),
.Y(n_491)
);

OR2x6_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_432),
.Y(n_492)
);

NAND3xp33_ASAP7_75t_SL g493 ( 
.A(n_395),
.B(n_403),
.C(n_352),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_425),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_455),
.Y(n_495)
);

NAND3xp33_ASAP7_75t_SL g496 ( 
.A(n_395),
.B(n_322),
.C(n_362),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_422),
.A2(n_322),
.B1(n_346),
.B2(n_357),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_425),
.B(n_357),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_428),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_397),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_R g501 ( 
.A(n_465),
.B(n_323),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_400),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_448),
.B(n_348),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_458),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_428),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_406),
.Y(n_506)
);

INVx3_ASAP7_75t_SL g507 ( 
.A(n_421),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_R g508 ( 
.A(n_471),
.B(n_353),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_406),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_448),
.B(n_357),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_430),
.B(n_434),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_426),
.B(n_16),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_434),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_440),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_435),
.Y(n_515)
);

OR2x6_ASAP7_75t_L g516 ( 
.A(n_472),
.B(n_319),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_R g517 ( 
.A(n_441),
.B(n_393),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_435),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_433),
.B(n_427),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_443),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_427),
.B(n_442),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_SL g522 ( 
.A1(n_467),
.A2(n_387),
.B1(n_388),
.B2(n_381),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_466),
.A2(n_346),
.B1(n_372),
.B2(n_393),
.Y(n_523)
);

A2O1A1Ixp33_ASAP7_75t_L g524 ( 
.A1(n_407),
.A2(n_372),
.B(n_371),
.C(n_346),
.Y(n_524)
);

NOR3xp33_ASAP7_75t_SL g525 ( 
.A(n_467),
.B(n_389),
.C(n_388),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_413),
.B(n_323),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_404),
.B(n_375),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_413),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_443),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_444),
.Y(n_530)
);

INVx5_ASAP7_75t_L g531 ( 
.A(n_456),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_R g532 ( 
.A(n_465),
.B(n_323),
.Y(n_532)
);

OR2x6_ASAP7_75t_L g533 ( 
.A(n_432),
.B(n_319),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_442),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_R g535 ( 
.A(n_441),
.B(n_393),
.Y(n_535)
);

NOR3xp33_ASAP7_75t_SL g536 ( 
.A(n_399),
.B(n_389),
.C(n_23),
.Y(n_536)
);

A2O1A1Ixp33_ASAP7_75t_SL g537 ( 
.A1(n_457),
.A2(n_338),
.B(n_374),
.C(n_365),
.Y(n_537)
);

NOR2xp67_ASAP7_75t_L g538 ( 
.A(n_441),
.B(n_338),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_416),
.B(n_420),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_452),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_492),
.B(n_456),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_482),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_476),
.B(n_416),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_482),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_526),
.B(n_420),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_516),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_492),
.B(n_456),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_476),
.B(n_444),
.Y(n_548)
);

OA21x2_ASAP7_75t_L g549 ( 
.A1(n_524),
.A2(n_390),
.B(n_436),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_483),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_526),
.B(n_456),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_489),
.B(n_449),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_534),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_492),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_492),
.Y(n_555)
);

A2O1A1Ixp33_ASAP7_75t_L g556 ( 
.A1(n_525),
.A2(n_417),
.B(n_407),
.C(n_457),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_533),
.B(n_456),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_483),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_490),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_490),
.Y(n_560)
);

AOI33xp33_ASAP7_75t_L g561 ( 
.A1(n_522),
.A2(n_463),
.A3(n_417),
.B1(n_25),
.B2(n_27),
.B3(n_24),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_488),
.Y(n_562)
);

AO21x2_ASAP7_75t_L g563 ( 
.A1(n_537),
.A2(n_436),
.B(n_461),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_488),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_485),
.B(n_449),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_500),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_500),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_516),
.B(n_456),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_516),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_506),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_506),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_509),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_509),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_528),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_528),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_493),
.A2(n_438),
.B1(n_427),
.B2(n_446),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_516),
.B(n_412),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_533),
.B(n_462),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_515),
.Y(n_579)
);

INVxp67_ASAP7_75t_SL g580 ( 
.A(n_491),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_518),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_498),
.B(n_412),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_520),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_533),
.B(n_477),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_529),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_533),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_530),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_479),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_481),
.B(n_451),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_494),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_499),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_498),
.B(n_450),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_505),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_513),
.B(n_451),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_488),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_524),
.B(n_450),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_539),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_480),
.B(n_469),
.Y(n_598)
);

INVx5_ASAP7_75t_L g599 ( 
.A(n_488),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_531),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_511),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_531),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_531),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_521),
.B(n_450),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_601),
.B(n_474),
.Y(n_605)
);

NAND3xp33_ASAP7_75t_L g606 ( 
.A(n_561),
.B(n_536),
.C(n_491),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_550),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_550),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_604),
.B(n_551),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_588),
.B(n_537),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_553),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_601),
.B(n_510),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_604),
.B(n_484),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_601),
.B(n_540),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_553),
.B(n_519),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_587),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_588),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_593),
.B(n_484),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_593),
.B(n_484),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_550),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_556),
.A2(n_484),
.B1(n_475),
.B2(n_438),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_587),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_604),
.B(n_503),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_548),
.B(n_486),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_597),
.B(n_531),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_599),
.B(n_531),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_548),
.B(n_507),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_551),
.B(n_478),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_587),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_565),
.Y(n_630)
);

INVxp67_ASAP7_75t_SL g631 ( 
.A(n_580),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_587),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_599),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_584),
.B(n_527),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_597),
.B(n_488),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_551),
.B(n_488),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_592),
.B(n_487),
.Y(n_637)
);

OAI22xp5_ASAP7_75t_L g638 ( 
.A1(n_556),
.A2(n_523),
.B1(n_497),
.B2(n_504),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_592),
.B(n_487),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_552),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_599),
.B(n_538),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_565),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_550),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_592),
.B(n_545),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_599),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_597),
.B(n_462),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_597),
.B(n_468),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_545),
.B(n_512),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_598),
.B(n_468),
.Y(n_649)
);

OAI21xp33_ASAP7_75t_L g650 ( 
.A1(n_561),
.A2(n_496),
.B(n_508),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_590),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_590),
.Y(n_652)
);

AND2x4_ASAP7_75t_SL g653 ( 
.A(n_562),
.B(n_432),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_598),
.B(n_469),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_545),
.B(n_461),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_590),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_598),
.B(n_470),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_582),
.B(n_532),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_590),
.Y(n_659)
);

NAND3xp33_ASAP7_75t_L g660 ( 
.A(n_549),
.B(n_532),
.C(n_501),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_582),
.B(n_501),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_609),
.B(n_596),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_616),
.Y(n_663)
);

OR2x6_ASAP7_75t_L g664 ( 
.A(n_660),
.B(n_595),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_637),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_631),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_609),
.B(n_596),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_616),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_640),
.B(n_591),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_644),
.B(n_596),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_644),
.B(n_580),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_617),
.Y(n_672)
);

AND2x2_ASAP7_75t_SL g673 ( 
.A(n_653),
.B(n_595),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_622),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_642),
.B(n_591),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_605),
.B(n_565),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_613),
.B(n_595),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_622),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_611),
.B(n_591),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_629),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_607),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_613),
.B(n_568),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_629),
.B(n_591),
.Y(n_683)
);

AND2x2_ASAP7_75t_SL g684 ( 
.A(n_653),
.B(n_562),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_637),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_632),
.B(n_589),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_623),
.B(n_568),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_607),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_607),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_605),
.B(n_552),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_623),
.B(n_568),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_634),
.B(n_584),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_655),
.B(n_546),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_634),
.B(n_584),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_612),
.B(n_543),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_633),
.B(n_599),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_632),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_633),
.B(n_599),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_651),
.B(n_652),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_651),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_610),
.Y(n_701)
);

OAI31xp33_ASAP7_75t_L g702 ( 
.A1(n_606),
.A2(n_578),
.A3(n_495),
.B(n_586),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_655),
.B(n_546),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_639),
.B(n_569),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_608),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_652),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_608),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_639),
.B(n_569),
.Y(n_708)
);

NAND2x1_ASAP7_75t_L g709 ( 
.A(n_633),
.B(n_562),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_608),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_620),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_636),
.B(n_557),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_610),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_656),
.B(n_589),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_636),
.B(n_557),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_656),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_615),
.B(n_543),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_659),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_658),
.B(n_661),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_620),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_620),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_658),
.B(n_557),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_661),
.B(n_557),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_628),
.B(n_557),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_628),
.B(n_557),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_614),
.B(n_578),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_659),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_648),
.B(n_577),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_654),
.B(n_579),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_630),
.Y(n_730)
);

A2O1A1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_702),
.A2(n_606),
.B(n_650),
.C(n_660),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_673),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_688),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_679),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_679),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_701),
.B(n_648),
.Y(n_736)
);

OAI322xp33_ASAP7_75t_L g737 ( 
.A1(n_690),
.A2(n_638),
.A3(n_654),
.B1(n_649),
.B2(n_621),
.C1(n_624),
.C2(n_657),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_688),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_662),
.B(n_627),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_669),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_692),
.B(n_618),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_669),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_672),
.Y(n_743)
);

OAI22xp33_ASAP7_75t_L g744 ( 
.A1(n_664),
.A2(n_638),
.B1(n_621),
.B2(n_599),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_702),
.A2(n_650),
.B1(n_576),
.B2(n_549),
.Y(n_745)
);

OAI31xp33_ASAP7_75t_L g746 ( 
.A1(n_701),
.A2(n_586),
.A3(n_657),
.B(n_635),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_662),
.B(n_618),
.Y(n_747)
);

AOI21xp33_ASAP7_75t_SL g748 ( 
.A1(n_730),
.A2(n_502),
.B(n_514),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_692),
.B(n_619),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_672),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_676),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_701),
.Y(n_752)
);

NAND2x2_ASAP7_75t_L g753 ( 
.A(n_709),
.B(n_554),
.Y(n_753)
);

OAI21xp33_ASAP7_75t_SL g754 ( 
.A1(n_662),
.A2(n_619),
.B(n_633),
.Y(n_754)
);

A2O1A1Ixp33_ASAP7_75t_L g755 ( 
.A1(n_666),
.A2(n_719),
.B(n_576),
.C(n_673),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_730),
.B(n_507),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_688),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_676),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_713),
.B(n_625),
.Y(n_759)
);

NAND4xp75_ASAP7_75t_L g760 ( 
.A(n_684),
.B(n_645),
.C(n_586),
.D(n_549),
.Y(n_760)
);

NAND5xp2_ASAP7_75t_L g761 ( 
.A(n_666),
.B(n_577),
.C(n_585),
.D(n_579),
.E(n_581),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_676),
.Y(n_762)
);

NAND4xp75_ASAP7_75t_L g763 ( 
.A(n_684),
.B(n_645),
.C(n_549),
.D(n_555),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_713),
.B(n_690),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_713),
.B(n_625),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_664),
.A2(n_577),
.B1(n_582),
.B2(n_555),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_724),
.B(n_626),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_692),
.B(n_578),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_690),
.B(n_646),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_705),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_686),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_666),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_729),
.B(n_646),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_705),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_664),
.A2(n_719),
.B1(n_684),
.B2(n_722),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_717),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_681),
.Y(n_777)
);

OAI322xp33_ASAP7_75t_L g778 ( 
.A1(n_717),
.A2(n_585),
.A3(n_579),
.B1(n_583),
.B2(n_581),
.C1(n_647),
.C2(n_594),
.Y(n_778)
);

NOR3x1_ASAP7_75t_L g779 ( 
.A(n_709),
.B(n_514),
.C(n_502),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_705),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_724),
.Y(n_781)
);

OAI211xp5_ASAP7_75t_L g782 ( 
.A1(n_729),
.A2(n_585),
.B(n_581),
.C(n_583),
.Y(n_782)
);

AOI33xp33_ASAP7_75t_L g783 ( 
.A1(n_671),
.A2(n_583),
.A3(n_24),
.B1(n_25),
.B2(n_27),
.B3(n_18),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_706),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_706),
.Y(n_785)
);

OAI33xp33_ASAP7_75t_L g786 ( 
.A1(n_686),
.A2(n_647),
.A3(n_594),
.B1(n_635),
.B2(n_559),
.B3(n_558),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_714),
.Y(n_787)
);

NAND4xp75_ASAP7_75t_L g788 ( 
.A(n_684),
.B(n_549),
.C(n_555),
.D(n_573),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_714),
.Y(n_789)
);

NAND5xp2_ASAP7_75t_L g790 ( 
.A(n_693),
.B(n_508),
.C(n_453),
.D(n_358),
.E(n_517),
.Y(n_790)
);

O2A1O1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_664),
.A2(n_549),
.B(n_563),
.C(n_602),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_663),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_663),
.Y(n_793)
);

OAI222xp33_ASAP7_75t_L g794 ( 
.A1(n_664),
.A2(n_562),
.B1(n_599),
.B2(n_544),
.C1(n_559),
.C2(n_558),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_695),
.B(n_458),
.Y(n_795)
);

OA222x2_ASAP7_75t_L g796 ( 
.A1(n_664),
.A2(n_554),
.B1(n_602),
.B2(n_603),
.C1(n_599),
.C2(n_564),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_776),
.B(n_694),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_731),
.A2(n_664),
.B1(n_719),
.B2(n_671),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_743),
.Y(n_799)
);

XOR2xp5_ASAP7_75t_L g800 ( 
.A(n_763),
.B(n_717),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_792),
.Y(n_801)
);

XOR2x2_ASAP7_75t_L g802 ( 
.A(n_795),
.B(n_671),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_731),
.A2(n_673),
.B(n_709),
.Y(n_803)
);

AOI21xp33_ASAP7_75t_L g804 ( 
.A1(n_791),
.A2(n_675),
.B(n_726),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_795),
.B(n_458),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_793),
.Y(n_806)
);

XNOR2x1_ASAP7_75t_L g807 ( 
.A(n_744),
.B(n_695),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_771),
.B(n_670),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_751),
.Y(n_809)
);

OAI21xp33_ASAP7_75t_L g810 ( 
.A1(n_761),
.A2(n_693),
.B(n_703),
.Y(n_810)
);

AOI21xp33_ASAP7_75t_SL g811 ( 
.A1(n_756),
.A2(n_673),
.B(n_667),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_787),
.B(n_670),
.Y(n_812)
);

OAI32xp33_ASAP7_75t_L g813 ( 
.A1(n_754),
.A2(n_694),
.A3(n_665),
.B1(n_685),
.B2(n_726),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_758),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_745),
.A2(n_667),
.B(n_670),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_768),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_762),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_789),
.B(n_695),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_L g819 ( 
.A(n_737),
.B(n_675),
.C(n_700),
.Y(n_819)
);

NAND3xp33_ASAP7_75t_L g820 ( 
.A(n_745),
.B(n_718),
.C(n_726),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_736),
.B(n_694),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_750),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_744),
.A2(n_698),
.B(n_696),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_L g824 ( 
.A(n_752),
.B(n_718),
.C(n_700),
.Y(n_824)
);

OAI21xp33_ASAP7_75t_L g825 ( 
.A1(n_783),
.A2(n_693),
.B(n_703),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_740),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_742),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_756),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_786),
.A2(n_722),
.B1(n_723),
.B2(n_667),
.Y(n_829)
);

OAI21xp5_ASAP7_75t_L g830 ( 
.A1(n_783),
.A2(n_755),
.B(n_752),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_755),
.A2(n_722),
.B(n_723),
.C(n_728),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_786),
.A2(n_723),
.B1(n_703),
.B2(n_728),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_766),
.A2(n_775),
.B1(n_753),
.B2(n_760),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_SL g834 ( 
.A1(n_778),
.A2(n_698),
.B(n_696),
.Y(n_834)
);

CKINVDCx16_ASAP7_75t_R g835 ( 
.A(n_739),
.Y(n_835)
);

AOI211xp5_ASAP7_75t_SL g836 ( 
.A1(n_772),
.A2(n_696),
.B(n_698),
.C(n_677),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_769),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_734),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_SL g839 ( 
.A(n_794),
.B(n_562),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_735),
.Y(n_840)
);

OAI211xp5_ASAP7_75t_SL g841 ( 
.A1(n_785),
.A2(n_685),
.B(n_665),
.C(n_700),
.Y(n_841)
);

OAI21xp33_ASAP7_75t_SL g842 ( 
.A1(n_772),
.A2(n_687),
.B(n_691),
.Y(n_842)
);

OAI21xp33_ASAP7_75t_L g843 ( 
.A1(n_764),
.A2(n_728),
.B(n_704),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_741),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_749),
.Y(n_845)
);

XOR2x2_ASAP7_75t_L g846 ( 
.A(n_788),
.B(n_724),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_782),
.A2(n_677),
.B1(n_725),
.B2(n_712),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_773),
.A2(n_677),
.B1(n_725),
.B2(n_712),
.Y(n_848)
);

XNOR2xp5_ASAP7_75t_L g849 ( 
.A(n_767),
.B(n_725),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_759),
.Y(n_850)
);

INVx1_ASAP7_75t_SL g851 ( 
.A(n_765),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_830),
.B(n_851),
.Y(n_852)
);

XNOR2x2_ASAP7_75t_L g853 ( 
.A(n_830),
.B(n_796),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_851),
.B(n_746),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_835),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_SL g856 ( 
.A1(n_836),
.A2(n_803),
.B(n_834),
.C(n_805),
.Y(n_856)
);

AND2x2_ASAP7_75t_SL g857 ( 
.A(n_839),
.B(n_779),
.Y(n_857)
);

OAI211xp5_ASAP7_75t_L g858 ( 
.A1(n_798),
.A2(n_748),
.B(n_784),
.C(n_785),
.Y(n_858)
);

OAI321xp33_ASAP7_75t_L g859 ( 
.A1(n_820),
.A2(n_784),
.A3(n_790),
.B1(n_747),
.B2(n_699),
.C(n_683),
.Y(n_859)
);

XNOR2xp5_ASAP7_75t_L g860 ( 
.A(n_800),
.B(n_807),
.Y(n_860)
);

OAI22xp33_ASAP7_75t_SL g861 ( 
.A1(n_815),
.A2(n_753),
.B1(n_732),
.B2(n_777),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_815),
.A2(n_732),
.B1(n_733),
.B2(n_780),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_831),
.A2(n_781),
.B1(n_767),
.B2(n_687),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_801),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_797),
.Y(n_865)
);

OAI21xp33_ASAP7_75t_SL g866 ( 
.A1(n_847),
.A2(n_691),
.B(n_687),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_806),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_819),
.B(n_825),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_839),
.A2(n_738),
.B1(n_774),
.B2(n_770),
.Y(n_869)
);

CKINVDCx16_ASAP7_75t_R g870 ( 
.A(n_833),
.Y(n_870)
);

OAI322xp33_ASAP7_75t_L g871 ( 
.A1(n_832),
.A2(n_699),
.A3(n_683),
.B1(n_680),
.B2(n_727),
.C1(n_678),
.C2(n_674),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_799),
.Y(n_872)
);

OAI31xp33_ASAP7_75t_L g873 ( 
.A1(n_804),
.A2(n_794),
.A3(n_777),
.B(n_757),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_850),
.B(n_691),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_844),
.Y(n_875)
);

O2A1O1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_813),
.A2(n_563),
.B(n_727),
.C(n_680),
.Y(n_876)
);

OAI221xp5_ASAP7_75t_L g877 ( 
.A1(n_846),
.A2(n_697),
.B1(n_668),
.B2(n_716),
.C(n_674),
.Y(n_877)
);

OAI311xp33_ASAP7_75t_L g878 ( 
.A1(n_842),
.A2(n_708),
.A3(n_704),
.B1(n_678),
.C1(n_668),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_837),
.B(n_697),
.Y(n_879)
);

NOR3xp33_ASAP7_75t_SL g880 ( 
.A(n_841),
.B(n_716),
.C(n_535),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_809),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_802),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_SL g883 ( 
.A1(n_836),
.A2(n_704),
.B(n_708),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_814),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_828),
.B(n_708),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_822),
.B(n_682),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_829),
.A2(n_682),
.B1(n_712),
.B2(n_715),
.Y(n_887)
);

OAI322xp33_ASAP7_75t_L g888 ( 
.A1(n_822),
.A2(n_721),
.A3(n_720),
.B1(n_681),
.B2(n_689),
.C1(n_710),
.C2(n_711),
.Y(n_888)
);

OAI22xp33_ASAP7_75t_L g889 ( 
.A1(n_848),
.A2(n_564),
.B1(n_562),
.B2(n_554),
.Y(n_889)
);

OR2x2_ASAP7_75t_L g890 ( 
.A(n_818),
.B(n_682),
.Y(n_890)
);

NOR2xp67_ASAP7_75t_SL g891 ( 
.A(n_824),
.B(n_447),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_810),
.A2(n_696),
.B(n_698),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_SL g893 ( 
.A1(n_811),
.A2(n_696),
.B(n_698),
.Y(n_893)
);

OAI21xp33_ASAP7_75t_SL g894 ( 
.A1(n_808),
.A2(n_715),
.B(n_720),
.Y(n_894)
);

OAI31xp33_ASAP7_75t_L g895 ( 
.A1(n_826),
.A2(n_715),
.A3(n_720),
.B(n_721),
.Y(n_895)
);

OAI211xp5_ASAP7_75t_L g896 ( 
.A1(n_843),
.A2(n_535),
.B(n_517),
.C(n_602),
.Y(n_896)
);

OAI21xp33_ASAP7_75t_L g897 ( 
.A1(n_827),
.A2(n_721),
.B(n_720),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_817),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_838),
.B(n_840),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_855),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_882),
.B(n_812),
.Y(n_901)
);

OAI221xp5_ASAP7_75t_L g902 ( 
.A1(n_860),
.A2(n_873),
.B1(n_868),
.B2(n_852),
.C(n_877),
.Y(n_902)
);

NAND3xp33_ASAP7_75t_L g903 ( 
.A(n_876),
.B(n_823),
.C(n_816),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_856),
.A2(n_849),
.B(n_845),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_865),
.B(n_821),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_899),
.Y(n_906)
);

AOI221xp5_ASAP7_75t_L g907 ( 
.A1(n_876),
.A2(n_721),
.B1(n_710),
.B2(n_681),
.C(n_689),
.Y(n_907)
);

NAND4xp75_ASAP7_75t_L g908 ( 
.A(n_857),
.B(n_710),
.C(n_689),
.D(n_681),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_859),
.A2(n_858),
.B(n_854),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_878),
.A2(n_563),
.B(n_710),
.C(n_689),
.Y(n_910)
);

AOI211xp5_ASAP7_75t_L g911 ( 
.A1(n_877),
.A2(n_641),
.B(n_564),
.C(n_626),
.Y(n_911)
);

OAI21xp33_ASAP7_75t_L g912 ( 
.A1(n_858),
.A2(n_711),
.B(n_707),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_872),
.B(n_711),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_SL g914 ( 
.A(n_870),
.B(n_861),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_880),
.B(n_564),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_864),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_885),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_867),
.B(n_707),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_881),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_880),
.B(n_564),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_884),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_898),
.B(n_707),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_875),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_874),
.B(n_563),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_853),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_879),
.Y(n_926)
);

NOR2x1_ASAP7_75t_L g927 ( 
.A(n_883),
.B(n_408),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_887),
.A2(n_564),
.B1(n_554),
.B2(n_653),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_890),
.B(n_641),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_896),
.B(n_564),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_886),
.Y(n_931)
);

OR2x2_ASAP7_75t_L g932 ( 
.A(n_863),
.B(n_563),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_871),
.B(n_600),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_866),
.B(n_600),
.Y(n_934)
);

OAI21xp33_ASAP7_75t_L g935 ( 
.A1(n_862),
.A2(n_547),
.B(n_541),
.Y(n_935)
);

NOR3x1_ASAP7_75t_L g936 ( 
.A(n_893),
.B(n_378),
.C(n_379),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_900),
.Y(n_937)
);

NAND3xp33_ASAP7_75t_L g938 ( 
.A(n_909),
.B(n_891),
.C(n_895),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_916),
.Y(n_939)
);

NOR3xp33_ASAP7_75t_L g940 ( 
.A(n_902),
.B(n_896),
.C(n_894),
.Y(n_940)
);

NOR3xp33_ASAP7_75t_SL g941 ( 
.A(n_904),
.B(n_892),
.C(n_889),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_900),
.B(n_897),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_914),
.A2(n_888),
.B(n_892),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_916),
.Y(n_944)
);

NAND3xp33_ASAP7_75t_L g945 ( 
.A(n_925),
.B(n_910),
.C(n_901),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_917),
.B(n_869),
.Y(n_946)
);

OAI211xp5_ASAP7_75t_L g947 ( 
.A1(n_910),
.A2(n_429),
.B(n_408),
.C(n_600),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_906),
.B(n_641),
.Y(n_948)
);

AOI211x1_ASAP7_75t_L g949 ( 
.A1(n_903),
.A2(n_572),
.B(n_544),
.C(n_558),
.Y(n_949)
);

NAND2x1_ASAP7_75t_L g950 ( 
.A(n_927),
.B(n_626),
.Y(n_950)
);

OAI22xp33_ASAP7_75t_L g951 ( 
.A1(n_933),
.A2(n_564),
.B1(n_602),
.B2(n_603),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_901),
.A2(n_547),
.B1(n_541),
.B2(n_641),
.Y(n_952)
);

AOI211x1_ASAP7_75t_L g953 ( 
.A1(n_912),
.A2(n_559),
.B(n_544),
.C(n_542),
.Y(n_953)
);

AO22x1_ASAP7_75t_L g954 ( 
.A1(n_933),
.A2(n_626),
.B1(n_429),
.B2(n_408),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_923),
.Y(n_955)
);

AOI31xp33_ASAP7_75t_L g956 ( 
.A1(n_919),
.A2(n_603),
.A3(n_547),
.B(n_541),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_907),
.A2(n_547),
.B(n_541),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_908),
.A2(n_603),
.B(n_541),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_911),
.A2(n_541),
.B(n_547),
.C(n_429),
.Y(n_959)
);

OAI21xp33_ASAP7_75t_L g960 ( 
.A1(n_931),
.A2(n_547),
.B(n_643),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_921),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_926),
.B(n_643),
.Y(n_962)
);

XOR2xp5_ASAP7_75t_L g963 ( 
.A(n_905),
.B(n_447),
.Y(n_963)
);

NOR3xp33_ASAP7_75t_L g964 ( 
.A(n_924),
.B(n_398),
.C(n_439),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_SL g965 ( 
.A1(n_934),
.A2(n_932),
.B(n_920),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_913),
.B(n_643),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_929),
.Y(n_967)
);

NOR3x1_ASAP7_75t_L g968 ( 
.A(n_915),
.B(n_378),
.C(n_379),
.Y(n_968)
);

NOR3xp33_ASAP7_75t_L g969 ( 
.A(n_934),
.B(n_379),
.C(n_378),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_918),
.B(n_572),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_922),
.Y(n_971)
);

NOR3xp33_ASAP7_75t_L g972 ( 
.A(n_935),
.B(n_390),
.C(n_374),
.Y(n_972)
);

AOI211xp5_ASAP7_75t_L g973 ( 
.A1(n_930),
.A2(n_600),
.B(n_447),
.C(n_398),
.Y(n_973)
);

AOI221xp5_ASAP7_75t_L g974 ( 
.A1(n_945),
.A2(n_928),
.B1(n_936),
.B2(n_542),
.C(n_572),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_937),
.B(n_542),
.Y(n_975)
);

OAI221xp5_ASAP7_75t_L g976 ( 
.A1(n_940),
.A2(n_573),
.B1(n_409),
.B2(n_574),
.C(n_575),
.Y(n_976)
);

AOI221xp5_ASAP7_75t_L g977 ( 
.A1(n_943),
.A2(n_573),
.B1(n_575),
.B2(n_574),
.C(n_560),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_955),
.B(n_600),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_942),
.B(n_600),
.Y(n_979)
);

NAND3xp33_ASAP7_75t_L g980 ( 
.A(n_941),
.B(n_447),
.C(n_600),
.Y(n_980)
);

NOR3xp33_ASAP7_75t_SL g981 ( 
.A(n_938),
.B(n_447),
.C(n_600),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_963),
.Y(n_982)
);

AOI32xp33_ASAP7_75t_L g983 ( 
.A1(n_951),
.A2(n_452),
.A3(n_427),
.B1(n_371),
.B2(n_398),
.Y(n_983)
);

OAI211xp5_ASAP7_75t_SL g984 ( 
.A1(n_939),
.A2(n_398),
.B(n_437),
.C(n_439),
.Y(n_984)
);

AOI221xp5_ASAP7_75t_L g985 ( 
.A1(n_949),
.A2(n_560),
.B1(n_575),
.B2(n_574),
.C(n_571),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_971),
.B(n_600),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_944),
.A2(n_439),
.B(n_437),
.C(n_387),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_961),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_947),
.A2(n_390),
.B(n_371),
.C(n_346),
.Y(n_989)
);

AOI221xp5_ASAP7_75t_L g990 ( 
.A1(n_971),
.A2(n_575),
.B1(n_574),
.B2(n_571),
.C(n_570),
.Y(n_990)
);

AOI321xp33_ASAP7_75t_L g991 ( 
.A1(n_946),
.A2(n_452),
.A3(n_570),
.B1(n_567),
.B2(n_566),
.C(n_560),
.Y(n_991)
);

NOR2x1_ASAP7_75t_R g992 ( 
.A(n_967),
.B(n_447),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_950),
.A2(n_437),
.B1(n_439),
.B2(n_460),
.Y(n_993)
);

OAI221xp5_ASAP7_75t_SL g994 ( 
.A1(n_965),
.A2(n_460),
.B1(n_432),
.B2(n_437),
.C(n_566),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_962),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_972),
.A2(n_387),
.B(n_432),
.C(n_374),
.Y(n_996)
);

OAI211xp5_ASAP7_75t_SL g997 ( 
.A1(n_973),
.A2(n_374),
.B(n_338),
.C(n_567),
.Y(n_997)
);

AOI221xp5_ASAP7_75t_L g998 ( 
.A1(n_953),
.A2(n_571),
.B1(n_570),
.B2(n_567),
.C(n_566),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_948),
.B(n_380),
.Y(n_999)
);

OAI21xp33_ASAP7_75t_SL g1000 ( 
.A1(n_956),
.A2(n_571),
.B(n_570),
.Y(n_1000)
);

OAI221xp5_ASAP7_75t_L g1001 ( 
.A1(n_972),
.A2(n_567),
.B1(n_566),
.B2(n_560),
.C(n_364),
.Y(n_1001)
);

OAI221xp5_ASAP7_75t_SL g1002 ( 
.A1(n_959),
.A2(n_338),
.B1(n_470),
.B2(n_459),
.C(n_445),
.Y(n_1002)
);

OAI221xp5_ASAP7_75t_L g1003 ( 
.A1(n_952),
.A2(n_364),
.B1(n_380),
.B2(n_450),
.C(n_365),
.Y(n_1003)
);

OAI222xp33_ASAP7_75t_L g1004 ( 
.A1(n_957),
.A2(n_375),
.B1(n_365),
.B2(n_464),
.C1(n_411),
.C2(n_410),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_969),
.A2(n_387),
.B1(n_347),
.B2(n_350),
.Y(n_1005)
);

OAI222xp33_ASAP7_75t_L g1006 ( 
.A1(n_954),
.A2(n_966),
.B1(n_970),
.B2(n_968),
.C1(n_969),
.C2(n_958),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_988),
.B(n_964),
.Y(n_1007)
);

AOI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_977),
.A2(n_960),
.B1(n_347),
.B2(n_350),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_978),
.B(n_361),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_995),
.Y(n_1010)
);

NOR2x1_ASAP7_75t_L g1011 ( 
.A(n_980),
.B(n_982),
.Y(n_1011)
);

OA22x2_ASAP7_75t_L g1012 ( 
.A1(n_975),
.A2(n_367),
.B1(n_333),
.B2(n_375),
.Y(n_1012)
);

NOR2x1_ASAP7_75t_L g1013 ( 
.A(n_986),
.B(n_337),
.Y(n_1013)
);

AO22x2_ASAP7_75t_L g1014 ( 
.A1(n_993),
.A2(n_361),
.B1(n_360),
.B2(n_445),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_976),
.Y(n_1015)
);

NOR2x1_ASAP7_75t_L g1016 ( 
.A(n_1006),
.B(n_337),
.Y(n_1016)
);

NOR2x1_ASAP7_75t_L g1017 ( 
.A(n_1006),
.B(n_337),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_987),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_999),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_992),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1001),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_974),
.A2(n_347),
.B1(n_350),
.B2(n_380),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_981),
.A2(n_380),
.B1(n_332),
.B2(n_334),
.Y(n_1023)
);

OR2x2_ASAP7_75t_L g1024 ( 
.A(n_979),
.B(n_337),
.Y(n_1024)
);

NOR2x1_ASAP7_75t_L g1025 ( 
.A(n_984),
.B(n_330),
.Y(n_1025)
);

AOI31xp33_ASAP7_75t_L g1026 ( 
.A1(n_1000),
.A2(n_361),
.A3(n_392),
.B(n_380),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_994),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_989),
.B(n_361),
.Y(n_1028)
);

NOR2x1_ASAP7_75t_L g1029 ( 
.A(n_997),
.B(n_330),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_1003),
.A2(n_347),
.B1(n_350),
.B2(n_367),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_996),
.Y(n_1031)
);

AOI221xp5_ASAP7_75t_L g1032 ( 
.A1(n_1018),
.A2(n_1004),
.B1(n_983),
.B2(n_1002),
.C(n_990),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_1010),
.B(n_1005),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1011),
.B(n_1020),
.Y(n_1034)
);

OAI221xp5_ASAP7_75t_L g1035 ( 
.A1(n_1016),
.A2(n_1017),
.B1(n_1031),
.B2(n_1022),
.C(n_1027),
.Y(n_1035)
);

NAND4xp75_ASAP7_75t_L g1036 ( 
.A(n_1021),
.B(n_1019),
.C(n_1015),
.D(n_1007),
.Y(n_1036)
);

AND4x1_ASAP7_75t_L g1037 ( 
.A(n_1025),
.B(n_985),
.C(n_998),
.D(n_991),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1029),
.B(n_330),
.Y(n_1038)
);

NAND3xp33_ASAP7_75t_L g1039 ( 
.A(n_1030),
.B(n_330),
.C(n_332),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_1009),
.B(n_361),
.Y(n_1040)
);

XOR2xp5_ASAP7_75t_SL g1041 ( 
.A(n_1013),
.B(n_392),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_1024),
.Y(n_1042)
);

NOR3xp33_ASAP7_75t_L g1043 ( 
.A(n_1026),
.B(n_1028),
.C(n_1008),
.Y(n_1043)
);

AOI222xp33_ASAP7_75t_L g1044 ( 
.A1(n_1014),
.A2(n_367),
.B1(n_360),
.B2(n_464),
.C1(n_445),
.C2(n_431),
.Y(n_1044)
);

NAND4xp75_ASAP7_75t_L g1045 ( 
.A(n_1014),
.B(n_392),
.C(n_464),
.D(n_402),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_1023),
.Y(n_1046)
);

NAND4xp75_ASAP7_75t_L g1047 ( 
.A(n_1012),
.B(n_392),
.C(n_459),
.D(n_401),
.Y(n_1047)
);

NAND4xp75_ASAP7_75t_L g1048 ( 
.A(n_1011),
.B(n_392),
.C(n_459),
.D(n_401),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1010),
.B(n_330),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_1011),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_1010),
.B(n_333),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_1034),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_1050),
.A2(n_333),
.B(n_376),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1049),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_1036),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_1046),
.B(n_332),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_1033),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_1042),
.Y(n_1058)
);

NAND2x1p5_ASAP7_75t_L g1059 ( 
.A(n_1040),
.B(n_332),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_1048),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1051),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_1040),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_1041),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1047),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1035),
.Y(n_1065)
);

XOR2xp5_ASAP7_75t_L g1066 ( 
.A(n_1045),
.B(n_332),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_R g1067 ( 
.A(n_1038),
.B(n_392),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1057),
.Y(n_1068)
);

XNOR2xp5_ASAP7_75t_L g1069 ( 
.A(n_1055),
.B(n_1043),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1052),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1052),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_1052),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1058),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_1055),
.Y(n_1074)
);

OA22x2_ASAP7_75t_L g1075 ( 
.A1(n_1058),
.A2(n_1032),
.B1(n_1037),
.B2(n_1039),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_1056),
.Y(n_1076)
);

OAI31xp33_ASAP7_75t_L g1077 ( 
.A1(n_1074),
.A2(n_1065),
.A3(n_1064),
.B(n_1060),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_1070),
.B(n_1054),
.Y(n_1078)
);

OAI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_1075),
.A2(n_1063),
.B1(n_1061),
.B2(n_1062),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1072),
.B(n_1056),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1068),
.B(n_1062),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1071),
.Y(n_1082)
);

OA22x2_ASAP7_75t_L g1083 ( 
.A1(n_1069),
.A2(n_1066),
.B1(n_1053),
.B2(n_1062),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1073),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_SL g1085 ( 
.A1(n_1084),
.A2(n_1076),
.B1(n_1075),
.B2(n_1059),
.Y(n_1085)
);

OR3x1_ASAP7_75t_L g1086 ( 
.A(n_1082),
.B(n_1067),
.C(n_1053),
.Y(n_1086)
);

OAI22x1_ASAP7_75t_L g1087 ( 
.A1(n_1078),
.A2(n_1059),
.B1(n_1037),
.B2(n_1044),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1080),
.A2(n_1081),
.B1(n_1079),
.B2(n_1083),
.Y(n_1088)
);

INVxp67_ASAP7_75t_L g1089 ( 
.A(n_1077),
.Y(n_1089)
);

AOI22x1_ASAP7_75t_L g1090 ( 
.A1(n_1084),
.A2(n_332),
.B1(n_334),
.B2(n_359),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1085),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1089),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1086),
.A2(n_334),
.B1(n_359),
.B2(n_358),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_R g1094 ( 
.A1(n_1087),
.A2(n_402),
.B1(n_415),
.B2(n_411),
.Y(n_1094)
);

AOI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1091),
.A2(n_1088),
.B(n_1090),
.Y(n_1095)
);

INVxp67_ASAP7_75t_SL g1096 ( 
.A(n_1092),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1096),
.A2(n_1093),
.B1(n_1094),
.B2(n_334),
.Y(n_1097)
);

OR2x6_ASAP7_75t_L g1098 ( 
.A(n_1097),
.B(n_1095),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1098),
.A2(n_334),
.B1(n_359),
.B2(n_402),
.Y(n_1099)
);


endmodule