module real_jpeg_30599_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_215;
wire n_166;
wire n_176;
wire n_292;
wire n_221;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_11;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_205;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_297;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_244;
wire n_133;
wire n_216;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_0),
.Y(n_160)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_0),
.Y(n_188)
);

INVx3_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_1),
.A2(n_47),
.B1(n_84),
.B2(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_1),
.A2(n_47),
.B1(n_150),
.B2(n_153),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_1),
.B(n_20),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_1),
.B(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_1),
.B(n_263),
.C(n_266),
.Y(n_262)
);

NAND2xp67_ASAP7_75t_L g278 ( 
.A(n_1),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_1),
.B(n_285),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_3),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_3),
.Y(n_110)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_4),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_4),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_5),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_5),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_6),
.Y(n_140)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_8),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_8),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_9),
.A2(n_192),
.B1(n_193),
.B2(n_197),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_9),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_207),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_205),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp67_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_167),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_15),
.B(n_167),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_122),
.C(n_162),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_16),
.B(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_55),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_18),
.B(n_56),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

AO22x2_ASAP7_75t_L g169 ( 
.A1(n_19),
.A2(n_92),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_19),
.Y(n_171)
);

OAI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_33),
.B(n_46),
.Y(n_19)
);

OAI22x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.B1(n_28),
.B2(n_31),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_23),
.Y(n_128)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_27),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_27),
.Y(n_145)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2x1_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_40),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_39),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_44),
.Y(n_136)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B(n_51),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_47),
.A2(n_116),
.B(n_120),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_47),
.B(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_51),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_55),
.B(n_214),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_91),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_56),
.B(n_92),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_56),
.A2(n_184),
.B1(n_203),
.B2(n_204),
.Y(n_183)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_56),
.Y(n_203)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_56),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_56),
.A2(n_147),
.B1(n_148),
.B2(n_203),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_56),
.A2(n_203),
.B1(n_257),
.B2(n_258),
.Y(n_288)
);

OA21x2_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_72),
.B(n_88),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_58),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B1(n_66),
.B2(n_68),
.Y(n_58)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_59),
.Y(n_161)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_59),
.Y(n_198)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_61),
.Y(n_196)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_65),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22x1_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_77),
.B1(n_81),
.B2(n_84),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_80),
.Y(n_222)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_87),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_92),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_92),
.B(n_171),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_102),
.B(n_115),
.Y(n_92)
);

NOR2x1p5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_103),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_93),
.Y(n_253)
);

OAI22x1_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_99),
.B2(n_101),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_96),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_96),
.Y(n_231)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_107),
.B1(n_111),
.B2(n_112),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_119),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_120),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_122),
.B(n_163),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_147),
.Y(n_122)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_132),
.B(n_137),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx4f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_141),
.B(n_146),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx2_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_164),
.C(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_147),
.B(n_173),
.Y(n_172)
);

NAND2x1p5_ASAP7_75t_L g242 ( 
.A(n_147),
.B(n_215),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_147),
.A2(n_148),
.B1(n_165),
.B2(n_166),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_147),
.B(n_243),
.C(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_147),
.B(n_288),
.Y(n_287)
);

CKINVDCx11_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_148),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_148),
.B(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_148),
.B(n_284),
.Y(n_283)
);

OR2x6_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_155),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_149),
.A2(n_185),
.B1(n_191),
.B2(n_199),
.Y(n_184)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx4f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_161),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_160),
.Y(n_279)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_SL g211 ( 
.A1(n_164),
.A2(n_212),
.B(n_214),
.C(n_238),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_164),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_176),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_168)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_182),
.B2(n_183),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_178),
.Y(n_177)
);

AND3x1_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.C(n_181),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_208),
.Y(n_207)
);

OAI21x1_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_293),
.B(n_297),
.Y(n_208)
);

AOI21x1_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_248),
.B(n_292),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_239),
.Y(n_210)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_211),
.B(n_239),
.Y(n_292)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_213),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_213),
.B(n_242),
.C(n_244),
.Y(n_294)
);

OAI21x1_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_219),
.B(n_227),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_232),
.B(n_236),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_244),
.B1(n_245),
.B2(n_247),
.Y(n_239)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI21x1_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_254),
.B(n_291),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_251),
.Y(n_291)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_274),
.B(n_289),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_270),
.Y(n_255)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_256),
.Y(n_290)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_287),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_283),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NOR2x1_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_295),
.Y(n_297)
);


endmodule