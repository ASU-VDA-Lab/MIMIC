module fake_ariane_1436_n_1681 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1681);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1681;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_SL g147 ( 
.A(n_82),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_16),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_93),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_13),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_60),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_90),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_80),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_3),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_35),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_14),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_6),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_101),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_7),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_105),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_37),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_54),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_57),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_136),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_48),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_143),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_95),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_62),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_51),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_32),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_137),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_32),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_142),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_8),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_20),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_5),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_140),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_1),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_8),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_85),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_28),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_117),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_33),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_42),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_49),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_38),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_0),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_134),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_44),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_106),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_14),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_42),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_103),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_73),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_99),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_78),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_118),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_50),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_114),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_35),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_121),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_41),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_107),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_38),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_65),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_97),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_75),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_46),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_144),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_91),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_145),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_89),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_130),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_92),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_124),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_64),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_36),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_26),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_71),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_81),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_109),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_131),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_52),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_25),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_2),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_47),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_17),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_31),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_25),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_98),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_146),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_58),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_7),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_40),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_59),
.Y(n_239)
);

BUFx2_ASAP7_75t_SL g240 ( 
.A(n_129),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_3),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_138),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_45),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_110),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_63),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_133),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_67),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_126),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_10),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_19),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_122),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_113),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_44),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_19),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_120),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_102),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_104),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_45),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_128),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_46),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_56),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_83),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_31),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_43),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_55),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_1),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_127),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_18),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_69),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_43),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_135),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_112),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_72),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_141),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_111),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_37),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_70),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_53),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_26),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_39),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_33),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_41),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_16),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_34),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_4),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_40),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_88),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_0),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_34),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_123),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_6),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_115),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_116),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_76),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_100),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_189),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_237),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_260),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_266),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_260),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_260),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_282),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_282),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_282),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_291),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_276),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_284),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_284),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_190),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_148),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_284),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_274),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_207),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_160),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_171),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_150),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_207),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_191),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_227),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_160),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_166),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_166),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_245),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_204),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_204),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_161),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_172),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_155),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_174),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_227),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_245),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_177),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_178),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_179),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_181),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_182),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_273),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_273),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_171),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_275),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_184),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_275),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_267),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_211),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_186),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_246),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_195),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_154),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_208),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_221),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_222),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_190),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_231),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_156),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_233),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_187),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_243),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_162),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_250),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_190),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_264),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_263),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_279),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_281),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_358),
.A2(n_232),
.B1(n_268),
.B2(n_228),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_165),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_319),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_319),
.Y(n_374)
);

INVx6_ASAP7_75t_L g375 ( 
.A(n_309),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_330),
.B(n_176),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_308),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_354),
.B(n_197),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_312),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_323),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_334),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_323),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_325),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_320),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_308),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_321),
.B(n_247),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_325),
.Y(n_387)
);

OAI21x1_ASAP7_75t_L g388 ( 
.A1(n_312),
.A2(n_202),
.B(n_199),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_R g389 ( 
.A(n_318),
.B(n_149),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_312),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_364),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_321),
.B(n_217),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_296),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_296),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_336),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_345),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_336),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_343),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_298),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_298),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_326),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_345),
.B(n_360),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_220),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_343),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_299),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_344),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_299),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_316),
.B(n_267),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_311),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_315),
.A2(n_268),
.B1(n_232),
.B2(n_254),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_300),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_331),
.B(n_267),
.Y(n_413)
);

NAND2xp33_ASAP7_75t_L g414 ( 
.A(n_322),
.B(n_292),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_327),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_328),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_346),
.Y(n_417)
);

BUFx8_ASAP7_75t_L g418 ( 
.A(n_349),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_346),
.B(n_223),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_300),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_301),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_348),
.B(n_200),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_301),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_302),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_351),
.B(n_289),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_348),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_302),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_304),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_304),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_305),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_305),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_329),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_351),
.B(n_264),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_306),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_306),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_335),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_337),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_307),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_307),
.B(n_244),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_324),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_427),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_390),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_390),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_411),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_408),
.Y(n_445)
);

BUFx6f_ASAP7_75t_SL g446 ( 
.A(n_422),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_418),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_350),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_390),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_411),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_396),
.Y(n_451)
);

BUFx4f_ASAP7_75t_L g452 ( 
.A(n_390),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_411),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_433),
.B(n_332),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_427),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_411),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_428),
.Y(n_458)
);

INVx8_ASAP7_75t_L g459 ( 
.A(n_433),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_413),
.B(n_352),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_408),
.B(n_338),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_408),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_411),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_429),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_410),
.B(n_297),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_429),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_390),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_390),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_430),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_421),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_433),
.A2(n_261),
.B1(n_228),
.B2(n_288),
.Y(n_471)
);

AO21x2_ASAP7_75t_L g472 ( 
.A1(n_388),
.A2(n_256),
.B(n_248),
.Y(n_472)
);

BUFx8_ASAP7_75t_SL g473 ( 
.A(n_384),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_418),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_396),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_390),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_396),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_421),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_SL g479 ( 
.A1(n_410),
.A2(n_280),
.B1(n_288),
.B2(n_254),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_430),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_421),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_390),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_402),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_391),
.B(n_372),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_421),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_421),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_423),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_379),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_423),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_376),
.B(n_339),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_423),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_423),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_423),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_434),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_377),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_434),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_434),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_434),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_389),
.B(n_341),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_434),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_379),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_379),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_409),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_379),
.Y(n_504)
);

NAND3xp33_ASAP7_75t_L g505 ( 
.A(n_414),
.B(n_194),
.C(n_342),
.Y(n_505)
);

CKINVDCx6p67_ASAP7_75t_R g506 ( 
.A(n_409),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_401),
.Y(n_507)
);

NAND3xp33_ASAP7_75t_L g508 ( 
.A(n_414),
.B(n_362),
.C(n_347),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_379),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_422),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_394),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_389),
.B(n_367),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_377),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_373),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_377),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_391),
.B(n_340),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_394),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_381),
.B(n_366),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_375),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_376),
.B(n_164),
.Y(n_520)
);

INVx5_ASAP7_75t_L g521 ( 
.A(n_377),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_372),
.B(n_357),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_373),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_399),
.Y(n_524)
);

AOI21x1_ASAP7_75t_L g525 ( 
.A1(n_388),
.A2(n_313),
.B(n_310),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_399),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_399),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_422),
.Y(n_528)
);

OR2x6_ASAP7_75t_L g529 ( 
.A(n_375),
.B(n_391),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_436),
.B(n_164),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_381),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_436),
.B(n_167),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_374),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_374),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_380),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_380),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_377),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_400),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_400),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_382),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_R g541 ( 
.A(n_418),
.B(n_303),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_382),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_377),
.Y(n_543)
);

INVxp33_ASAP7_75t_SL g544 ( 
.A(n_432),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_377),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_L g546 ( 
.A(n_425),
.B(n_167),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_375),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_383),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_418),
.B(n_168),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_400),
.Y(n_550)
);

INVx8_ASAP7_75t_L g551 ( 
.A(n_422),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_383),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_377),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_405),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_393),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_387),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_405),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_387),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_405),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_375),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_395),
.Y(n_561)
);

OR2x6_ASAP7_75t_L g562 ( 
.A(n_375),
.B(n_353),
.Y(n_562)
);

OAI22xp33_ASAP7_75t_L g563 ( 
.A1(n_371),
.A2(n_280),
.B1(n_258),
.B2(n_261),
.Y(n_563)
);

BUFx10_ASAP7_75t_L g564 ( 
.A(n_375),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_372),
.B(n_310),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_420),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_418),
.B(n_168),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_420),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_378),
.B(n_169),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_378),
.A2(n_264),
.B1(n_157),
.B2(n_155),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_386),
.B(n_333),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_420),
.Y(n_572)
);

BUFx10_ASAP7_75t_L g573 ( 
.A(n_386),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_378),
.B(n_353),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_393),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_424),
.Y(n_576)
);

NAND2xp33_ASAP7_75t_SL g577 ( 
.A(n_425),
.B(n_157),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_424),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_424),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_431),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_395),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_397),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_431),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_425),
.A2(n_158),
.B1(n_159),
.B2(n_163),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_397),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_422),
.Y(n_586)
);

INVxp33_ASAP7_75t_L g587 ( 
.A(n_371),
.Y(n_587)
);

AOI21x1_ASAP7_75t_L g588 ( 
.A1(n_388),
.A2(n_314),
.B(n_317),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_573),
.B(n_169),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_479),
.A2(n_398),
.B1(n_412),
.B2(n_406),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_573),
.B(n_170),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_483),
.B(n_571),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_503),
.B(n_402),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g594 ( 
.A(n_558),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_503),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_574),
.B(n_392),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_573),
.B(n_170),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_558),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_558),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_518),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_441),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_445),
.B(n_392),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_501),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_518),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_459),
.Y(n_605)
);

AND2x6_ASAP7_75t_SL g606 ( 
.A(n_544),
.B(n_355),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_501),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_484),
.A2(n_454),
.B1(n_516),
.B2(n_514),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_445),
.B(n_403),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_573),
.B(n_239),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_L g611 ( 
.A(n_459),
.B(n_239),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_490),
.B(n_403),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_461),
.B(n_462),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_531),
.B(n_159),
.C(n_158),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_462),
.B(n_398),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_459),
.B(n_404),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_459),
.B(n_404),
.Y(n_617)
);

NAND3xp33_ASAP7_75t_L g618 ( 
.A(n_546),
.B(n_238),
.C(n_163),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_473),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_L g620 ( 
.A(n_459),
.B(n_287),
.Y(n_620)
);

O2A1O1Ixp33_ASAP7_75t_L g621 ( 
.A1(n_520),
.A2(n_523),
.B(n_533),
.C(n_514),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_454),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_510),
.B(n_528),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_510),
.B(n_406),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_506),
.B(n_355),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_440),
.B(n_412),
.Y(n_626)
);

BUFx8_ASAP7_75t_L g627 ( 
.A(n_446),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_510),
.B(n_417),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_510),
.B(n_417),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_L g630 ( 
.A1(n_471),
.A2(n_584),
.B1(n_587),
.B2(n_529),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_528),
.B(n_426),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_528),
.B(n_586),
.Y(n_632)
);

NOR3xp33_ASAP7_75t_L g633 ( 
.A(n_448),
.B(n_286),
.C(n_238),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_451),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_455),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_511),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_451),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_564),
.B(n_426),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_528),
.A2(n_286),
.B1(n_253),
.B2(n_192),
.Y(n_639)
);

AO22x2_ASAP7_75t_L g640 ( 
.A1(n_465),
.A2(n_356),
.B1(n_369),
.B2(n_368),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_455),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_586),
.B(n_484),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_460),
.B(n_419),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_586),
.B(n_419),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_522),
.B(n_508),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_586),
.B(n_516),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g647 ( 
.A1(n_481),
.A2(n_439),
.B(n_262),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_517),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_507),
.Y(n_649)
);

O2A1O1Ixp5_ASAP7_75t_L g650 ( 
.A1(n_523),
.A2(n_439),
.B(n_438),
.C(n_435),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_505),
.A2(n_200),
.B1(n_271),
.B2(n_240),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_508),
.B(n_206),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_564),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_551),
.B(n_533),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_551),
.B(n_534),
.Y(n_655)
);

OR2x6_ASAP7_75t_L g656 ( 
.A(n_529),
.B(n_356),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_551),
.B(n_147),
.Y(n_657)
);

OAI22xp33_ASAP7_75t_L g658 ( 
.A1(n_471),
.A2(n_359),
.B1(n_370),
.B2(n_369),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_505),
.A2(n_212),
.B1(n_270),
.B2(n_283),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_456),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_551),
.B(n_229),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_517),
.Y(n_662)
);

BUFx5_ASAP7_75t_L g663 ( 
.A(n_564),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_551),
.B(n_255),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_534),
.B(n_431),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_529),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_535),
.B(n_435),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_535),
.B(n_435),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_536),
.B(n_438),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_536),
.B(n_438),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_519),
.B(n_241),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_456),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_540),
.B(n_359),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_458),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_458),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_451),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_541),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_540),
.B(n_361),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_547),
.B(n_249),
.Y(n_679)
);

NOR2xp67_ASAP7_75t_L g680 ( 
.A(n_447),
.B(n_361),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_584),
.B(n_363),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_512),
.B(n_363),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_542),
.B(n_365),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_547),
.B(n_285),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_465),
.B(n_384),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_542),
.B(n_365),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_562),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_446),
.A2(n_259),
.B1(n_272),
.B2(n_277),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_548),
.A2(n_385),
.B1(n_368),
.B2(n_370),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_548),
.B(n_151),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_552),
.B(n_556),
.Y(n_691)
);

NOR2xp67_ASAP7_75t_L g692 ( 
.A(n_447),
.B(n_385),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_SL g693 ( 
.A1(n_570),
.A2(n_437),
.B1(n_416),
.B2(n_415),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_552),
.A2(n_385),
.B1(n_278),
.B2(n_290),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_560),
.B(n_152),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_464),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_529),
.B(n_415),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_446),
.A2(n_293),
.B1(n_224),
.B2(n_219),
.Y(n_698)
);

O2A1O1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_556),
.A2(n_313),
.B(n_314),
.C(n_317),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_464),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_466),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_466),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_524),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_526),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_529),
.A2(n_153),
.B1(n_173),
.B2(n_175),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_562),
.Y(n_706)
);

O2A1O1Ixp5_ASAP7_75t_L g707 ( 
.A1(n_561),
.A2(n_393),
.B(n_407),
.C(n_292),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_474),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_562),
.Y(n_709)
);

OR2x6_ASAP7_75t_L g710 ( 
.A(n_562),
.B(n_437),
.Y(n_710)
);

AO22x2_ASAP7_75t_L g711 ( 
.A1(n_563),
.A2(n_416),
.B1(n_4),
.B2(n_5),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_476),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_569),
.B(n_2),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_562),
.A2(n_218),
.B1(n_183),
.B2(n_295),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_530),
.B(n_9),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_581),
.A2(n_407),
.B1(n_393),
.B2(n_226),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_475),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_582),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_499),
.B(n_180),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_526),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_469),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_527),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_577),
.A2(n_225),
.B1(n_188),
.B2(n_294),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_532),
.B(n_185),
.Y(n_724)
);

NAND2x1_ASAP7_75t_L g725 ( 
.A(n_443),
.B(n_407),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_469),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_475),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_549),
.A2(n_193),
.B1(n_196),
.B2(n_198),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_582),
.B(n_234),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_527),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_476),
.B(n_292),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_567),
.A2(n_230),
.B1(n_203),
.B2(n_205),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_480),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_585),
.B(n_236),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_538),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_488),
.B(n_11),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_475),
.Y(n_737)
);

AO22x2_ASAP7_75t_L g738 ( 
.A1(n_565),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_585),
.A2(n_235),
.B1(n_209),
.B2(n_269),
.Y(n_739)
);

A2O1A1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_481),
.A2(n_407),
.B(n_393),
.C(n_265),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_474),
.B(n_12),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_488),
.B(n_201),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_477),
.B(n_407),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_480),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_538),
.A2(n_407),
.B1(n_393),
.B2(n_226),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_539),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_488),
.B(n_15),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_502),
.Y(n_748)
);

NOR3xp33_ASAP7_75t_L g749 ( 
.A(n_595),
.B(n_502),
.C(n_504),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_612),
.B(n_504),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_601),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_649),
.Y(n_752)
);

INVx8_ASAP7_75t_L g753 ( 
.A(n_656),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_612),
.B(n_509),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_656),
.B(n_477),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_643),
.B(n_509),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_643),
.B(n_444),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_600),
.B(n_477),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_592),
.B(n_444),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_596),
.B(n_450),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_666),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_645),
.B(n_450),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_656),
.B(n_666),
.Y(n_763)
);

INVxp33_ASAP7_75t_L g764 ( 
.A(n_625),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_635),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_645),
.B(n_646),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_666),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_604),
.B(n_593),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_SL g769 ( 
.A1(n_640),
.A2(n_711),
.B1(n_693),
.B2(n_681),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_666),
.B(n_476),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_712),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_622),
.A2(n_489),
.B1(n_498),
.B2(n_497),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_619),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_743),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_608),
.B(n_453),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_622),
.B(n_453),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_641),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_R g778 ( 
.A(n_708),
.B(n_468),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_608),
.B(n_457),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_687),
.B(n_476),
.Y(n_780)
);

NAND2xp33_ASAP7_75t_L g781 ( 
.A(n_663),
.B(n_482),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_660),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_626),
.B(n_457),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_672),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_697),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_613),
.B(n_605),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_697),
.Y(n_787)
);

CKINVDCx8_ASAP7_75t_R g788 ( 
.A(n_606),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_674),
.B(n_675),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_613),
.A2(n_652),
.B1(n_630),
.B2(n_715),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_696),
.B(n_463),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_640),
.B(n_470),
.Y(n_792)
);

BUFx4f_ASAP7_75t_L g793 ( 
.A(n_710),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_650),
.A2(n_496),
.B(n_500),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_685),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_700),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_743),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_701),
.B(n_470),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_702),
.B(n_721),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_636),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_726),
.B(n_478),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_627),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_709),
.B(n_478),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_733),
.B(n_485),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_744),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_652),
.A2(n_489),
.B1(n_485),
.B2(n_491),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_627),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_648),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_748),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_677),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_634),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_710),
.Y(n_812)
);

AND3x1_ASAP7_75t_SL g813 ( 
.A(n_658),
.B(n_496),
.C(n_494),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_594),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_737),
.A2(n_452),
.B(n_487),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_712),
.Y(n_816)
);

AND2x6_ASAP7_75t_L g817 ( 
.A(n_634),
.B(n_486),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_706),
.B(n_491),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_594),
.B(n_492),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_590),
.B(n_492),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_712),
.Y(n_821)
);

INVxp67_ASAP7_75t_L g822 ( 
.A(n_682),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_673),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_678),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_642),
.B(n_443),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_662),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_644),
.B(n_497),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_741),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_691),
.B(n_498),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_663),
.B(n_482),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_715),
.A2(n_493),
.B1(n_500),
.B2(n_494),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_737),
.B(n_486),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_590),
.A2(n_658),
.B1(n_711),
.B2(n_640),
.Y(n_833)
);

INVx2_ASAP7_75t_SL g834 ( 
.A(n_719),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_711),
.B(n_633),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_680),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_712),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_683),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_686),
.Y(n_839)
);

NOR2x1p5_ASAP7_75t_L g840 ( 
.A(n_614),
.B(n_442),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_615),
.B(n_487),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_609),
.B(n_618),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_602),
.B(n_443),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_650),
.A2(n_493),
.B(n_588),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_713),
.A2(n_566),
.B1(n_583),
.B2(n_580),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_665),
.Y(n_846)
);

AND2x6_ASAP7_75t_L g847 ( 
.A(n_637),
.B(n_442),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_713),
.A2(n_633),
.B1(n_598),
.B2(n_599),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_667),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_663),
.B(n_482),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_668),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_736),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_615),
.B(n_539),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_727),
.B(n_550),
.Y(n_854)
);

INVx3_ASAP7_75t_L g855 ( 
.A(n_637),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_639),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_669),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_670),
.Y(n_858)
);

AND2x6_ASAP7_75t_SL g859 ( 
.A(n_736),
.B(n_17),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_663),
.B(n_482),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_703),
.Y(n_861)
);

OAI221xp5_ASAP7_75t_L g862 ( 
.A1(n_659),
.A2(n_550),
.B1(n_583),
.B2(n_580),
.C(n_579),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_704),
.A2(n_568),
.B1(n_579),
.B2(n_578),
.Y(n_863)
);

NAND2x1p5_ASAP7_75t_L g864 ( 
.A(n_676),
.B(n_449),
.Y(n_864)
);

BUFx8_ASAP7_75t_L g865 ( 
.A(n_603),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_676),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_727),
.B(n_554),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_720),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_589),
.B(n_449),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_591),
.B(n_449),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_597),
.B(n_449),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_607),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_689),
.B(n_554),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_722),
.Y(n_874)
);

NOR3xp33_ASAP7_75t_SL g875 ( 
.A(n_724),
.B(n_216),
.C(n_257),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_717),
.B(n_557),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_730),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_663),
.B(n_482),
.Y(n_878)
);

INVx4_ASAP7_75t_L g879 ( 
.A(n_717),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_725),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_735),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_621),
.B(n_557),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_654),
.B(n_559),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_671),
.Y(n_884)
);

NOR3xp33_ASAP7_75t_SL g885 ( 
.A(n_610),
.B(n_214),
.C(n_252),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_657),
.A2(n_575),
.B1(n_467),
.B2(n_468),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_664),
.B(n_452),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_746),
.A2(n_572),
.B1(n_578),
.B2(n_576),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_624),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_653),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_653),
.B(n_705),
.Y(n_891)
);

OAI21xp33_ASAP7_75t_SL g892 ( 
.A1(n_655),
.A2(n_628),
.B(n_631),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_629),
.B(n_568),
.Y(n_893)
);

OR2x6_ASAP7_75t_L g894 ( 
.A(n_692),
.B(n_566),
.Y(n_894)
);

INVx4_ASAP7_75t_L g895 ( 
.A(n_738),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_623),
.B(n_576),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_632),
.B(n_467),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_731),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_616),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_738),
.A2(n_559),
.B1(n_572),
.B2(n_472),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_651),
.A2(n_575),
.B1(n_467),
.B2(n_468),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_617),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_731),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_647),
.B(n_442),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_699),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_714),
.B(n_467),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_661),
.A2(n_611),
.B1(n_620),
.B2(n_739),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_689),
.B(n_442),
.Y(n_908)
);

INVx5_ASAP7_75t_L g909 ( 
.A(n_638),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_707),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_747),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_738),
.A2(n_472),
.B1(n_575),
.B2(n_555),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_688),
.B(n_515),
.Y(n_913)
);

NOR2xp67_ASAP7_75t_L g914 ( 
.A(n_698),
.B(n_723),
.Y(n_914)
);

NAND2x1p5_ASAP7_75t_L g915 ( 
.A(n_638),
.B(n_543),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_707),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_679),
.B(n_495),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_690),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_747),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_742),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_684),
.B(n_495),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_728),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_729),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_732),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_734),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_751),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_810),
.Y(n_927)
);

NAND3xp33_ASAP7_75t_L g928 ( 
.A(n_790),
.B(n_718),
.C(n_695),
.Y(n_928)
);

AO32x1_ASAP7_75t_L g929 ( 
.A1(n_895),
.A2(n_740),
.A3(n_472),
.B1(n_588),
.B2(n_525),
.Y(n_929)
);

INVx4_ASAP7_75t_L g930 ( 
.A(n_753),
.Y(n_930)
);

O2A1O1Ixp5_ASAP7_75t_L g931 ( 
.A1(n_891),
.A2(n_515),
.B(n_495),
.C(n_543),
.Y(n_931)
);

NOR2x1_ASAP7_75t_R g932 ( 
.A(n_773),
.B(n_215),
.Y(n_932)
);

AO21x2_ASAP7_75t_L g933 ( 
.A1(n_882),
.A2(n_525),
.B(n_694),
.Y(n_933)
);

BUFx12f_ASAP7_75t_L g934 ( 
.A(n_802),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_768),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_764),
.B(n_822),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_766),
.A2(n_515),
.B(n_495),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_795),
.B(n_785),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_756),
.B(n_694),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_756),
.A2(n_716),
.B1(n_745),
.B2(n_513),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_828),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_781),
.A2(n_513),
.B(n_553),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_787),
.B(n_716),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_SL g944 ( 
.A(n_924),
.B(n_210),
.C(n_213),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_844),
.A2(n_537),
.B(n_553),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_750),
.A2(n_545),
.B(n_555),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_833),
.A2(n_745),
.B1(n_545),
.B2(n_555),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_793),
.B(n_393),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_765),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_SL g950 ( 
.A1(n_788),
.A2(n_242),
.B1(n_251),
.B2(n_226),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_750),
.A2(n_555),
.B(n_521),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_754),
.A2(n_757),
.B(n_783),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_793),
.B(n_393),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_800),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_767),
.Y(n_955)
);

OR2x6_ASAP7_75t_L g956 ( 
.A(n_753),
.B(n_226),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_808),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_777),
.Y(n_958)
);

INVx3_ASAP7_75t_SL g959 ( 
.A(n_807),
.Y(n_959)
);

BUFx12f_ASAP7_75t_L g960 ( 
.A(n_865),
.Y(n_960)
);

NOR3xp33_ASAP7_75t_L g961 ( 
.A(n_914),
.B(n_18),
.C(n_20),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_754),
.B(n_757),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_826),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_R g964 ( 
.A(n_812),
.B(n_79),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_782),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_783),
.A2(n_521),
.B(n_77),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_753),
.B(n_521),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_823),
.B(n_824),
.Y(n_968)
);

OAI22xp33_ASAP7_75t_L g969 ( 
.A1(n_895),
.A2(n_521),
.B1(n_22),
.B2(n_23),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_784),
.Y(n_970)
);

OAI22x1_ASAP7_75t_L g971 ( 
.A1(n_835),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_789),
.A2(n_21),
.B1(n_24),
.B2(n_27),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_842),
.A2(n_292),
.B(n_28),
.C(n_29),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_769),
.B(n_792),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_752),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_796),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_755),
.B(n_292),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_758),
.B(n_292),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_805),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_838),
.B(n_292),
.Y(n_980)
);

NOR2xp67_ASAP7_75t_SL g981 ( 
.A(n_890),
.B(n_27),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_SL g982 ( 
.A1(n_922),
.A2(n_30),
.B1(n_36),
.B2(n_39),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_R g983 ( 
.A(n_865),
.B(n_761),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_771),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_778),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_816),
.Y(n_986)
);

INVx8_ASAP7_75t_L g987 ( 
.A(n_763),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_923),
.A2(n_61),
.B(n_66),
.C(n_68),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_763),
.B(n_918),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_761),
.B(n_74),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_809),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_SL g992 ( 
.A1(n_911),
.A2(n_84),
.B(n_86),
.C(n_87),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_874),
.Y(n_993)
);

O2A1O1Ixp5_ASAP7_75t_L g994 ( 
.A1(n_887),
.A2(n_94),
.B(n_96),
.C(n_108),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_877),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_881),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_834),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_892),
.A2(n_925),
.B(n_919),
.C(n_839),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_820),
.A2(n_797),
.B1(n_774),
.B2(n_861),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_852),
.A2(n_789),
.B(n_799),
.C(n_786),
.Y(n_1000)
);

BUFx12f_ASAP7_75t_L g1001 ( 
.A(n_859),
.Y(n_1001)
);

O2A1O1Ixp5_ASAP7_75t_L g1002 ( 
.A1(n_906),
.A2(n_871),
.B(n_870),
.C(n_869),
.Y(n_1002)
);

NOR3xp33_ASAP7_75t_SL g1003 ( 
.A(n_799),
.B(n_921),
.C(n_917),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_907),
.A2(n_841),
.B1(n_814),
.B2(n_760),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_872),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_836),
.B(n_884),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_868),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_846),
.B(n_849),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_776),
.B(n_803),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_818),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_920),
.B(n_774),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_759),
.A2(n_762),
.B(n_853),
.Y(n_1012)
);

OAI21xp33_ASAP7_75t_L g1013 ( 
.A1(n_889),
.A2(n_848),
.B(n_841),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_760),
.A2(n_853),
.B1(n_858),
.B2(n_857),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_851),
.B(n_762),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_749),
.A2(n_759),
.B(n_920),
.C(n_829),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_854),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_775),
.B(n_779),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_913),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_819),
.A2(n_832),
.B(n_829),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_791),
.Y(n_1021)
);

INVx11_ASAP7_75t_L g1022 ( 
.A(n_817),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_SL g1023 ( 
.A1(n_912),
.A2(n_913),
.B1(n_813),
.B2(n_909),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_775),
.B(n_779),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_819),
.A2(n_832),
.B(n_843),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_791),
.A2(n_804),
.B(n_798),
.C(n_801),
.Y(n_1026)
);

CKINVDCx10_ASAP7_75t_R g1027 ( 
.A(n_894),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_798),
.Y(n_1028)
);

NOR3xp33_ASAP7_75t_SL g1029 ( 
.A(n_794),
.B(n_844),
.C(n_804),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_902),
.B(n_899),
.Y(n_1030)
);

OR2x6_ASAP7_75t_L g1031 ( 
.A(n_894),
.B(n_902),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_893),
.A2(n_827),
.B(n_825),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_854),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_873),
.B(n_899),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_893),
.A2(n_896),
.B(n_883),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_771),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_771),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_840),
.B(n_885),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_905),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_909),
.B(n_879),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_831),
.A2(n_806),
.B(n_904),
.C(n_772),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_821),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_909),
.B(n_879),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_875),
.Y(n_1044)
);

BUFx12f_ASAP7_75t_SL g1045 ( 
.A(n_894),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_908),
.A2(n_867),
.B1(n_883),
.B2(n_896),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_908),
.A2(n_909),
.B1(n_901),
.B2(n_876),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_811),
.B(n_866),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_897),
.B(n_866),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_815),
.A2(n_878),
.B(n_860),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_897),
.B(n_855),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_882),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_941),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_973),
.A2(n_855),
.B(n_780),
.C(n_770),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_960),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_927),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_926),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_1025),
.A2(n_850),
.B(n_830),
.Y(n_1058)
);

OAI22x1_ASAP7_75t_L g1059 ( 
.A1(n_1039),
.A2(n_915),
.B1(n_898),
.B2(n_916),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_1003),
.A2(n_886),
.B(n_862),
.C(n_845),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1032),
.A2(n_876),
.B(n_910),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_1013),
.A2(n_903),
.B(n_900),
.C(n_890),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_1035),
.A2(n_915),
.B(n_864),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1041),
.A2(n_863),
.B(n_888),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_998),
.A2(n_864),
.B(n_847),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_SL g1066 ( 
.A1(n_1000),
.A2(n_1015),
.B(n_962),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_952),
.A2(n_821),
.B(n_837),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_1020),
.A2(n_837),
.B(n_880),
.Y(n_1068)
);

BUFx4_ASAP7_75t_SL g1069 ( 
.A(n_997),
.Y(n_1069)
);

AO31x2_ASAP7_75t_L g1070 ( 
.A1(n_1046),
.A2(n_903),
.A3(n_817),
.B(n_847),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1004),
.A2(n_847),
.B(n_817),
.Y(n_1071)
);

OAI22x1_ASAP7_75t_L g1072 ( 
.A1(n_1044),
.A2(n_880),
.B1(n_903),
.B2(n_1019),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_928),
.A2(n_1016),
.B(n_939),
.C(n_1026),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1008),
.B(n_1009),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_966),
.A2(n_937),
.B(n_931),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_946),
.A2(n_1047),
.B(n_951),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1008),
.B(n_935),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1014),
.A2(n_1002),
.B(n_939),
.Y(n_1078)
);

NOR4xp25_ASAP7_75t_L g1079 ( 
.A(n_972),
.B(n_969),
.C(n_1014),
.D(n_1015),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_1047),
.A2(n_945),
.B(n_942),
.Y(n_1080)
);

OA21x2_ASAP7_75t_L g1081 ( 
.A1(n_1029),
.A2(n_945),
.B(n_1024),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_949),
.Y(n_1082)
);

BUFx2_ASAP7_75t_R g1083 ( 
.A(n_959),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_1022),
.A2(n_1033),
.B1(n_1023),
.B2(n_1021),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_1046),
.A2(n_1024),
.A3(n_1018),
.B(n_1052),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_975),
.B(n_1011),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_983),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1028),
.A2(n_985),
.B1(n_1049),
.B2(n_1051),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_958),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_967),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_965),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_970),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_976),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_938),
.B(n_989),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1049),
.A2(n_1051),
.B1(n_982),
.B2(n_1010),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_961),
.A2(n_1038),
.B(n_1034),
.C(n_1017),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_979),
.Y(n_1097)
);

AOI21x1_ASAP7_75t_SL g1098 ( 
.A1(n_980),
.A2(n_990),
.B(n_1034),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_991),
.Y(n_1099)
);

AOI221xp5_ASAP7_75t_L g1100 ( 
.A1(n_971),
.A2(n_972),
.B1(n_944),
.B2(n_950),
.C(n_1006),
.Y(n_1100)
);

BUFx4_ASAP7_75t_SL g1101 ( 
.A(n_956),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_936),
.B(n_974),
.Y(n_1102)
);

NOR2x1_ASAP7_75t_SL g1103 ( 
.A(n_967),
.B(n_1031),
.Y(n_1103)
);

AOI221xp5_ASAP7_75t_SL g1104 ( 
.A1(n_1048),
.A2(n_940),
.B1(n_999),
.B2(n_988),
.C(n_977),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_993),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_948),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_940),
.A2(n_1043),
.B(n_1040),
.Y(n_1107)
);

OR2x6_ASAP7_75t_L g1108 ( 
.A(n_987),
.B(n_967),
.Y(n_1108)
);

AO21x2_ASAP7_75t_L g1109 ( 
.A1(n_933),
.A2(n_1030),
.B(n_995),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_933),
.A2(n_992),
.B(n_929),
.Y(n_1110)
);

OA21x2_ASAP7_75t_L g1111 ( 
.A1(n_994),
.A2(n_947),
.B(n_996),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1005),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_990),
.B(n_1036),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1001),
.B(n_943),
.Y(n_1114)
);

NOR2xp67_ASAP7_75t_L g1115 ( 
.A(n_1042),
.B(n_986),
.Y(n_1115)
);

OAI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_981),
.A2(n_964),
.B(n_956),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_1031),
.B(n_953),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1007),
.B(n_963),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_1027),
.B(n_932),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_954),
.B(n_957),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1037),
.A2(n_955),
.B(n_929),
.Y(n_1121)
);

AOI221x1_ASAP7_75t_L g1122 ( 
.A1(n_1042),
.A2(n_984),
.B1(n_1036),
.B2(n_1045),
.C(n_934),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_984),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_987),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1009),
.B(n_768),
.Y(n_1125)
);

AO32x2_ASAP7_75t_L g1126 ( 
.A1(n_1046),
.A2(n_895),
.A3(n_1004),
.B1(n_1023),
.B2(n_1014),
.Y(n_1126)
);

OR2x6_ASAP7_75t_L g1127 ( 
.A(n_987),
.B(n_753),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1009),
.B(n_768),
.Y(n_1128)
);

INVx4_ASAP7_75t_L g1129 ( 
.A(n_1022),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_938),
.Y(n_1130)
);

AO32x2_ASAP7_75t_L g1131 ( 
.A1(n_1046),
.A2(n_895),
.A3(n_1004),
.B1(n_1023),
.B2(n_1014),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_927),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_926),
.Y(n_1133)
);

NAND2x1p5_ASAP7_75t_L g1134 ( 
.A(n_930),
.B(n_773),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_968),
.B(n_600),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1009),
.B(n_768),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_927),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_927),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1050),
.A2(n_1035),
.B(n_1012),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1014),
.B(n_790),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_973),
.B(n_790),
.C(n_961),
.Y(n_1141)
);

OR2x2_ASAP7_75t_L g1142 ( 
.A(n_938),
.B(n_795),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_941),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_968),
.B(n_600),
.Y(n_1144)
);

AO32x2_ASAP7_75t_L g1145 ( 
.A1(n_1046),
.A2(n_895),
.A3(n_1004),
.B1(n_1023),
.B2(n_1014),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1009),
.B(n_768),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1050),
.A2(n_1035),
.B(n_1012),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_968),
.B(n_600),
.Y(n_1148)
);

AO22x2_ASAP7_75t_L g1149 ( 
.A1(n_974),
.A2(n_895),
.B1(n_835),
.B2(n_465),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1050),
.A2(n_1035),
.B(n_1012),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_973),
.A2(n_490),
.B(n_856),
.C(n_961),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1039),
.A2(n_790),
.B(n_592),
.Y(n_1152)
);

NOR2xp67_ASAP7_75t_L g1153 ( 
.A(n_968),
.B(n_816),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_973),
.A2(n_490),
.B(n_856),
.C(n_961),
.Y(n_1154)
);

OAI21xp33_ASAP7_75t_L g1155 ( 
.A1(n_928),
.A2(n_790),
.B(n_612),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_968),
.B(n_600),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1050),
.A2(n_1035),
.B(n_1012),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_968),
.B(n_600),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_968),
.B(n_600),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1025),
.A2(n_1032),
.B(n_952),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_926),
.Y(n_1161)
);

INVx3_ASAP7_75t_SL g1162 ( 
.A(n_927),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1050),
.A2(n_1035),
.B(n_1012),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1022),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1003),
.A2(n_790),
.B(n_612),
.C(n_645),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1025),
.A2(n_1032),
.B(n_952),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_968),
.B(n_600),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_926),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1050),
.A2(n_1035),
.B(n_1012),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1050),
.A2(n_1035),
.B(n_1012),
.Y(n_1170)
);

AOI31xp67_ASAP7_75t_L g1171 ( 
.A1(n_978),
.A2(n_910),
.A3(n_916),
.B(n_887),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1025),
.A2(n_1032),
.B(n_952),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_968),
.B(n_600),
.Y(n_1173)
);

CKINVDCx11_ASAP7_75t_R g1174 ( 
.A(n_960),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1041),
.A2(n_790),
.B(n_1025),
.Y(n_1175)
);

AND2x6_ASAP7_75t_L g1176 ( 
.A(n_990),
.B(n_666),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1057),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1134),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1076),
.A2(n_1147),
.B(n_1139),
.Y(n_1179)
);

INVx5_ASAP7_75t_L g1180 ( 
.A(n_1176),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1082),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1075),
.A2(n_1157),
.B(n_1150),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1163),
.A2(n_1170),
.B(n_1169),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1089),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_1110),
.A2(n_1166),
.B(n_1160),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_1069),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1155),
.A2(n_1165),
.B(n_1140),
.C(n_1175),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1091),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1164),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1058),
.A2(n_1172),
.B(n_1061),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_1109),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1092),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1063),
.A2(n_1068),
.B(n_1121),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1093),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1053),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1080),
.A2(n_1098),
.B(n_1067),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1149),
.A2(n_1084),
.B1(n_1141),
.B2(n_1095),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1097),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1149),
.A2(n_1155),
.B1(n_1141),
.B2(n_1100),
.Y(n_1199)
);

OA21x2_ASAP7_75t_L g1200 ( 
.A1(n_1078),
.A2(n_1073),
.B(n_1104),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1074),
.B(n_1135),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1144),
.B(n_1148),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1099),
.Y(n_1203)
);

AOI332xp33_ASAP7_75t_L g1204 ( 
.A1(n_1133),
.A2(n_1168),
.A3(n_1161),
.B1(n_1125),
.B2(n_1128),
.B3(n_1146),
.C1(n_1136),
.C2(n_1077),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1085),
.Y(n_1205)
);

NAND3xp33_ASAP7_75t_L g1206 ( 
.A(n_1151),
.B(n_1154),
.C(n_1096),
.Y(n_1206)
);

OR2x6_ASAP7_75t_L g1207 ( 
.A(n_1108),
.B(n_1072),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_SL g1208 ( 
.A1(n_1066),
.A2(n_1152),
.B(n_1071),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1105),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1143),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1107),
.A2(n_1065),
.B(n_1064),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1112),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1085),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1114),
.B(n_1086),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1118),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1120),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_SL g1217 ( 
.A1(n_1102),
.A2(n_1064),
.B1(n_1176),
.B2(n_1131),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1054),
.A2(n_1081),
.B(n_1111),
.Y(n_1218)
);

NAND2x1p5_ASAP7_75t_L g1219 ( 
.A(n_1090),
.B(n_1113),
.Y(n_1219)
);

OR2x2_ASAP7_75t_L g1220 ( 
.A(n_1094),
.B(n_1130),
.Y(n_1220)
);

INVxp67_ASAP7_75t_L g1221 ( 
.A(n_1088),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1117),
.B(n_1103),
.Y(n_1222)
);

CKINVDCx16_ASAP7_75t_R g1223 ( 
.A(n_1055),
.Y(n_1223)
);

OAI222xp33_ASAP7_75t_L g1224 ( 
.A1(n_1130),
.A2(n_1106),
.B1(n_1173),
.B2(n_1159),
.C1(n_1158),
.C2(n_1167),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1153),
.A2(n_1171),
.B(n_1115),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1116),
.A2(n_1156),
.B1(n_1176),
.B2(n_1142),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1070),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1117),
.B(n_1108),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1162),
.B(n_1056),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1060),
.A2(n_1079),
.B(n_1062),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1122),
.A2(n_1164),
.B(n_1059),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1124),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1233)
);

AOI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1108),
.A2(n_1127),
.B(n_1079),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1106),
.Y(n_1235)
);

NAND2x1p5_ASAP7_75t_L g1236 ( 
.A(n_1124),
.B(n_1129),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1083),
.A2(n_1127),
.B1(n_1131),
.B2(n_1126),
.Y(n_1237)
);

AO21x2_ASAP7_75t_L g1238 ( 
.A1(n_1126),
.A2(n_1145),
.B(n_1131),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1124),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1070),
.Y(n_1240)
);

BUFx12f_ASAP7_75t_L g1241 ( 
.A(n_1174),
.Y(n_1241)
);

NAND2x1p5_ASAP7_75t_L g1242 ( 
.A(n_1123),
.B(n_1101),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1126),
.A2(n_1145),
.B(n_1123),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1137),
.B(n_1145),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1123),
.Y(n_1245)
);

BUFx4_ASAP7_75t_SL g1246 ( 
.A(n_1127),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1119),
.Y(n_1247)
);

OA21x2_ASAP7_75t_L g1248 ( 
.A1(n_1110),
.A2(n_1166),
.B(n_1160),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1057),
.Y(n_1249)
);

INVx4_ASAP7_75t_L g1250 ( 
.A(n_1056),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_SL g1251 ( 
.A1(n_1066),
.A2(n_1152),
.B(n_1175),
.Y(n_1251)
);

BUFx8_ASAP7_75t_L g1252 ( 
.A(n_1087),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1110),
.A2(n_1059),
.A3(n_1172),
.B(n_1166),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1057),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1109),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1174),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1057),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1174),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1076),
.A2(n_1147),
.B(n_1139),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1123),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1155),
.A2(n_790),
.B1(n_924),
.B2(n_1140),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1117),
.B(n_1090),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1057),
.Y(n_1263)
);

INVxp67_ASAP7_75t_SL g1264 ( 
.A(n_1140),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1117),
.B(n_1090),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1069),
.Y(n_1266)
);

NAND2x1p5_ASAP7_75t_L g1267 ( 
.A(n_1090),
.B(n_1010),
.Y(n_1267)
);

NOR2xp67_ASAP7_75t_R g1268 ( 
.A(n_1129),
.B(n_985),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1110),
.A2(n_1059),
.A3(n_1172),
.B(n_1166),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1110),
.A2(n_1166),
.B(n_1160),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1076),
.A2(n_1147),
.B(n_1139),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1057),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1076),
.A2(n_1147),
.B(n_1139),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1076),
.A2(n_1147),
.B(n_1139),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1123),
.Y(n_1275)
);

OA21x2_ASAP7_75t_L g1276 ( 
.A1(n_1110),
.A2(n_1166),
.B(n_1160),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1125),
.B(n_1128),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1165),
.A2(n_790),
.B1(n_1155),
.B2(n_1141),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1057),
.Y(n_1279)
);

XOR2xp5_ASAP7_75t_L g1280 ( 
.A(n_1083),
.B(n_384),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1110),
.A2(n_1166),
.B(n_1160),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1155),
.B(n_1140),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1165),
.A2(n_790),
.B1(n_1155),
.B2(n_1141),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1074),
.B(n_1135),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1149),
.A2(n_769),
.B1(n_833),
.B2(n_640),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1155),
.A2(n_1165),
.B(n_790),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1102),
.B(n_1094),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1155),
.A2(n_1165),
.B(n_790),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_SL g1289 ( 
.A1(n_1066),
.A2(n_1152),
.B(n_1175),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1057),
.Y(n_1290)
);

AND2x2_ASAP7_75t_SL g1291 ( 
.A(n_1200),
.B(n_1199),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1244),
.B(n_1277),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1177),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1241),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1220),
.B(n_1287),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1261),
.A2(n_1187),
.B1(n_1282),
.B2(n_1199),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_SL g1297 ( 
.A1(n_1187),
.A2(n_1283),
.B(n_1278),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_SL g1298 ( 
.A(n_1256),
.B(n_1258),
.Y(n_1298)
);

O2A1O1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1286),
.A2(n_1288),
.B(n_1282),
.C(n_1251),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1284),
.B(n_1202),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1214),
.B(n_1195),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_SL g1302 ( 
.A1(n_1237),
.A2(n_1200),
.B(n_1264),
.Y(n_1302)
);

OAI31xp33_ASAP7_75t_L g1303 ( 
.A1(n_1206),
.A2(n_1230),
.A3(n_1224),
.B(n_1285),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1289),
.A2(n_1208),
.B(n_1221),
.C(n_1264),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1235),
.B(n_1210),
.Y(n_1305)
);

AOI21x1_ASAP7_75t_SL g1306 ( 
.A1(n_1229),
.A2(n_1268),
.B(n_1233),
.Y(n_1306)
);

BUFx2_ASAP7_75t_R g1307 ( 
.A(n_1256),
.Y(n_1307)
);

INVx2_ASAP7_75t_SL g1308 ( 
.A(n_1252),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1221),
.B(n_1215),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1262),
.B(n_1265),
.Y(n_1310)
);

AOI221x1_ASAP7_75t_SL g1311 ( 
.A1(n_1247),
.A2(n_1194),
.B1(n_1212),
.B2(n_1209),
.C(n_1181),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1184),
.B(n_1188),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1197),
.A2(n_1204),
.B(n_1217),
.C(n_1211),
.Y(n_1313)
);

O2A1O1Ixp5_ASAP7_75t_L g1314 ( 
.A1(n_1234),
.A2(n_1205),
.B(n_1213),
.C(n_1227),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1192),
.B(n_1198),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1207),
.A2(n_1178),
.B(n_1242),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1203),
.B(n_1249),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1254),
.B(n_1257),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_R g1319 ( 
.A(n_1258),
.B(n_1180),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1228),
.B(n_1222),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1197),
.A2(n_1217),
.B1(n_1285),
.B2(n_1226),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1218),
.A2(n_1190),
.B(n_1182),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1226),
.A2(n_1189),
.B1(n_1242),
.B2(n_1236),
.Y(n_1323)
);

O2A1O1Ixp5_ASAP7_75t_L g1324 ( 
.A1(n_1240),
.A2(n_1224),
.B(n_1260),
.C(n_1275),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1263),
.B(n_1279),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1272),
.B(n_1290),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1216),
.B(n_1238),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1189),
.A2(n_1236),
.B1(n_1280),
.B2(n_1180),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_SL g1329 ( 
.A1(n_1207),
.A2(n_1238),
.B(n_1246),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1179),
.A2(n_1259),
.B(n_1274),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1180),
.A2(n_1223),
.B1(n_1186),
.B2(n_1266),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1245),
.B(n_1260),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1180),
.A2(n_1219),
.B1(n_1250),
.B2(n_1239),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1253),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1275),
.B(n_1243),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_SL g1336 ( 
.A1(n_1246),
.A2(n_1239),
.B(n_1232),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1252),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1191),
.A2(n_1267),
.B(n_1281),
.C(n_1276),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1232),
.B(n_1239),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1232),
.B(n_1239),
.Y(n_1340)
);

O2A1O1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1267),
.A2(n_1270),
.B(n_1281),
.C(n_1276),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1231),
.B(n_1225),
.Y(n_1342)
);

AOI211xp5_ASAP7_75t_L g1343 ( 
.A1(n_1196),
.A2(n_1193),
.B(n_1255),
.C(n_1179),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1252),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_SL g1345 ( 
.A1(n_1241),
.A2(n_1248),
.B1(n_1185),
.B2(n_1269),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_1185),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1259),
.B(n_1271),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1273),
.A2(n_790),
.B(n_1155),
.C(n_1230),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1183),
.B(n_1201),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1278),
.A2(n_1165),
.B(n_1283),
.C(n_1187),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1244),
.B(n_1277),
.Y(n_1351)
);

NOR2xp67_ASAP7_75t_L g1352 ( 
.A(n_1180),
.B(n_1250),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1244),
.B(n_1277),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1261),
.A2(n_1187),
.B1(n_790),
.B2(n_1282),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1244),
.B(n_1277),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1222),
.Y(n_1356)
);

O2A1O1Ixp5_ASAP7_75t_L g1357 ( 
.A1(n_1278),
.A2(n_1140),
.B(n_1175),
.C(n_1283),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1218),
.A2(n_1190),
.B(n_1182),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1218),
.A2(n_1190),
.B(n_1182),
.Y(n_1359)
);

O2A1O1Ixp5_ASAP7_75t_L g1360 ( 
.A1(n_1278),
.A2(n_1140),
.B(n_1175),
.C(n_1283),
.Y(n_1360)
);

O2A1O1Ixp5_ASAP7_75t_L g1361 ( 
.A1(n_1278),
.A2(n_1140),
.B(n_1175),
.C(n_1283),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1218),
.A2(n_1190),
.B(n_1182),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1244),
.B(n_1277),
.Y(n_1363)
);

OR2x6_ASAP7_75t_L g1364 ( 
.A(n_1207),
.B(n_1230),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1244),
.B(n_1277),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1187),
.A2(n_1165),
.B(n_1116),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1330),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1349),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1297),
.B(n_1354),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1293),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1327),
.B(n_1309),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1292),
.B(n_1351),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1353),
.B(n_1355),
.Y(n_1373)
);

CKINVDCx11_ASAP7_75t_R g1374 ( 
.A(n_1344),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1342),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1347),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1346),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1311),
.B(n_1325),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1363),
.B(n_1365),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1300),
.B(n_1291),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1314),
.A2(n_1348),
.B(n_1324),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1341),
.A2(n_1348),
.B(n_1338),
.Y(n_1382)
);

NAND2x1p5_ASAP7_75t_L g1383 ( 
.A(n_1291),
.B(n_1322),
.Y(n_1383)
);

BUFx2_ASAP7_75t_L g1384 ( 
.A(n_1335),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1312),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1315),
.B(n_1317),
.Y(n_1386)
);

AO21x2_ASAP7_75t_L g1387 ( 
.A1(n_1334),
.A2(n_1313),
.B(n_1302),
.Y(n_1387)
);

NAND3xp33_ASAP7_75t_L g1388 ( 
.A(n_1350),
.B(n_1296),
.C(n_1361),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1318),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1326),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1358),
.B(n_1359),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1358),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1358),
.Y(n_1393)
);

NOR2x1_ASAP7_75t_R g1394 ( 
.A(n_1294),
.B(n_1337),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1362),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1345),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1366),
.A2(n_1299),
.B1(n_1321),
.B2(n_1364),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1305),
.B(n_1295),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1343),
.B(n_1356),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1364),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1357),
.A2(n_1361),
.B(n_1360),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1304),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1301),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1368),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1374),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1374),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1368),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1368),
.B(n_1303),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1375),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1384),
.B(n_1320),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1367),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1375),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1371),
.B(n_1332),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1371),
.B(n_1329),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1371),
.B(n_1340),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1370),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1376),
.B(n_1372),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1370),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1370),
.Y(n_1419)
);

INVx5_ASAP7_75t_L g1420 ( 
.A(n_1400),
.Y(n_1420)
);

NAND3xp33_ASAP7_75t_L g1421 ( 
.A(n_1388),
.B(n_1323),
.C(n_1328),
.Y(n_1421)
);

INVx2_ASAP7_75t_R g1422 ( 
.A(n_1391),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1375),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1385),
.B(n_1339),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1399),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1398),
.B(n_1310),
.Y(n_1426)
);

OAI221xp5_ASAP7_75t_L g1427 ( 
.A1(n_1408),
.A2(n_1397),
.B1(n_1388),
.B2(n_1369),
.C(n_1396),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1425),
.B(n_1398),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1425),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1408),
.B(n_1378),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1416),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1425),
.B(n_1373),
.Y(n_1432)
);

AND2x6_ASAP7_75t_SL g1433 ( 
.A(n_1406),
.B(n_1307),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1413),
.B(n_1378),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1413),
.B(n_1385),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1425),
.B(n_1373),
.Y(n_1436)
);

OAI221xp5_ASAP7_75t_L g1437 ( 
.A1(n_1421),
.A2(n_1397),
.B1(n_1369),
.B2(n_1396),
.C(n_1380),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1406),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1421),
.A2(n_1387),
.B1(n_1396),
.B2(n_1401),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1415),
.B(n_1385),
.Y(n_1440)
);

NAND4xp25_ASAP7_75t_L g1441 ( 
.A(n_1421),
.B(n_1402),
.C(n_1409),
.D(n_1412),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1417),
.B(n_1373),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1404),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1416),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1415),
.B(n_1398),
.Y(n_1445)
);

INVxp67_ASAP7_75t_SL g1446 ( 
.A(n_1404),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1416),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1411),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1426),
.B(n_1403),
.Y(n_1449)
);

OAI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1414),
.A2(n_1380),
.B1(n_1377),
.B2(n_1383),
.C(n_1381),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1407),
.B(n_1402),
.C(n_1401),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1417),
.B(n_1379),
.Y(n_1452)
);

OA21x2_ASAP7_75t_L g1453 ( 
.A1(n_1411),
.A2(n_1392),
.B(n_1395),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1411),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1414),
.A2(n_1387),
.B1(n_1401),
.B2(n_1377),
.Y(n_1455)
);

OAI31xp33_ASAP7_75t_L g1456 ( 
.A1(n_1414),
.A2(n_1377),
.A3(n_1383),
.B(n_1399),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1423),
.B(n_1399),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1405),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1426),
.B(n_1403),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1407),
.B(n_1389),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1418),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1417),
.B(n_1379),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1418),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1418),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1426),
.A2(n_1401),
.B1(n_1383),
.B2(n_1352),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1410),
.B(n_1379),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1424),
.A2(n_1389),
.B1(n_1386),
.B2(n_1382),
.C(n_1387),
.Y(n_1467)
);

AOI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1424),
.A2(n_1389),
.B1(n_1382),
.B2(n_1387),
.C(n_1390),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1420),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1453),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1443),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1453),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1431),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1444),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1447),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1453),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1448),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1461),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_L g1479 ( 
.A(n_1430),
.B(n_1405),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1463),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1451),
.A2(n_1393),
.B(n_1392),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1454),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1464),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1438),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1460),
.Y(n_1485)
);

INVxp67_ASAP7_75t_SL g1486 ( 
.A(n_1439),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1428),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1445),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1429),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1438),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1445),
.Y(n_1491)
);

INVx4_ASAP7_75t_SL g1492 ( 
.A(n_1469),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1429),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1446),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1458),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1449),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1427),
.B(n_1394),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1434),
.B(n_1419),
.Y(n_1498)
);

INVx4_ASAP7_75t_SL g1499 ( 
.A(n_1469),
.Y(n_1499)
);

INVxp67_ASAP7_75t_SL g1500 ( 
.A(n_1455),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1428),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1449),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1432),
.B(n_1422),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1456),
.B(n_1409),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1504),
.B(n_1432),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1492),
.B(n_1457),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1504),
.B(n_1436),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1492),
.B(n_1436),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1484),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1484),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1478),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1486),
.B(n_1485),
.Y(n_1512)
);

NOR3xp33_ASAP7_75t_L g1513 ( 
.A(n_1486),
.B(n_1437),
.C(n_1441),
.Y(n_1513)
);

AND4x1_ASAP7_75t_L g1514 ( 
.A(n_1497),
.B(n_1298),
.C(n_1467),
.D(n_1468),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1498),
.B(n_1459),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1478),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1473),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1484),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1472),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1473),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1492),
.B(n_1457),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1490),
.B(n_1458),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1492),
.B(n_1457),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1490),
.B(n_1433),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1474),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1498),
.B(n_1459),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1474),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1485),
.B(n_1442),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1492),
.B(n_1442),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1484),
.B(n_1465),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1475),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1492),
.B(n_1469),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1488),
.B(n_1452),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1475),
.Y(n_1534)
);

NOR2x1_ASAP7_75t_L g1535 ( 
.A(n_1495),
.B(n_1331),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1480),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1488),
.B(n_1452),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1472),
.Y(n_1538)
);

INVxp67_ASAP7_75t_SL g1539 ( 
.A(n_1479),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1480),
.Y(n_1540)
);

OR2x6_ASAP7_75t_L g1541 ( 
.A(n_1472),
.B(n_1316),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1499),
.B(n_1462),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1499),
.B(n_1462),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1491),
.B(n_1435),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1491),
.B(n_1440),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1499),
.B(n_1466),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1519),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1512),
.B(n_1496),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1517),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1513),
.B(n_1496),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1517),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1532),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1546),
.B(n_1499),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1520),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1520),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1522),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1510),
.B(n_1502),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1525),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1525),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1527),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1527),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1509),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1531),
.Y(n_1563)
);

NAND2x1_ASAP7_75t_SL g1564 ( 
.A(n_1535),
.B(n_1497),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1531),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1534),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1510),
.B(n_1502),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1535),
.A2(n_1500),
.B(n_1514),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1534),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1536),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1536),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1506),
.B(n_1499),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1540),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1519),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1540),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1546),
.B(n_1499),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1544),
.B(n_1487),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1511),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1545),
.B(n_1487),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1511),
.Y(n_1580)
);

OAI31xp33_ASAP7_75t_L g1581 ( 
.A1(n_1505),
.A2(n_1500),
.A3(n_1450),
.B(n_1507),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1548),
.B(n_1515),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1562),
.B(n_1518),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1562),
.B(n_1539),
.Y(n_1584)
);

NOR2x1p5_ASAP7_75t_L g1585 ( 
.A(n_1552),
.B(n_1550),
.Y(n_1585)
);

AOI221xp5_ASAP7_75t_L g1586 ( 
.A1(n_1568),
.A2(n_1538),
.B1(n_1507),
.B2(n_1505),
.C(n_1530),
.Y(n_1586)
);

BUFx12f_ASAP7_75t_L g1587 ( 
.A(n_1572),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1549),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1553),
.B(n_1521),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1548),
.B(n_1515),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_SL g1591 ( 
.A1(n_1581),
.A2(n_1524),
.B1(n_1481),
.B2(n_1538),
.Y(n_1591)
);

INVx1_ASAP7_75t_SL g1592 ( 
.A(n_1564),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1564),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1572),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1552),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1551),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1554),
.Y(n_1597)
);

INVx3_ASAP7_75t_SL g1598 ( 
.A(n_1572),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1555),
.Y(n_1599)
);

INVx2_ASAP7_75t_SL g1600 ( 
.A(n_1552),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1547),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1557),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1553),
.B(n_1521),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1577),
.B(n_1533),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1567),
.Y(n_1605)
);

AND2x4_ASAP7_75t_SL g1606 ( 
.A(n_1576),
.B(n_1506),
.Y(n_1606)
);

INVx1_ASAP7_75t_SL g1607 ( 
.A(n_1598),
.Y(n_1607)
);

AOI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1592),
.A2(n_1556),
.B(n_1547),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1586),
.B(n_1532),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1591),
.A2(n_1574),
.B1(n_1541),
.B2(n_1387),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1598),
.A2(n_1508),
.B1(n_1543),
.B2(n_1542),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1602),
.B(n_1578),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1594),
.A2(n_1508),
.B1(n_1542),
.B2(n_1543),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1589),
.B(n_1576),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1582),
.B(n_1577),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1605),
.B(n_1580),
.Y(n_1616)
);

AOI22x1_ASAP7_75t_L g1617 ( 
.A1(n_1587),
.A2(n_1506),
.B1(n_1523),
.B2(n_1495),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1582),
.B(n_1579),
.Y(n_1618)
);

OAI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1593),
.A2(n_1541),
.B1(n_1574),
.B2(n_1579),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1590),
.B(n_1558),
.Y(n_1620)
);

OAI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1590),
.A2(n_1541),
.B1(n_1481),
.B2(n_1472),
.Y(n_1621)
);

A2O1A1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1585),
.A2(n_1479),
.B(n_1532),
.C(n_1476),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1601),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1584),
.B(n_1559),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1600),
.B(n_1560),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1607),
.B(n_1587),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1608),
.B(n_1600),
.Y(n_1627)
);

CKINVDCx16_ASAP7_75t_R g1628 ( 
.A(n_1614),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1615),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1610),
.A2(n_1601),
.B1(n_1596),
.B2(n_1597),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1608),
.B(n_1595),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1618),
.B(n_1606),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1620),
.B(n_1595),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1609),
.B(n_1589),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1623),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1612),
.B(n_1583),
.Y(n_1636)
);

AOI311xp33_ASAP7_75t_L g1637 ( 
.A1(n_1632),
.A2(n_1624),
.A3(n_1625),
.B(n_1616),
.C(n_1613),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1628),
.B(n_1617),
.Y(n_1638)
);

OAI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1630),
.A2(n_1631),
.B1(n_1622),
.B2(n_1627),
.C(n_1633),
.Y(n_1639)
);

NAND3xp33_ASAP7_75t_SL g1640 ( 
.A(n_1629),
.B(n_1603),
.C(n_1611),
.Y(n_1640)
);

OAI21xp33_ASAP7_75t_SL g1641 ( 
.A1(n_1634),
.A2(n_1603),
.B(n_1599),
.Y(n_1641)
);

NOR3xp33_ASAP7_75t_SL g1642 ( 
.A(n_1626),
.B(n_1619),
.C(n_1588),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1630),
.A2(n_1621),
.B(n_1604),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1635),
.A2(n_1563),
.B1(n_1561),
.B2(n_1575),
.C(n_1573),
.Y(n_1644)
);

AOI211xp5_ASAP7_75t_L g1645 ( 
.A1(n_1636),
.A2(n_1566),
.B(n_1565),
.C(n_1571),
.Y(n_1645)
);

AOI221x1_ASAP7_75t_L g1646 ( 
.A1(n_1626),
.A2(n_1570),
.B1(n_1569),
.B2(n_1516),
.C(n_1506),
.Y(n_1646)
);

AOI21xp33_ASAP7_75t_L g1647 ( 
.A1(n_1639),
.A2(n_1606),
.B(n_1476),
.Y(n_1647)
);

NOR2x1_ASAP7_75t_L g1648 ( 
.A(n_1638),
.B(n_1532),
.Y(n_1648)
);

XNOR2xp5_ASAP7_75t_L g1649 ( 
.A(n_1640),
.B(n_1308),
.Y(n_1649)
);

AOI221x1_ASAP7_75t_L g1650 ( 
.A1(n_1643),
.A2(n_1516),
.B1(n_1493),
.B2(n_1489),
.C(n_1494),
.Y(n_1650)
);

OAI31xp33_ASAP7_75t_L g1651 ( 
.A1(n_1642),
.A2(n_1476),
.A3(n_1470),
.B(n_1523),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1646),
.B(n_1471),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1650),
.B(n_1641),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1652),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1649),
.Y(n_1655)
);

OR3x1_ASAP7_75t_L g1656 ( 
.A(n_1647),
.B(n_1637),
.C(n_1645),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1651),
.B(n_1526),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1648),
.Y(n_1658)
);

NOR2x1_ASAP7_75t_L g1659 ( 
.A(n_1648),
.B(n_1529),
.Y(n_1659)
);

OAI21xp33_ASAP7_75t_SL g1660 ( 
.A1(n_1653),
.A2(n_1644),
.B(n_1529),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1654),
.A2(n_1541),
.B1(n_1476),
.B2(n_1470),
.Y(n_1661)
);

NOR4xp75_ASAP7_75t_L g1662 ( 
.A(n_1656),
.B(n_1537),
.C(n_1528),
.D(n_1503),
.Y(n_1662)
);

NOR2x1p5_ASAP7_75t_L g1663 ( 
.A(n_1655),
.B(n_1657),
.Y(n_1663)
);

OAI221xp5_ASAP7_75t_L g1664 ( 
.A1(n_1658),
.A2(n_1541),
.B1(n_1481),
.B2(n_1470),
.C(n_1501),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1660),
.B(n_1659),
.Y(n_1665)
);

NAND3x1_ASAP7_75t_L g1666 ( 
.A(n_1662),
.B(n_1494),
.C(n_1503),
.Y(n_1666)
);

AOI211xp5_ASAP7_75t_SL g1667 ( 
.A1(n_1663),
.A2(n_1471),
.B(n_1489),
.C(n_1493),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1666),
.Y(n_1668)
);

AOI322xp5_ASAP7_75t_L g1669 ( 
.A1(n_1668),
.A2(n_1665),
.A3(n_1661),
.B1(n_1667),
.B2(n_1664),
.C1(n_1503),
.C2(n_1501),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1669),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1669),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1670),
.B(n_1394),
.Y(n_1672)
);

A2O1A1Ixp33_ASAP7_75t_L g1673 ( 
.A1(n_1671),
.A2(n_1493),
.B(n_1489),
.C(n_1501),
.Y(n_1673)
);

XNOR2xp5_ASAP7_75t_L g1674 ( 
.A(n_1672),
.B(n_1487),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1673),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1675),
.A2(n_1481),
.B1(n_1477),
.B2(n_1482),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1676),
.A2(n_1674),
.B1(n_1481),
.B2(n_1501),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1677),
.B(n_1489),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_SL g1679 ( 
.A1(n_1678),
.A2(n_1493),
.B1(n_1481),
.B2(n_1319),
.Y(n_1679)
);

AO22x1_ASAP7_75t_L g1680 ( 
.A1(n_1679),
.A2(n_1306),
.B1(n_1483),
.B2(n_1333),
.Y(n_1680)
);

AOI211xp5_ASAP7_75t_L g1681 ( 
.A1(n_1680),
.A2(n_1336),
.B(n_1319),
.C(n_1526),
.Y(n_1681)
);


endmodule