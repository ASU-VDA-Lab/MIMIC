module fake_jpeg_9467_n_277 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_24),
.Y(n_50)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_33),
.B1(n_29),
.B2(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_58),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_33),
.B1(n_19),
.B2(n_24),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_62),
.B1(n_37),
.B2(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_55),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_32),
.B(n_34),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_8),
.C(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_25),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_65),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_61),
.B1(n_21),
.B2(n_19),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_33),
.B1(n_19),
.B2(n_21),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_33),
.B1(n_19),
.B2(n_21),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_71),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_40),
.B1(n_21),
.B2(n_42),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_72),
.B1(n_93),
.B2(n_63),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_68),
.B(n_77),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_29),
.B1(n_28),
.B2(n_20),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_75),
.A2(n_79),
.B1(n_82),
.B2(n_89),
.Y(n_119)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_81),
.Y(n_104)
);

AO22x1_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_38),
.B1(n_37),
.B2(n_36),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_29),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_87),
.Y(n_118)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_29),
.B1(n_28),
.B2(n_20),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_83),
.Y(n_117)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_90),
.Y(n_110)
);

AO22x1_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_28),
.B1(n_17),
.B2(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_65),
.A2(n_17),
.B1(n_22),
.B2(n_23),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_95),
.Y(n_112)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_54),
.A2(n_23),
.B1(n_20),
.B2(n_31),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_56),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_98),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_53),
.B(n_17),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_54),
.A2(n_31),
.B1(n_22),
.B2(n_23),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_22),
.B1(n_26),
.B2(n_32),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_63),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_101),
.B(n_114),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_103),
.A2(n_120),
.B1(n_125),
.B2(n_74),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_107),
.B(n_113),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_63),
.B1(n_54),
.B2(n_46),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_123),
.B1(n_80),
.B2(n_77),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_124),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_122),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_86),
.A2(n_47),
.B1(n_38),
.B2(n_46),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_139),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_130),
.B(n_131),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_104),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_133),
.B1(n_137),
.B2(n_145),
.Y(n_160)
);

AOI22x1_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_77),
.B1(n_68),
.B2(n_78),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_134),
.B(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_108),
.A2(n_85),
.B1(n_78),
.B2(n_83),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_26),
.B(n_27),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_95),
.B1(n_81),
.B2(n_66),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_47),
.B(n_70),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_138),
.A2(n_149),
.B(n_152),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_141),
.Y(n_166)
);

AO22x1_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_87),
.B1(n_76),
.B2(n_38),
.Y(n_142)
);

AO22x1_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_84),
.B1(n_38),
.B2(n_39),
.Y(n_168)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_146),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_121),
.B1(n_124),
.B2(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_39),
.B(n_87),
.C(n_27),
.D(n_41),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_30),
.C(n_18),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_123),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_32),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_165),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_153),
.B(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_158),
.B(n_183),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_125),
.B1(n_117),
.B2(n_107),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_169),
.B1(n_180),
.B2(n_128),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_SL g165 ( 
.A1(n_136),
.A2(n_117),
.A3(n_102),
.B1(n_116),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_168),
.A2(n_172),
.B(n_179),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_102),
.B1(n_100),
.B2(n_90),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_133),
.A2(n_70),
.B1(n_94),
.B2(n_38),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_131),
.B1(n_154),
.B2(n_155),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_26),
.B(n_111),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_152),
.B(n_139),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_41),
.C(n_111),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_178),
.C(n_184),
.Y(n_198)
);

XNOR2x1_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_148),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_18),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_156),
.A2(n_18),
.B(n_1),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_132),
.A2(n_18),
.B1(n_92),
.B2(n_0),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_143),
.C(n_135),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_188),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_186),
.B(n_194),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_189),
.B(n_203),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_160),
.A2(n_180),
.B1(n_182),
.B2(n_184),
.Y(n_190)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_199),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_200),
.B1(n_206),
.B2(n_179),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_160),
.B(n_146),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_150),
.Y(n_196)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_162),
.Y(n_214)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_171),
.A2(n_137),
.B1(n_142),
.B2(n_129),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_158),
.Y(n_201)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_204),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_172),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_150),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_161),
.A2(n_129),
.B1(n_142),
.B2(n_127),
.Y(n_206)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_178),
.C(n_175),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_213),
.C(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_167),
.C(n_162),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_220),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_173),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_176),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_167),
.B1(n_166),
.B2(n_177),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_222),
.B1(n_200),
.B2(n_199),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_192),
.A2(n_177),
.B1(n_159),
.B2(n_166),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_168),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_205),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_209),
.B(n_185),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_231),
.Y(n_244)
);

FAx1_ASAP7_75t_SL g226 ( 
.A(n_224),
.B(n_204),
.CI(n_197),
.CON(n_226),
.SN(n_226)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_226),
.B(n_234),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_215),
.A2(n_186),
.B(n_191),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_227),
.A2(n_232),
.B1(n_233),
.B2(n_223),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_207),
.A2(n_217),
.B1(n_208),
.B2(n_219),
.Y(n_230)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_218),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_188),
.B(n_206),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_205),
.B(n_189),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_229),
.C(n_224),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_196),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_220),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_236),
.A2(n_195),
.B(n_193),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_242),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_240),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_211),
.B(n_164),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_233),
.B(n_230),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_246),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_247),
.C(n_249),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_214),
.C(n_216),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_232),
.Y(n_248)
);

OAI221xp5_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_227),
.B1(n_237),
.B2(n_226),
.C(n_4),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_168),
.C(n_18),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_254),
.C(n_259),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_241),
.A2(n_226),
.B1(n_10),
.B2(n_3),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_11),
.Y(n_264)
);

AOI31xp33_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_240),
.A3(n_250),
.B(n_249),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_92),
.C(n_9),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_258),
.C(n_10),
.Y(n_262)
);

OAI221xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_16),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_255),
.A2(n_4),
.B(n_6),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_264),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_256),
.B(n_9),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_261),
.B(n_262),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_252),
.B(n_11),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_11),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_253),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_269),
.C(n_253),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_257),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_12),
.B(n_13),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_271),
.A2(n_268),
.B(n_266),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_273),
.C(n_12),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_12),
.C(n_13),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_275),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_14),
.C(n_16),
.Y(n_277)
);


endmodule