module real_jpeg_23092_n_32 (n_17, n_8, n_0, n_21, n_2, n_29, n_10, n_31, n_9, n_12, n_154, n_152, n_147, n_24, n_146, n_6, n_28, n_153, n_151, n_23, n_11, n_14, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_150, n_1, n_26, n_27, n_20, n_19, n_148, n_30, n_149, n_16, n_15, n_13, n_155, n_32);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_29;
input n_10;
input n_31;
input n_9;
input n_12;
input n_154;
input n_152;
input n_147;
input n_24;
input n_146;
input n_6;
input n_28;
input n_153;
input n_151;
input n_23;
input n_11;
input n_14;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_150;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_148;
input n_30;
input n_149;
input n_16;
input n_15;
input n_13;
input n_155;

output n_32;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_0),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_1),
.Y(n_102)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_4),
.B(n_52),
.C(n_101),
.Y(n_51)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_6),
.B(n_60),
.C(n_70),
.Y(n_59)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_7),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_8),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_9),
.B(n_54),
.C(n_94),
.Y(n_53)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_10),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_11),
.A2(n_33),
.B(n_144),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_11),
.B(n_37),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_12),
.Y(n_140)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_13),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_14),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_50),
.C(n_110),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_16),
.Y(n_129)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_17),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_18),
.Y(n_126)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_19),
.Y(n_115)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_22),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_24),
.B(n_58),
.C(n_77),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_25),
.B(n_48),
.C(n_121),
.Y(n_47)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_26),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_27),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_28),
.B(n_56),
.C(n_86),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_42),
.C(n_139),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_44),
.C(n_134),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_46),
.C(n_128),
.Y(n_45)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_41),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_38),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_38),
.B(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_38),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_38),
.B(n_122),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_39),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_43),
.C(n_136),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_45),
.C(n_130),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_123),
.C(n_124),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_112),
.C(n_113),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_104),
.C(n_105),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_97),
.C(n_98),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_89),
.C(n_90),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_80),
.C(n_81),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_73),
.C(n_74),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.C(n_65),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_138),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_146),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_147),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_148),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_149),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_150),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_151),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_152),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_153),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_154),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_155),
.Y(n_100)
);


endmodule