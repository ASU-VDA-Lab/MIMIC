module fake_netlist_6_3324_n_2073 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2073);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2073;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_322;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_474;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_206;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g205 ( 
.A(n_34),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_41),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_120),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_90),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_118),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_200),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_127),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_131),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_188),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_43),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_77),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_116),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_132),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_74),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_21),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_84),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_33),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_89),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_38),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_153),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_32),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_87),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_133),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_129),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_203),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_73),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_170),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_148),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_97),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_139),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_163),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_178),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_42),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_40),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_67),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_28),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_38),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_52),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_10),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_86),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_109),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_48),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_186),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_144),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_62),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_121),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_159),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_114),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_174),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_137),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_69),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_150),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_88),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_78),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_183),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_92),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_172),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_143),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_192),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_138),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_164),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_101),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_18),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_155),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_27),
.Y(n_273)
);

BUFx5_ASAP7_75t_L g274 ( 
.A(n_98),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_31),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_75),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_91),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_55),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_8),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_99),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_191),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_173),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_175),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_180),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_141),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_96),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_100),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_21),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_61),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_46),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_83),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_122),
.Y(n_292)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_69),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_43),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_46),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_16),
.Y(n_296)
);

BUFx8_ASAP7_75t_SL g297 ( 
.A(n_0),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_55),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_147),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_156),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_161),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_187),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_135),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_47),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_12),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_31),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_13),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_167),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_176),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_201),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_48),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_112),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_146),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_184),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_157),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_134),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_47),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_102),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_11),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_76),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_36),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_185),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_158),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_160),
.Y(n_324)
);

BUFx8_ASAP7_75t_SL g325 ( 
.A(n_166),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_16),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_93),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_51),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_6),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_94),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_204),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_72),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_6),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_113),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_123),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_72),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_35),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_7),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_51),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_35),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_140),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_45),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_63),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_106),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_8),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_9),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_103),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_64),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_126),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_18),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_57),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_1),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_169),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_154),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_190),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_14),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_145),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_67),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_29),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_52),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_26),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_57),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_165),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_189),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_49),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_22),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_108),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_42),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_2),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_54),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_162),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_197),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_115),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_66),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_56),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_32),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_15),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_66),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_22),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_71),
.Y(n_380)
);

CKINVDCx12_ASAP7_75t_R g381 ( 
.A(n_105),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_168),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_34),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_25),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_29),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_177),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_23),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_124),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_142),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_24),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_3),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_12),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_117),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_2),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_59),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_62),
.Y(n_396)
);

BUFx8_ASAP7_75t_SL g397 ( 
.A(n_179),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_15),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_64),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_107),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_54),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_61),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_136),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_104),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_10),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_194),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_130),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_356),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_405),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_356),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_356),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_261),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_356),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_325),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_356),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_395),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_405),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_395),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_395),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_395),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_266),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_395),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_205),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_351),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_268),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_351),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_276),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_334),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_397),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_384),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_384),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_365),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_274),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_205),
.Y(n_434)
);

INVxp33_ASAP7_75t_SL g435 ( 
.A(n_342),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_206),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_206),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_247),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_365),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_362),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_224),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_224),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_297),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_274),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_360),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_243),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_243),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_271),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_302),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_309),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_271),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_207),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_275),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_211),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_212),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_213),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_214),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_275),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_216),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_289),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_220),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_289),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_221),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_290),
.Y(n_464)
);

INVxp33_ASAP7_75t_L g465 ( 
.A(n_290),
.Y(n_465)
);

INVxp33_ASAP7_75t_L g466 ( 
.A(n_295),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_222),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_217),
.Y(n_468)
);

INVxp33_ASAP7_75t_SL g469 ( 
.A(n_226),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_223),
.Y(n_470)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_280),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_209),
.Y(n_472)
);

INVxp33_ASAP7_75t_SL g473 ( 
.A(n_228),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_295),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_305),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_305),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_306),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_225),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_227),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_280),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_209),
.Y(n_481)
);

INVxp33_ASAP7_75t_L g482 ( 
.A(n_306),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_241),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_329),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_242),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_252),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_329),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_232),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_332),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_233),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_332),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_234),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_336),
.Y(n_493)
);

BUFx2_ASAP7_75t_SL g494 ( 
.A(n_273),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_252),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_244),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_336),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_210),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_338),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_235),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_274),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_236),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_338),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_237),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_238),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_339),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_239),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_240),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_248),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_246),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_245),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_433),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_481),
.B(n_407),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_440),
.Y(n_514)
);

INVx6_ASAP7_75t_L g515 ( 
.A(n_472),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_440),
.Y(n_516)
);

BUFx8_ASAP7_75t_L g517 ( 
.A(n_417),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_408),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_486),
.B(n_251),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_408),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_410),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_410),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_411),
.B(n_406),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_411),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_433),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_413),
.B(n_256),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_413),
.B(n_404),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_415),
.B(n_284),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_415),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_433),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_416),
.B(n_258),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_416),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_418),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_418),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_472),
.B(n_284),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_472),
.B(n_495),
.Y(n_536)
);

NOR2x1_ASAP7_75t_L g537 ( 
.A(n_419),
.B(n_285),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_419),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_438),
.B(n_210),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_495),
.B(n_285),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_432),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_420),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_444),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_420),
.B(n_313),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_422),
.Y(n_545)
);

AND2x6_ASAP7_75t_L g546 ( 
.A(n_444),
.B(n_249),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_422),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_452),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_444),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_501),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_498),
.B(n_293),
.Y(n_551)
);

OA21x2_ASAP7_75t_L g552 ( 
.A1(n_501),
.A2(n_426),
.B(n_424),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_439),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_495),
.B(n_313),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_412),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_494),
.B(n_391),
.Y(n_556)
);

CKINVDCx6p67_ASAP7_75t_R g557 ( 
.A(n_438),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_434),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_501),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_454),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_423),
.B(n_318),
.Y(n_561)
);

AND2x6_ASAP7_75t_L g562 ( 
.A(n_436),
.B(n_249),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_494),
.B(n_318),
.Y(n_563)
);

BUFx8_ASAP7_75t_L g564 ( 
.A(n_417),
.Y(n_564)
);

CKINVDCx16_ASAP7_75t_R g565 ( 
.A(n_445),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_424),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_436),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_426),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_423),
.B(n_349),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_430),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_430),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_437),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_471),
.A2(n_250),
.B1(n_399),
.B2(n_401),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_456),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_475),
.B(n_349),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_437),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_431),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_467),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_431),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_441),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_441),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_435),
.B(n_229),
.Y(n_582)
);

AND3x1_ASAP7_75t_L g583 ( 
.A(n_409),
.B(n_340),
.C(n_339),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_475),
.B(n_355),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_442),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_442),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_468),
.A2(n_510),
.B1(n_425),
.B2(n_427),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_446),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_446),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_447),
.B(n_355),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_447),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_483),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_514),
.B(n_480),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_543),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_549),
.Y(n_595)
);

INVxp67_ASAP7_75t_SL g596 ( 
.A(n_514),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_552),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_549),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_552),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_549),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_559),
.Y(n_601)
);

AO21x2_ASAP7_75t_L g602 ( 
.A1(n_513),
.A2(n_215),
.B(n_208),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_559),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_552),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_546),
.Y(n_605)
);

BUFx4f_ASAP7_75t_L g606 ( 
.A(n_552),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_559),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_R g608 ( 
.A(n_548),
.B(n_414),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_516),
.B(n_428),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_556),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_543),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_516),
.B(n_445),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_543),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_513),
.B(n_469),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_536),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_517),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_551),
.B(n_498),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_512),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_515),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_512),
.Y(n_620)
);

AND2x2_ASAP7_75t_SL g621 ( 
.A(n_583),
.B(n_257),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_552),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_517),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_512),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_548),
.Y(n_625)
);

OAI22xp33_ASAP7_75t_L g626 ( 
.A1(n_551),
.A2(n_466),
.B1(n_482),
.B2(n_465),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_518),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_518),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_512),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_L g630 ( 
.A(n_573),
.B(n_587),
.C(n_582),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_519),
.B(n_473),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_520),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_582),
.B(n_455),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_512),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_543),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_520),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_563),
.B(n_461),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_525),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_525),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_556),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_519),
.B(n_463),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_578),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_543),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_525),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_525),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_543),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_525),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_536),
.B(n_470),
.Y(n_648)
);

OAI22x1_ASAP7_75t_L g649 ( 
.A1(n_539),
.A2(n_510),
.B1(n_468),
.B2(n_345),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_536),
.B(n_478),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_530),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_563),
.B(n_479),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_530),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_530),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_546),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_530),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_561),
.B(n_485),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_530),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_517),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_563),
.B(n_488),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_556),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_521),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_543),
.Y(n_663)
);

OR2x6_ASAP7_75t_L g664 ( 
.A(n_539),
.B(n_208),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_550),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_546),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_521),
.Y(n_667)
);

CKINVDCx6p67_ASAP7_75t_R g668 ( 
.A(n_557),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_561),
.B(n_492),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_542),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_550),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_550),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_L g673 ( 
.A(n_569),
.B(n_218),
.C(n_215),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_561),
.A2(n_391),
.B1(n_345),
.B2(n_358),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_550),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_542),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_550),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_545),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_522),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_515),
.B(n_561),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_545),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_575),
.B(n_500),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_515),
.B(n_502),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_522),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_592),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_575),
.B(n_504),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_515),
.B(n_575),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_546),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_560),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_575),
.B(n_505),
.Y(n_690)
);

INVx4_ASAP7_75t_L g691 ( 
.A(n_546),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_515),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_575),
.B(n_496),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_584),
.B(n_507),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_522),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_581),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_515),
.B(n_508),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_541),
.B(n_511),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_581),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_524),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_584),
.A2(n_358),
.B1(n_359),
.B2(n_340),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_524),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_581),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_581),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_560),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_541),
.B(n_443),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_524),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_583),
.A2(n_459),
.B1(n_490),
.B2(n_457),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_584),
.B(n_509),
.Y(n_709)
);

BUFx6f_ASAP7_75t_SL g710 ( 
.A(n_584),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_529),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_569),
.B(n_429),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_529),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_581),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_565),
.B(n_592),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_529),
.Y(n_716)
);

XOR2xp5_ASAP7_75t_L g717 ( 
.A(n_573),
.B(n_421),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_581),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_517),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_532),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_535),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_590),
.B(n_218),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_581),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_558),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_558),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_532),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_532),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_567),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_553),
.B(n_449),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_567),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_572),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_565),
.B(n_210),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_553),
.B(n_450),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_533),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_523),
.B(n_526),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_533),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_526),
.B(n_262),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_533),
.Y(n_738)
);

AND3x2_ASAP7_75t_L g739 ( 
.A(n_592),
.B(n_327),
.C(n_257),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_578),
.B(n_210),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_534),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_535),
.B(n_260),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_618),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_618),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_593),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_608),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_661),
.B(n_517),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_615),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_597),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_735),
.B(n_527),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_610),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_661),
.B(n_564),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_724),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_724),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_597),
.B(n_535),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_599),
.B(n_540),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_725),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_610),
.B(n_564),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_599),
.B(n_540),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_604),
.B(n_540),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_604),
.B(n_554),
.Y(n_761)
);

NOR2xp67_ASAP7_75t_L g762 ( 
.A(n_642),
.B(n_574),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_640),
.B(n_564),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_609),
.B(n_554),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_609),
.B(n_554),
.Y(n_765)
);

AO22x2_ASAP7_75t_L g766 ( 
.A1(n_630),
.A2(n_230),
.B1(n_231),
.B2(n_219),
.Y(n_766)
);

NAND2x1_ASAP7_75t_L g767 ( 
.A(n_605),
.B(n_546),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_640),
.B(n_564),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_725),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_626),
.B(n_527),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_701),
.A2(n_361),
.B1(n_379),
.B2(n_359),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_721),
.B(n_590),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_596),
.B(n_557),
.Y(n_773)
);

NOR3xp33_ASAP7_75t_L g774 ( 
.A(n_617),
.B(n_587),
.C(n_708),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_614),
.B(n_531),
.Y(n_775)
);

NAND2x1p5_ASAP7_75t_L g776 ( 
.A(n_606),
.B(n_528),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_728),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_631),
.B(n_528),
.Y(n_778)
);

BUFx2_ASAP7_75t_L g779 ( 
.A(n_685),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_721),
.B(n_528),
.Y(n_780)
);

BUFx5_ASAP7_75t_L g781 ( 
.A(n_622),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_737),
.B(n_544),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_618),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_641),
.B(n_557),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_620),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_685),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_693),
.B(n_574),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_622),
.B(n_544),
.Y(n_788)
);

OR2x2_ASAP7_75t_SL g789 ( 
.A(n_706),
.B(n_361),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_648),
.B(n_555),
.Y(n_790)
);

BUFx8_ASAP7_75t_L g791 ( 
.A(n_616),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_657),
.B(n_669),
.Y(n_792)
);

BUFx5_ASAP7_75t_L g793 ( 
.A(n_619),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_682),
.B(n_331),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_693),
.B(n_590),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_730),
.B(n_544),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_698),
.Y(n_797)
);

NOR3xp33_ASAP7_75t_L g798 ( 
.A(n_612),
.B(n_259),
.C(n_253),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_620),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_698),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_712),
.B(n_590),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_625),
.Y(n_802)
);

OR2x6_ASAP7_75t_L g803 ( 
.A(n_616),
.B(n_379),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_706),
.B(n_576),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_650),
.B(n_555),
.Y(n_805)
);

NOR2x1p5_ASAP7_75t_L g806 ( 
.A(n_668),
.B(n_278),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_729),
.B(n_586),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_606),
.B(n_544),
.Y(n_808)
);

BUFx8_ASAP7_75t_L g809 ( 
.A(n_623),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_621),
.B(n_263),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_606),
.B(n_544),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_621),
.B(n_264),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_606),
.B(n_602),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_620),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_624),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_680),
.A2(n_537),
.B(n_546),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_730),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_731),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_L g819 ( 
.A(n_709),
.B(n_715),
.C(n_733),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_621),
.B(n_267),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_637),
.B(n_269),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_602),
.B(n_566),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_652),
.B(n_270),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_731),
.B(n_566),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_633),
.B(n_279),
.Y(n_825)
);

OR2x6_ASAP7_75t_L g826 ( 
.A(n_623),
.B(n_385),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_660),
.B(n_288),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_686),
.B(n_282),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_664),
.A2(n_283),
.B1(n_286),
.B2(n_291),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_690),
.B(n_300),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_694),
.B(n_294),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_673),
.A2(n_589),
.B(n_586),
.C(n_394),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_627),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_602),
.A2(n_327),
.B1(n_364),
.B2(n_400),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_674),
.B(n_303),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_628),
.B(n_566),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_659),
.B(n_719),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_722),
.B(n_589),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_632),
.B(n_636),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_664),
.B(n_296),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_619),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_636),
.B(n_566),
.Y(n_842)
);

NAND2x1p5_ASAP7_75t_L g843 ( 
.A(n_605),
.B(n_219),
.Y(n_843)
);

BUFx6f_ASAP7_75t_SL g844 ( 
.A(n_664),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_649),
.B(n_308),
.Y(n_845)
);

BUFx5_ASAP7_75t_L g846 ( 
.A(n_619),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_602),
.A2(n_364),
.B1(n_400),
.B2(n_353),
.Y(n_847)
);

OAI221xp5_ASAP7_75t_L g848 ( 
.A1(n_664),
.A2(n_385),
.B1(n_394),
.B2(n_398),
.C(n_396),
.Y(n_848)
);

O2A1O1Ixp5_ASAP7_75t_L g849 ( 
.A1(n_687),
.A2(n_265),
.B(n_255),
.C(n_254),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_662),
.B(n_566),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_664),
.B(n_448),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_624),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_662),
.B(n_667),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_667),
.B(n_568),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_689),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_659),
.B(n_448),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_740),
.B(n_298),
.Y(n_857)
);

BUFx5_ASAP7_75t_L g858 ( 
.A(n_692),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_710),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_649),
.B(n_310),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_670),
.B(n_568),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_719),
.B(n_312),
.Y(n_862)
);

BUFx5_ASAP7_75t_L g863 ( 
.A(n_692),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_742),
.B(n_314),
.Y(n_864)
);

NAND2xp33_ASAP7_75t_L g865 ( 
.A(n_683),
.B(n_274),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_624),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_670),
.B(n_676),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_710),
.A2(n_315),
.B1(n_324),
.B2(n_363),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_676),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_722),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_739),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_732),
.B(n_304),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_605),
.B(n_344),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_629),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_678),
.B(n_568),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_668),
.B(n_451),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_678),
.B(n_568),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_629),
.Y(n_878)
);

NAND2xp33_ASAP7_75t_L g879 ( 
.A(n_697),
.B(n_681),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_710),
.A2(n_353),
.B1(n_231),
.B2(n_254),
.Y(n_880)
);

OR2x6_ASAP7_75t_L g881 ( 
.A(n_722),
.B(n_396),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_629),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_671),
.B(n_568),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_681),
.Y(n_884)
);

OR2x6_ASAP7_75t_L g885 ( 
.A(n_722),
.B(n_398),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_710),
.A2(n_354),
.B1(n_371),
.B2(n_382),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_605),
.B(n_372),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_692),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_671),
.B(n_571),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_717),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_722),
.B(n_307),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_705),
.B(n_311),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_671),
.A2(n_373),
.B1(n_388),
.B2(n_389),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_671),
.B(n_571),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_679),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_595),
.B(n_571),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_679),
.Y(n_897)
);

AO22x2_ASAP7_75t_L g898 ( 
.A1(n_717),
.A2(n_230),
.B1(n_255),
.B2(n_265),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_679),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_594),
.B(n_317),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_634),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_655),
.B(n_249),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_594),
.B(n_319),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_655),
.A2(n_376),
.B1(n_321),
.B2(n_326),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_594),
.B(n_571),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_595),
.B(n_571),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_655),
.B(n_666),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_838),
.B(n_451),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_779),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_753),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_807),
.B(n_453),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_751),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_750),
.B(n_594),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_772),
.Y(n_914)
);

BUFx4f_ASAP7_75t_L g915 ( 
.A(n_786),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_743),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_754),
.Y(n_917)
);

INVx8_ASAP7_75t_L g918 ( 
.A(n_881),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_744),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_757),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_841),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_838),
.B(n_453),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_775),
.B(n_613),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_781),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_769),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_783),
.Y(n_926)
);

AO22x1_ASAP7_75t_L g927 ( 
.A1(n_774),
.A2(n_377),
.B1(n_380),
.B2(n_378),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_781),
.B(n_655),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_841),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_777),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_770),
.A2(n_691),
.B1(n_666),
.B2(n_688),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_764),
.B(n_613),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_772),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_781),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_802),
.Y(n_935)
);

NAND2xp33_ASAP7_75t_SL g936 ( 
.A(n_844),
.B(n_328),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_781),
.B(n_813),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_745),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_785),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_781),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_841),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_799),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_781),
.B(n_813),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_797),
.B(n_458),
.Y(n_944)
);

NOR3xp33_ASAP7_75t_SL g945 ( 
.A(n_845),
.B(n_337),
.C(n_333),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_765),
.B(n_613),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_895),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_748),
.B(n_458),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_871),
.B(n_460),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_749),
.B(n_778),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_755),
.B(n_613),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_808),
.B(n_688),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_804),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_755),
.B(n_635),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_888),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_817),
.Y(n_956)
);

INVx4_ASAP7_75t_L g957 ( 
.A(n_888),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_876),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_818),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_800),
.B(n_635),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_833),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_756),
.B(n_635),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_789),
.B(n_787),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_756),
.B(n_635),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_R g965 ( 
.A(n_746),
.B(n_381),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_856),
.B(n_460),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_814),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_773),
.B(n_462),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_792),
.A2(n_718),
.B1(n_696),
.B2(n_699),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_815),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_870),
.B(n_462),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_888),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_759),
.B(n_643),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_811),
.B(n_611),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_790),
.B(n_643),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_801),
.A2(n_795),
.B1(n_812),
.B2(n_810),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_820),
.A2(n_718),
.B1(n_696),
.B2(n_699),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_869),
.Y(n_978)
);

AND2x2_ASAP7_75t_SL g979 ( 
.A(n_847),
.B(n_272),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_884),
.B(n_881),
.Y(n_980)
);

BUFx8_ASAP7_75t_SL g981 ( 
.A(n_855),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_859),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_852),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_866),
.Y(n_984)
);

NOR3xp33_ASAP7_75t_SL g985 ( 
.A(n_860),
.B(n_346),
.C(n_343),
.Y(n_985)
);

NAND2xp33_ASAP7_75t_L g986 ( 
.A(n_793),
.B(n_611),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_759),
.B(n_643),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_883),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_851),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_892),
.B(n_464),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_805),
.B(n_643),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_881),
.B(n_464),
.Y(n_992)
);

OAI221xp5_ASAP7_75t_L g993 ( 
.A1(n_840),
.A2(n_348),
.B1(n_350),
.B2(n_352),
.C(n_366),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_791),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_889),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_782),
.B(n_611),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_885),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_819),
.B(n_611),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_760),
.B(n_611),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_760),
.B(n_646),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_766),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_766),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_889),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_885),
.B(n_474),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_803),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_761),
.A2(n_393),
.B1(n_281),
.B2(n_272),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_784),
.B(n_663),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_761),
.B(n_663),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_R g1009 ( 
.A(n_859),
.B(n_381),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_794),
.B(n_663),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_776),
.B(n_646),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_839),
.B(n_663),
.Y(n_1012)
);

NAND2x1p5_ASAP7_75t_L g1013 ( 
.A(n_767),
.B(n_723),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_885),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_897),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_766),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_890),
.B(n_474),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_776),
.B(n_646),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_853),
.B(n_646),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_803),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_894),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_874),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_780),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_894),
.Y(n_1024)
);

OR2x4_ASAP7_75t_L g1025 ( 
.A(n_872),
.B(n_476),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_825),
.B(n_703),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_791),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_837),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_878),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_867),
.B(n_646),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_882),
.Y(n_1031)
);

OR2x6_ASAP7_75t_L g1032 ( 
.A(n_758),
.B(n_281),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_824),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_836),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_796),
.B(n_788),
.Y(n_1035)
);

BUFx4f_ASAP7_75t_L g1036 ( 
.A(n_803),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_842),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_809),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_848),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_899),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_821),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_879),
.A2(n_704),
.B1(n_714),
.B2(n_644),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_843),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_809),
.Y(n_1044)
);

OR2x6_ASAP7_75t_L g1045 ( 
.A(n_763),
.B(n_287),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_834),
.A2(n_771),
.B1(n_822),
.B2(n_898),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_907),
.A2(n_723),
.B(n_714),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_831),
.A2(n_704),
.B1(n_639),
.B2(n_644),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_768),
.B(n_747),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_827),
.A2(n_638),
.B1(n_639),
.B2(n_644),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_816),
.B(n_723),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_901),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_SL g1053 ( 
.A(n_904),
.B(n_369),
.C(n_368),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_850),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_752),
.B(n_476),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_843),
.Y(n_1056)
);

NAND3xp33_ASAP7_75t_L g1057 ( 
.A(n_857),
.B(n_374),
.C(n_370),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_896),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_844),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_896),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_854),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_806),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_861),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_900),
.B(n_903),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_891),
.A2(n_638),
.B1(n_639),
.B2(n_645),
.Y(n_1065)
);

NOR2xp67_ASAP7_75t_L g1066 ( 
.A(n_829),
.B(n_638),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_823),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_771),
.A2(n_330),
.B1(n_403),
.B2(n_393),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_816),
.B(n_723),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_904),
.B(n_645),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_822),
.B(n_723),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_798),
.A2(n_645),
.B1(n_647),
.B2(n_651),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_875),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_877),
.Y(n_1074)
);

OR2x6_ASAP7_75t_L g1075 ( 
.A(n_826),
.B(n_287),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_826),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_826),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_906),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_906),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_862),
.B(n_477),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_793),
.B(n_723),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_793),
.B(n_647),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_898),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_828),
.B(n_647),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_793),
.B(n_598),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_793),
.B(n_598),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_793),
.B(n_651),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_846),
.B(n_598),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_873),
.A2(n_653),
.B(n_651),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_846),
.B(n_600),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_L g1091 ( 
.A(n_990),
.B(n_968),
.C(n_993),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_958),
.B(n_762),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_986),
.A2(n_887),
.B(n_902),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1046),
.A2(n_880),
.B1(n_898),
.B2(n_830),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_915),
.B(n_868),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_910),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1046),
.A2(n_886),
.B1(n_835),
.B2(n_832),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1064),
.A2(n_865),
.B(n_858),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_980),
.B(n_864),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_981),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_979),
.A2(n_905),
.B1(n_330),
.B2(n_335),
.Y(n_1101)
);

OAI21xp33_ASAP7_75t_SL g1102 ( 
.A1(n_937),
.A2(n_299),
.B(n_292),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_909),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_1026),
.A2(n_849),
.B(n_893),
.C(n_323),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_917),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_950),
.B(n_863),
.Y(n_1106)
);

XNOR2xp5_ASAP7_75t_L g1107 ( 
.A(n_935),
.B(n_537),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_920),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1035),
.A2(n_858),
.B(n_846),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1051),
.A2(n_601),
.B(n_600),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1049),
.A2(n_863),
.B1(n_858),
.B2(n_846),
.Y(n_1111)
);

INVx4_ASAP7_75t_L g1112 ( 
.A(n_921),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_928),
.A2(n_858),
.B(n_846),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1026),
.A2(n_322),
.B(n_323),
.C(n_341),
.Y(n_1114)
);

INVx1_ASAP7_75t_SL g1115 ( 
.A(n_909),
.Y(n_1115)
);

O2A1O1Ixp5_ASAP7_75t_SL g1116 ( 
.A1(n_998),
.A2(n_477),
.B(n_484),
.C(n_487),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_979),
.A2(n_320),
.B1(n_403),
.B2(n_292),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_921),
.Y(n_1118)
);

NAND2x1p5_ASAP7_75t_L g1119 ( 
.A(n_957),
.B(n_726),
.Y(n_1119)
);

BUFx8_ASAP7_75t_L g1120 ( 
.A(n_994),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_980),
.B(n_484),
.Y(n_1121)
);

INVx6_ASAP7_75t_L g1122 ( 
.A(n_994),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_921),
.Y(n_1123)
);

OAI21xp33_ASAP7_75t_L g1124 ( 
.A1(n_911),
.A2(n_966),
.B(n_953),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_1028),
.B(n_375),
.Y(n_1125)
);

AOI21x1_ASAP7_75t_L g1126 ( 
.A1(n_974),
.A2(n_695),
.B(n_684),
.Y(n_1126)
);

BUFx4_ASAP7_75t_SL g1127 ( 
.A(n_1027),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1068),
.A2(n_316),
.B1(n_301),
.B2(n_320),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1068),
.A2(n_301),
.B1(n_299),
.B2(n_316),
.Y(n_1129)
);

OAI22x1_ASAP7_75t_L g1130 ( 
.A1(n_1083),
.A2(n_402),
.B1(n_383),
.B2(n_387),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_915),
.B(n_863),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_947),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_908),
.B(n_487),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_908),
.B(n_489),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1023),
.B(n_846),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1023),
.B(n_988),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_928),
.A2(n_863),
.B(n_858),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_929),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_952),
.A2(n_863),
.B(n_858),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_925),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1001),
.A2(n_367),
.B1(n_357),
.B2(n_347),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_912),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_995),
.B(n_600),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1003),
.B(n_601),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_966),
.B(n_489),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_929),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_976),
.A2(n_322),
.B(n_367),
.C(n_357),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1049),
.B(n_989),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_912),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_1044),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1021),
.B(n_601),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_952),
.A2(n_656),
.B(n_675),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_929),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1024),
.B(n_603),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_914),
.B(n_653),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1002),
.A2(n_1016),
.B1(n_1039),
.B2(n_913),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_SL g1157 ( 
.A1(n_918),
.A2(n_1036),
.B1(n_1041),
.B2(n_1032),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_914),
.B(n_653),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_930),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_975),
.B(n_603),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_975),
.B(n_603),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_938),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_956),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_929),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_922),
.B(n_491),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_933),
.A2(n_1080),
.B1(n_922),
.B2(n_1055),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_982),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1039),
.A2(n_335),
.B(n_341),
.C(n_347),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_937),
.A2(n_654),
.B(n_675),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_933),
.B(n_654),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_947),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1055),
.B(n_656),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_991),
.B(n_607),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_943),
.A2(n_658),
.B(n_665),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_971),
.B(n_491),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_959),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_991),
.A2(n_658),
.B(n_672),
.C(n_665),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_963),
.B(n_390),
.Y(n_1178)
);

INVx2_ASAP7_75t_SL g1179 ( 
.A(n_944),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1078),
.B(n_607),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_1017),
.Y(n_1181)
);

CKINVDCx6p67_ASAP7_75t_R g1182 ( 
.A(n_1027),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_943),
.A2(n_658),
.B(n_665),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_938),
.Y(n_1184)
);

NAND4xp25_ASAP7_75t_SL g1185 ( 
.A(n_1057),
.B(n_493),
.C(n_497),
.D(n_499),
.Y(n_1185)
);

OR2x6_ASAP7_75t_SL g1186 ( 
.A(n_1059),
.B(n_392),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_982),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1070),
.A2(n_672),
.B(n_677),
.C(n_607),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1080),
.A2(n_249),
.B1(n_277),
.B2(n_386),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1079),
.B(n_580),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1019),
.A2(n_1030),
.B(n_1085),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_998),
.A2(n_591),
.B(n_588),
.C(n_585),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1086),
.A2(n_672),
.B(n_677),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_1038),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1060),
.B(n_580),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1025),
.B(n_726),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1088),
.A2(n_726),
.B(n_734),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_982),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1090),
.A2(n_1081),
.B(n_996),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1015),
.Y(n_1200)
);

BUFx5_ASAP7_75t_L g1201 ( 
.A(n_1033),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1067),
.A2(n_734),
.B1(n_726),
.B2(n_588),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1006),
.A2(n_591),
.B(n_580),
.C(n_585),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1032),
.A2(n_734),
.B1(n_588),
.B2(n_591),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1032),
.A2(n_585),
.B(n_497),
.C(n_499),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1015),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_961),
.Y(n_1207)
);

OR2x6_ASAP7_75t_L g1208 ( 
.A(n_918),
.B(n_493),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_SL g1209 ( 
.A(n_965),
.B(n_503),
.C(n_506),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_R g1210 ( 
.A(n_1062),
.B(n_79),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1045),
.A2(n_503),
.B(n_506),
.C(n_736),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1025),
.B(n_734),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_971),
.B(n_570),
.Y(n_1213)
);

NOR3xp33_ASAP7_75t_SL g1214 ( 
.A(n_936),
.B(n_0),
.C(n_1),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1060),
.B(n_684),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1058),
.B(n_923),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1051),
.A2(n_741),
.B(n_738),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1077),
.Y(n_1218)
);

BUFx8_ASAP7_75t_SL g1219 ( 
.A(n_1005),
.Y(n_1219)
);

O2A1O1Ixp5_ASAP7_75t_SL g1220 ( 
.A1(n_1071),
.A2(n_274),
.B(n_4),
.C(n_5),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_978),
.B(n_684),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1045),
.A2(n_741),
.B(n_738),
.C(n_736),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_982),
.Y(n_1223)
);

AOI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1045),
.A2(n_736),
.B1(n_727),
.B2(n_720),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1066),
.A2(n_727),
.B1(n_720),
.B2(n_716),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1040),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1034),
.B(n_695),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_948),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_948),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1081),
.A2(n_727),
.B(n_720),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_SL g1231 ( 
.A(n_1036),
.B(n_249),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_SL g1232 ( 
.A1(n_1007),
.A2(n_716),
.B(n_713),
.C(n_711),
.Y(n_1232)
);

INVxp67_ASAP7_75t_L g1233 ( 
.A(n_949),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1040),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_965),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1077),
.B(n_3),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1020),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_997),
.B(n_570),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1014),
.B(n_4),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1076),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_957),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1022),
.Y(n_1242)
);

BUFx8_ASAP7_75t_SL g1243 ( 
.A(n_1075),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1014),
.B(n_5),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1037),
.B(n_695),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1126),
.A2(n_1089),
.B(n_1047),
.Y(n_1246)
);

NOR4xp25_ASAP7_75t_L g1247 ( 
.A(n_1094),
.B(n_1071),
.C(n_1070),
.D(n_1069),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1147),
.A2(n_1007),
.A3(n_1084),
.B(n_1010),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1136),
.B(n_1054),
.Y(n_1249)
);

NOR2x1_ASAP7_75t_L g1250 ( 
.A(n_1100),
.B(n_1241),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1216),
.B(n_1156),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1156),
.B(n_1061),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1118),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1096),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1109),
.A2(n_934),
.B(n_924),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1201),
.B(n_1063),
.Y(n_1256)
);

OA22x2_ASAP7_75t_L g1257 ( 
.A1(n_1181),
.A2(n_1075),
.B1(n_949),
.B2(n_1004),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1091),
.A2(n_985),
.B(n_945),
.C(n_1053),
.Y(n_1258)
);

INVx5_ASAP7_75t_L g1259 ( 
.A(n_1118),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1091),
.A2(n_1069),
.B(n_1000),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1181),
.B(n_1075),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1115),
.B(n_992),
.Y(n_1262)
);

AO21x2_ASAP7_75t_L g1263 ( 
.A1(n_1232),
.A2(n_1018),
.B(n_1011),
.Y(n_1263)
);

NOR2x1_ASAP7_75t_SL g1264 ( 
.A(n_1131),
.B(n_1043),
.Y(n_1264)
);

OR2x6_ASAP7_75t_L g1265 ( 
.A(n_1208),
.B(n_918),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1106),
.A2(n_934),
.B(n_924),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1201),
.B(n_1073),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1104),
.A2(n_1084),
.A3(n_1010),
.B(n_940),
.Y(n_1268)
);

AOI22x1_ASAP7_75t_L g1269 ( 
.A1(n_1098),
.A2(n_1074),
.B1(n_1056),
.B2(n_916),
.Y(n_1269)
);

AOI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1191),
.A2(n_1199),
.B(n_1161),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1093),
.A2(n_1139),
.B(n_1137),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1113),
.A2(n_940),
.B(n_1011),
.Y(n_1272)
);

AO21x2_ASAP7_75t_L g1273 ( 
.A1(n_1160),
.A2(n_1018),
.B(n_999),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1111),
.A2(n_1043),
.B(n_1012),
.Y(n_1274)
);

INVx4_ASAP7_75t_L g1275 ( 
.A(n_1118),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1132),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1169),
.A2(n_1087),
.B(n_1082),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1171),
.Y(n_1278)
);

AOI221xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1094),
.A2(n_960),
.B1(n_946),
.B2(n_932),
.C(n_987),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1173),
.A2(n_1043),
.B(n_1056),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1145),
.B(n_992),
.Y(n_1281)
);

NAND2xp33_ASAP7_75t_R g1282 ( 
.A(n_1235),
.B(n_1053),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1175),
.B(n_1004),
.Y(n_1283)
);

NAND2xp33_ASAP7_75t_SL g1284 ( 
.A(n_1210),
.B(n_945),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1200),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1105),
.Y(n_1286)
);

OAI22x1_ASAP7_75t_L g1287 ( 
.A1(n_1239),
.A2(n_1244),
.B1(n_1236),
.B2(n_1099),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1201),
.B(n_951),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1177),
.A2(n_977),
.B(n_954),
.Y(n_1289)
);

OAI21xp33_ASAP7_75t_L g1290 ( 
.A1(n_1178),
.A2(n_985),
.B(n_1009),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1206),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1174),
.A2(n_1087),
.B(n_1082),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1115),
.B(n_927),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1201),
.B(n_962),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1117),
.A2(n_1166),
.B1(n_1101),
.B2(n_1189),
.Y(n_1295)
);

NAND3xp33_ASAP7_75t_L g1296 ( 
.A(n_1097),
.B(n_960),
.C(n_969),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1114),
.A2(n_964),
.A3(n_973),
.B(n_1008),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1146),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1183),
.A2(n_1042),
.B(n_1013),
.Y(n_1299)
);

NOR4xp25_ASAP7_75t_L g1300 ( 
.A(n_1168),
.B(n_942),
.C(n_1052),
.D(n_1029),
.Y(n_1300)
);

CKINVDCx11_ASAP7_75t_R g1301 ( 
.A(n_1186),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1142),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1108),
.Y(n_1303)
);

AO21x2_ASAP7_75t_L g1304 ( 
.A1(n_1217),
.A2(n_1048),
.B(n_1065),
.Y(n_1304)
);

NOR2xp67_ASAP7_75t_SL g1305 ( 
.A(n_1122),
.B(n_941),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_SL g1306 ( 
.A1(n_1222),
.A2(n_1072),
.B(n_1050),
.Y(n_1306)
);

AOI31xp67_ASAP7_75t_L g1307 ( 
.A1(n_1225),
.A2(n_926),
.A3(n_939),
.B(n_967),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1201),
.B(n_1022),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1226),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1135),
.A2(n_931),
.B(n_1013),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1099),
.A2(n_941),
.B1(n_955),
.B2(n_972),
.Y(n_1311)
);

INVxp67_ASAP7_75t_L g1312 ( 
.A(n_1149),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1195),
.A2(n_972),
.B(n_955),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1101),
.A2(n_1031),
.B1(n_919),
.B2(n_984),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1175),
.B(n_1009),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1230),
.A2(n_1031),
.B(n_983),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1110),
.A2(n_970),
.B(n_711),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1179),
.B(n_577),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1245),
.A2(n_707),
.B(n_702),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1110),
.A2(n_707),
.B(n_702),
.Y(n_1320)
);

OAI21xp33_ASAP7_75t_L g1321 ( 
.A1(n_1125),
.A2(n_277),
.B(n_386),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1127),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1217),
.A2(n_707),
.B(n_702),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1245),
.A2(n_700),
.B(n_386),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1229),
.B(n_577),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1116),
.A2(n_700),
.B(n_534),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1234),
.B(n_700),
.Y(n_1327)
);

AO31x2_ASAP7_75t_L g1328 ( 
.A1(n_1097),
.A2(n_538),
.A3(n_534),
.B(n_547),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1190),
.B(n_577),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1188),
.A2(n_538),
.B(n_547),
.Y(n_1330)
);

INVx1_ASAP7_75t_SL g1331 ( 
.A(n_1162),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1140),
.B(n_579),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1159),
.B(n_579),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1103),
.B(n_7),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1133),
.B(n_579),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1228),
.B(n_171),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1163),
.B(n_579),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_1120),
.Y(n_1338)
);

AOI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1197),
.A2(n_538),
.B(n_547),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1133),
.B(n_579),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1124),
.B(n_9),
.Y(n_1341)
);

AO32x2_ASAP7_75t_L g1342 ( 
.A1(n_1128),
.A2(n_11),
.A3(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1176),
.B(n_579),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1122),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1107),
.B(n_579),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1215),
.A2(n_1227),
.B(n_1180),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1152),
.A2(n_274),
.B(n_277),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1193),
.A2(n_274),
.B(n_277),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1148),
.B(n_151),
.Y(n_1349)
);

OAI22x1_ASAP7_75t_L g1350 ( 
.A1(n_1218),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1237),
.Y(n_1351)
);

AND2x6_ASAP7_75t_L g1352 ( 
.A(n_1167),
.B(n_386),
.Y(n_1352)
);

AOI221xp5_ASAP7_75t_L g1353 ( 
.A1(n_1128),
.A2(n_1129),
.B1(n_1130),
.B2(n_1209),
.C(n_1233),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_SL g1354 ( 
.A(n_1121),
.B(n_274),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1143),
.A2(n_277),
.B(n_386),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1144),
.A2(n_274),
.B(n_562),
.Y(n_1356)
);

AOI221x1_ASAP7_75t_L g1357 ( 
.A1(n_1129),
.A2(n_19),
.B1(n_20),
.B2(n_23),
.C(n_24),
.Y(n_1357)
);

INVxp67_ASAP7_75t_L g1358 ( 
.A(n_1184),
.Y(n_1358)
);

BUFx10_ASAP7_75t_L g1359 ( 
.A(n_1150),
.Y(n_1359)
);

AOI211x1_ASAP7_75t_L g1360 ( 
.A1(n_1207),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1134),
.B(n_28),
.Y(n_1361)
);

O2A1O1Ixp33_ASAP7_75t_SL g1362 ( 
.A1(n_1095),
.A2(n_202),
.B(n_199),
.C(n_198),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1213),
.B(n_30),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_SL g1364 ( 
.A(n_1121),
.B(n_30),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1213),
.B(n_33),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1240),
.Y(n_1366)
);

NAND3xp33_ASAP7_75t_SL g1367 ( 
.A(n_1157),
.B(n_36),
.C(n_37),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1151),
.B(n_546),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1192),
.A2(n_119),
.B(n_81),
.Y(n_1369)
);

AO31x2_ASAP7_75t_L g1370 ( 
.A1(n_1196),
.A2(n_562),
.A3(n_546),
.B(n_40),
.Y(n_1370)
);

AO31x2_ASAP7_75t_L g1371 ( 
.A1(n_1212),
.A2(n_562),
.A3(n_546),
.B(n_41),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1154),
.B(n_562),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1221),
.A2(n_111),
.B(n_196),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1238),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1242),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1165),
.B(n_1208),
.Y(n_1376)
);

NOR2x1_ASAP7_75t_SL g1377 ( 
.A(n_1146),
.B(n_193),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1219),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1223),
.B(n_1141),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1165),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1231),
.B(n_37),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1223),
.B(n_562),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1102),
.A2(n_39),
.B(n_44),
.C(n_45),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1231),
.A2(n_39),
.B(n_44),
.C(n_49),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1194),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1241),
.Y(n_1386)
);

INVx5_ASAP7_75t_L g1387 ( 
.A(n_1146),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_R g1388 ( 
.A(n_1182),
.B(n_181),
.Y(n_1388)
);

OAI22x1_ASAP7_75t_L g1389 ( 
.A1(n_1185),
.A2(n_50),
.B1(n_53),
.B2(n_56),
.Y(n_1389)
);

AOI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1155),
.A2(n_562),
.B(n_152),
.Y(n_1390)
);

AO32x2_ASAP7_75t_L g1391 ( 
.A1(n_1220),
.A2(n_50),
.A3(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1172),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1203),
.A2(n_562),
.B(n_80),
.Y(n_1393)
);

AO21x2_ASAP7_75t_L g1394 ( 
.A1(n_1224),
.A2(n_125),
.B(n_110),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1120),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1119),
.A2(n_95),
.B(n_85),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1119),
.A2(n_82),
.B(n_562),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1158),
.A2(n_1170),
.B(n_1202),
.Y(n_1398)
);

AND2x6_ASAP7_75t_L g1399 ( 
.A(n_1167),
.B(n_1187),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1211),
.A2(n_58),
.B(n_60),
.C(n_63),
.Y(n_1400)
);

AO31x2_ASAP7_75t_L g1401 ( 
.A1(n_1112),
.A2(n_562),
.A3(n_65),
.B(n_68),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1208),
.A2(n_60),
.B1(n_65),
.B2(n_68),
.Y(n_1402)
);

INVx6_ASAP7_75t_L g1403 ( 
.A(n_1167),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1123),
.B(n_562),
.Y(n_1404)
);

OAI21xp33_ASAP7_75t_L g1405 ( 
.A1(n_1214),
.A2(n_70),
.B(n_71),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1092),
.B(n_1112),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1123),
.A2(n_70),
.B(n_1138),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1138),
.A2(n_1153),
.B(n_1164),
.Y(n_1408)
);

AO21x2_ASAP7_75t_L g1409 ( 
.A1(n_1271),
.A2(n_1204),
.B(n_1205),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1254),
.Y(n_1410)
);

OR3x4_ASAP7_75t_SL g1411 ( 
.A(n_1402),
.B(n_1243),
.C(n_1187),
.Y(n_1411)
);

AO31x2_ASAP7_75t_L g1412 ( 
.A1(n_1357),
.A2(n_1153),
.A3(n_1164),
.B(n_1187),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1296),
.A2(n_1198),
.B(n_1258),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1246),
.A2(n_1198),
.B(n_1339),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1331),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1249),
.B(n_1198),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1286),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1296),
.A2(n_1295),
.B(n_1290),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1303),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1344),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1268),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1367),
.A2(n_1405),
.B1(n_1402),
.B2(n_1287),
.Y(n_1422)
);

INVx5_ASAP7_75t_L g1423 ( 
.A(n_1399),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1269),
.A2(n_1255),
.B(n_1272),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1300),
.A2(n_1260),
.B(n_1270),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1295),
.A2(n_1260),
.B(n_1310),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_SL g1427 ( 
.A1(n_1264),
.A2(n_1252),
.B(n_1377),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1374),
.B(n_1380),
.Y(n_1428)
);

NAND3xp33_ASAP7_75t_L g1429 ( 
.A(n_1353),
.B(n_1341),
.C(n_1293),
.Y(n_1429)
);

NAND2x1p5_ASAP7_75t_L g1430 ( 
.A(n_1259),
.B(n_1387),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1276),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1278),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1285),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1291),
.Y(n_1434)
);

INVx5_ASAP7_75t_SL g1435 ( 
.A(n_1265),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1327),
.Y(n_1436)
);

BUFx12f_ASAP7_75t_L g1437 ( 
.A(n_1322),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1257),
.A2(n_1349),
.B1(n_1261),
.B2(n_1393),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1327),
.Y(n_1439)
);

CKINVDCx11_ASAP7_75t_R g1440 ( 
.A(n_1338),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1299),
.A2(n_1347),
.B(n_1348),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1317),
.A2(n_1320),
.B(n_1323),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1328),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1328),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1283),
.B(n_1361),
.Y(n_1445)
);

OR2x6_ASAP7_75t_L g1446 ( 
.A(n_1274),
.B(n_1265),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1277),
.A2(n_1292),
.B(n_1316),
.Y(n_1447)
);

NAND3xp33_ASAP7_75t_L g1448 ( 
.A(n_1384),
.B(n_1400),
.C(n_1383),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1406),
.B(n_1349),
.Y(n_1449)
);

OA21x2_ASAP7_75t_L g1450 ( 
.A1(n_1279),
.A2(n_1324),
.B(n_1326),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1259),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1380),
.B(n_1331),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1389),
.A2(n_1350),
.B1(n_1251),
.B2(n_1252),
.Y(n_1453)
);

AOI221xp5_ASAP7_75t_L g1454 ( 
.A1(n_1247),
.A2(n_1364),
.B1(n_1360),
.B2(n_1279),
.C(n_1284),
.Y(n_1454)
);

O2A1O1Ixp5_ASAP7_75t_L g1455 ( 
.A1(n_1393),
.A2(n_1381),
.B(n_1251),
.C(n_1345),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_1395),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1369),
.A2(n_1266),
.B(n_1326),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1319),
.A2(n_1330),
.B(n_1397),
.Y(n_1458)
);

INVx8_ASAP7_75t_L g1459 ( 
.A(n_1399),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1375),
.Y(n_1460)
);

OAI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1280),
.A2(n_1321),
.B(n_1346),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1312),
.A2(n_1311),
.B1(n_1358),
.B2(n_1262),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1256),
.A2(n_1267),
.B(n_1294),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1328),
.Y(n_1464)
);

INVx5_ASAP7_75t_L g1465 ( 
.A(n_1399),
.Y(n_1465)
);

OAI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1265),
.A2(n_1365),
.B1(n_1363),
.B2(n_1267),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1315),
.B(n_1302),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1330),
.A2(n_1373),
.B(n_1407),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1355),
.A2(n_1294),
.B(n_1288),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1392),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1288),
.A2(n_1256),
.B(n_1306),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1398),
.A2(n_1313),
.B(n_1396),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1366),
.B(n_1379),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1282),
.B(n_1334),
.C(n_1354),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1376),
.B(n_1318),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1308),
.A2(n_1329),
.B(n_1390),
.Y(n_1476)
);

INVxp67_ASAP7_75t_L g1477 ( 
.A(n_1351),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_1359),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1385),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1259),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1247),
.B(n_1406),
.Y(n_1481)
);

INVx2_ASAP7_75t_SL g1482 ( 
.A(n_1359),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1378),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1301),
.Y(n_1484)
);

AOI221xp5_ASAP7_75t_L g1485 ( 
.A1(n_1300),
.A2(n_1362),
.B1(n_1314),
.B2(n_1379),
.C(n_1325),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1308),
.A2(n_1304),
.B(n_1289),
.Y(n_1486)
);

O2A1O1Ixp33_ASAP7_75t_SL g1487 ( 
.A1(n_1332),
.A2(n_1333),
.B(n_1337),
.C(n_1343),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1335),
.B(n_1340),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1307),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1250),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1356),
.A2(n_1329),
.B(n_1408),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1333),
.Y(n_1492)
);

AO21x2_ASAP7_75t_L g1493 ( 
.A1(n_1263),
.A2(n_1304),
.B(n_1273),
.Y(n_1493)
);

INVx2_ASAP7_75t_SL g1494 ( 
.A(n_1403),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1356),
.A2(n_1337),
.B(n_1343),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1273),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1394),
.A2(n_1336),
.B1(n_1314),
.B2(n_1289),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1386),
.B(n_1253),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1275),
.B(n_1253),
.Y(n_1499)
);

BUFx10_ASAP7_75t_L g1500 ( 
.A(n_1399),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1372),
.A2(n_1368),
.B(n_1382),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1372),
.A2(n_1368),
.B(n_1382),
.Y(n_1502)
);

AOI21xp33_ASAP7_75t_L g1503 ( 
.A1(n_1263),
.A2(n_1394),
.B(n_1404),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1404),
.A2(n_1305),
.B(n_1352),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1401),
.Y(n_1505)
);

NAND3xp33_ASAP7_75t_L g1506 ( 
.A(n_1275),
.B(n_1387),
.C(n_1253),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1268),
.A2(n_1297),
.B(n_1248),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1268),
.A2(n_1297),
.B(n_1248),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_SL g1509 ( 
.A1(n_1342),
.A2(n_1401),
.B(n_1391),
.Y(n_1509)
);

OA21x2_ASAP7_75t_L g1510 ( 
.A1(n_1297),
.A2(n_1401),
.B(n_1370),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1370),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1370),
.A2(n_1371),
.B(n_1391),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_1403),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1298),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1388),
.A2(n_1342),
.B1(n_1352),
.B2(n_1391),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1342),
.A2(n_1352),
.B1(n_1298),
.B2(n_1371),
.Y(n_1516)
);

NAND3xp33_ASAP7_75t_L g1517 ( 
.A(n_1371),
.B(n_774),
.C(n_825),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1352),
.A2(n_1279),
.B(n_1271),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1367),
.A2(n_774),
.B1(n_630),
.B2(n_664),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1302),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_SL g1521 ( 
.A1(n_1264),
.A2(n_1252),
.B(n_1377),
.Y(n_1521)
);

BUFx2_ASAP7_75t_SL g1522 ( 
.A(n_1344),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1246),
.A2(n_1339),
.B(n_1271),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1246),
.A2(n_1339),
.B(n_1271),
.Y(n_1524)
);

CKINVDCx11_ASAP7_75t_R g1525 ( 
.A(n_1338),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1254),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1281),
.B(n_412),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1281),
.B(n_412),
.Y(n_1528)
);

AO21x2_ASAP7_75t_L g1529 ( 
.A1(n_1271),
.A2(n_1300),
.B(n_1260),
.Y(n_1529)
);

O2A1O1Ixp33_ASAP7_75t_SL g1530 ( 
.A1(n_1258),
.A2(n_1384),
.B(n_1383),
.C(n_1147),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1254),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1275),
.Y(n_1532)
);

NAND3xp33_ASAP7_75t_L g1533 ( 
.A(n_1258),
.B(n_774),
.C(n_825),
.Y(n_1533)
);

INVx2_ASAP7_75t_SL g1534 ( 
.A(n_1344),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1246),
.A2(n_1339),
.B(n_1271),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_SL g1536 ( 
.A1(n_1264),
.A2(n_1252),
.B(n_1377),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1309),
.Y(n_1537)
);

AO31x2_ASAP7_75t_L g1538 ( 
.A1(n_1271),
.A2(n_1147),
.A3(n_1156),
.B(n_1064),
.Y(n_1538)
);

OR2x6_ASAP7_75t_L g1539 ( 
.A(n_1274),
.B(n_1265),
.Y(n_1539)
);

NAND2x1p5_ASAP7_75t_L g1540 ( 
.A(n_1259),
.B(n_1387),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1246),
.A2(n_1339),
.B(n_1271),
.Y(n_1541)
);

AO21x2_ASAP7_75t_L g1542 ( 
.A1(n_1271),
.A2(n_1300),
.B(n_1260),
.Y(n_1542)
);

OAI221xp5_ASAP7_75t_L g1543 ( 
.A1(n_1290),
.A2(n_631),
.B1(n_614),
.B2(n_774),
.C(n_551),
.Y(n_1543)
);

OAI221xp5_ASAP7_75t_L g1544 ( 
.A1(n_1290),
.A2(n_631),
.B1(n_614),
.B2(n_774),
.C(n_551),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1290),
.A2(n_560),
.B1(n_574),
.B2(n_548),
.Y(n_1545)
);

OAI222xp33_ASAP7_75t_L g1546 ( 
.A1(n_1295),
.A2(n_664),
.B1(n_1094),
.B2(n_514),
.C1(n_516),
.C2(n_717),
.Y(n_1546)
);

AOI221xp5_ASAP7_75t_L g1547 ( 
.A1(n_1247),
.A2(n_630),
.B1(n_582),
.B2(n_774),
.C(n_649),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1309),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1254),
.Y(n_1549)
);

BUFx12f_ASAP7_75t_L g1550 ( 
.A(n_1322),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1249),
.B(n_990),
.Y(n_1551)
);

NAND2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1259),
.B(n_1387),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1246),
.A2(n_1339),
.B(n_1271),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1249),
.B(n_990),
.Y(n_1554)
);

NAND3xp33_ASAP7_75t_L g1555 ( 
.A(n_1258),
.B(n_774),
.C(n_825),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1344),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1302),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1338),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_SL g1559 ( 
.A1(n_1402),
.A2(n_551),
.B1(n_564),
.B2(n_517),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_SL g1560 ( 
.A1(n_1264),
.A2(n_1252),
.B(n_1377),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1246),
.A2(n_1339),
.B(n_1271),
.Y(n_1561)
);

OAI21xp33_ASAP7_75t_SL g1562 ( 
.A1(n_1252),
.A2(n_979),
.B(n_1046),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1271),
.A2(n_1064),
.B(n_986),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1246),
.A2(n_1339),
.B(n_1271),
.Y(n_1564)
);

O2A1O1Ixp33_ASAP7_75t_SL g1565 ( 
.A1(n_1258),
.A2(n_1384),
.B(n_1383),
.C(n_1147),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1249),
.B(n_990),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_SL g1567 ( 
.A1(n_1264),
.A2(n_1252),
.B(n_1377),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1331),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1309),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1246),
.A2(n_1339),
.B(n_1271),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1367),
.A2(n_774),
.B1(n_630),
.B2(n_664),
.Y(n_1571)
);

OA22x2_ASAP7_75t_L g1572 ( 
.A1(n_1418),
.A2(n_1413),
.B1(n_1509),
.B2(n_1462),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1410),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1559),
.A2(n_1429),
.B1(n_1422),
.B2(n_1519),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1551),
.B(n_1554),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1445),
.B(n_1475),
.Y(n_1576)
);

O2A1O1Ixp5_ASAP7_75t_L g1577 ( 
.A1(n_1426),
.A2(n_1546),
.B(n_1455),
.C(n_1461),
.Y(n_1577)
);

BUFx4f_ASAP7_75t_L g1578 ( 
.A(n_1437),
.Y(n_1578)
);

OA21x2_ASAP7_75t_L g1579 ( 
.A1(n_1457),
.A2(n_1508),
.B(n_1507),
.Y(n_1579)
);

AOI211xp5_ASAP7_75t_L g1580 ( 
.A1(n_1543),
.A2(n_1544),
.B(n_1533),
.C(n_1555),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1481),
.B(n_1452),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1422),
.A2(n_1519),
.B1(n_1571),
.B2(n_1438),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1563),
.A2(n_1424),
.B(n_1463),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1428),
.B(n_1473),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1417),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1562),
.A2(n_1486),
.B(n_1487),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1449),
.B(n_1415),
.Y(n_1587)
);

INVxp33_ASAP7_75t_L g1588 ( 
.A(n_1467),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1568),
.B(n_1488),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1419),
.Y(n_1590)
);

NOR2x1_ASAP7_75t_SL g1591 ( 
.A(n_1446),
.B(n_1539),
.Y(n_1591)
);

O2A1O1Ixp5_ASAP7_75t_L g1592 ( 
.A1(n_1503),
.A2(n_1453),
.B(n_1517),
.C(n_1448),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1527),
.B(n_1528),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1484),
.A2(n_1571),
.B1(n_1411),
.B2(n_1558),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1474),
.A2(n_1545),
.B1(n_1547),
.B2(n_1490),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1527),
.B(n_1528),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1446),
.A2(n_1539),
.B(n_1430),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1446),
.B(n_1539),
.Y(n_1598)
);

OA21x2_ASAP7_75t_L g1599 ( 
.A1(n_1457),
.A2(n_1541),
.B(n_1570),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1526),
.B(n_1531),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1416),
.B(n_1433),
.Y(n_1601)
);

O2A1O1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1530),
.A2(n_1565),
.B(n_1466),
.C(n_1454),
.Y(n_1602)
);

O2A1O1Ixp5_ASAP7_75t_L g1603 ( 
.A1(n_1466),
.A2(n_1511),
.B(n_1505),
.C(n_1444),
.Y(n_1603)
);

O2A1O1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1530),
.A2(n_1565),
.B(n_1487),
.C(n_1567),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1518),
.A2(n_1497),
.B(n_1469),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1515),
.A2(n_1477),
.B1(n_1478),
.B2(n_1497),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1518),
.A2(n_1469),
.B(n_1471),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1470),
.B(n_1460),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1549),
.B(n_1537),
.Y(n_1609)
);

OA21x2_ASAP7_75t_L g1610 ( 
.A1(n_1523),
.A2(n_1535),
.B(n_1564),
.Y(n_1610)
);

O2A1O1Ixp5_ASAP7_75t_L g1611 ( 
.A1(n_1443),
.A2(n_1464),
.B(n_1496),
.C(n_1489),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1478),
.A2(n_1435),
.B1(n_1557),
.B2(n_1520),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1548),
.B(n_1569),
.Y(n_1613)
);

A2O1A1Ixp33_ASAP7_75t_L g1614 ( 
.A1(n_1485),
.A2(n_1504),
.B(n_1468),
.C(n_1516),
.Y(n_1614)
);

AOI21x1_ASAP7_75t_SL g1615 ( 
.A1(n_1499),
.A2(n_1412),
.B(n_1538),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1514),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_SL g1617 ( 
.A1(n_1430),
.A2(n_1552),
.B(n_1540),
.Y(n_1617)
);

INVx3_ASAP7_75t_L g1618 ( 
.A(n_1500),
.Y(n_1618)
);

AND2x4_ASAP7_75t_SL g1619 ( 
.A(n_1456),
.B(n_1558),
.Y(n_1619)
);

OA21x2_ASAP7_75t_L g1620 ( 
.A1(n_1541),
.A2(n_1553),
.B(n_1564),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1548),
.B(n_1569),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1431),
.B(n_1432),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1506),
.B(n_1423),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1518),
.A2(n_1469),
.B(n_1471),
.Y(n_1624)
);

OA21x2_ASAP7_75t_L g1625 ( 
.A1(n_1553),
.A2(n_1561),
.B(n_1524),
.Y(n_1625)
);

AOI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1502),
.A2(n_1536),
.B1(n_1560),
.B2(n_1521),
.C(n_1427),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_SL g1627 ( 
.A1(n_1540),
.A2(n_1552),
.B(n_1451),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1434),
.B(n_1498),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1514),
.Y(n_1629)
);

A2O1A1Ixp33_ASAP7_75t_SL g1630 ( 
.A1(n_1516),
.A2(n_1532),
.B(n_1496),
.C(n_1492),
.Y(n_1630)
);

O2A1O1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1436),
.A2(n_1439),
.B(n_1479),
.C(n_1494),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1471),
.B(n_1436),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1423),
.A2(n_1465),
.B1(n_1483),
.B2(n_1522),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1412),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1451),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1480),
.B(n_1513),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1534),
.B(n_1556),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1420),
.B(n_1483),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1451),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1420),
.B(n_1451),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1501),
.B(n_1542),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1529),
.B(n_1542),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1423),
.A2(n_1465),
.B1(n_1459),
.B2(n_1484),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1412),
.B(n_1538),
.Y(n_1644)
);

AOI21x1_ASAP7_75t_SL g1645 ( 
.A1(n_1538),
.A2(n_1500),
.B(n_1425),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1472),
.B(n_1414),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1529),
.A2(n_1450),
.B(n_1458),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1538),
.B(n_1425),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1459),
.A2(n_1450),
.B1(n_1550),
.B2(n_1437),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1414),
.B(n_1476),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1500),
.B(n_1510),
.Y(n_1651)
);

AOI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1409),
.A2(n_1489),
.B1(n_1493),
.B2(n_1512),
.C(n_1510),
.Y(n_1652)
);

O2A1O1Ixp33_ASAP7_75t_L g1653 ( 
.A1(n_1409),
.A2(n_1493),
.B(n_1510),
.C(n_1512),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1491),
.Y(n_1654)
);

AOI21x1_ASAP7_75t_SL g1655 ( 
.A1(n_1512),
.A2(n_1495),
.B(n_1491),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_SL g1656 ( 
.A1(n_1550),
.A2(n_1440),
.B(n_1525),
.Y(n_1656)
);

OA21x2_ASAP7_75t_L g1657 ( 
.A1(n_1447),
.A2(n_1441),
.B(n_1442),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_SL g1658 ( 
.A1(n_1440),
.A2(n_1554),
.B(n_1551),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1525),
.A2(n_1559),
.B1(n_1429),
.B2(n_1422),
.Y(n_1659)
);

NAND2x1p5_ASAP7_75t_L g1660 ( 
.A(n_1423),
.B(n_1465),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1429),
.A2(n_1555),
.B1(n_1533),
.B2(n_1544),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1449),
.B(n_1446),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1551),
.B(n_1554),
.Y(n_1663)
);

NOR2xp67_ASAP7_75t_L g1664 ( 
.A(n_1482),
.B(n_1474),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1551),
.B(n_1554),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1420),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1559),
.A2(n_1429),
.B1(n_1422),
.B2(n_1519),
.Y(n_1667)
);

O2A1O1Ixp33_ASAP7_75t_L g1668 ( 
.A1(n_1543),
.A2(n_1544),
.B(n_1546),
.C(n_1530),
.Y(n_1668)
);

BUFx3_ASAP7_75t_L g1669 ( 
.A(n_1420),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1481),
.B(n_1452),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1481),
.B(n_1452),
.Y(n_1671)
);

O2A1O1Ixp33_ASAP7_75t_L g1672 ( 
.A1(n_1543),
.A2(n_1544),
.B(n_1546),
.C(n_1530),
.Y(n_1672)
);

CKINVDCx16_ASAP7_75t_R g1673 ( 
.A(n_1456),
.Y(n_1673)
);

O2A1O1Ixp33_ASAP7_75t_L g1674 ( 
.A1(n_1543),
.A2(n_1544),
.B(n_1546),
.C(n_1530),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1449),
.B(n_1446),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1445),
.B(n_1475),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1551),
.B(n_1554),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_SL g1678 ( 
.A1(n_1551),
.A2(n_1566),
.B(n_1554),
.Y(n_1678)
);

A2O1A1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1543),
.A2(n_1544),
.B(n_1555),
.C(n_1533),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_L g1680 ( 
.A1(n_1543),
.A2(n_1544),
.B(n_1546),
.C(n_1530),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1415),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1445),
.B(n_1475),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1445),
.B(n_1475),
.Y(n_1683)
);

OA21x2_ASAP7_75t_L g1684 ( 
.A1(n_1457),
.A2(n_1508),
.B(n_1507),
.Y(n_1684)
);

O2A1O1Ixp33_ASAP7_75t_L g1685 ( 
.A1(n_1543),
.A2(n_1544),
.B(n_1546),
.C(n_1530),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_SL g1686 ( 
.A1(n_1551),
.A2(n_1566),
.B(n_1554),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1445),
.B(n_1475),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1551),
.B(n_1554),
.Y(n_1688)
);

NOR2x1_ASAP7_75t_SL g1689 ( 
.A(n_1446),
.B(n_1539),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1551),
.B(n_1554),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1551),
.B(n_1554),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1563),
.A2(n_1064),
.B(n_1461),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1563),
.A2(n_1064),
.B(n_1461),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1421),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1445),
.B(n_1475),
.Y(n_1695)
);

O2A1O1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1543),
.A2(n_1544),
.B(n_1546),
.C(n_1530),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_1440),
.Y(n_1697)
);

OR2x6_ASAP7_75t_L g1698 ( 
.A(n_1597),
.B(n_1586),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1632),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1573),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1598),
.B(n_1591),
.Y(n_1701)
);

INVx3_ASAP7_75t_L g1702 ( 
.A(n_1650),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1585),
.Y(n_1703)
);

BUFx2_ASAP7_75t_L g1704 ( 
.A(n_1651),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1581),
.B(n_1670),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1611),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1681),
.Y(n_1707)
);

OAI21x1_ASAP7_75t_L g1708 ( 
.A1(n_1655),
.A2(n_1647),
.B(n_1624),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1590),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1598),
.Y(n_1710)
);

OAI21x1_ASAP7_75t_SL g1711 ( 
.A1(n_1689),
.A2(n_1602),
.B(n_1631),
.Y(n_1711)
);

OAI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1577),
.A2(n_1679),
.B(n_1592),
.Y(n_1712)
);

OA21x2_ASAP7_75t_L g1713 ( 
.A1(n_1607),
.A2(n_1605),
.B(n_1586),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1694),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1642),
.B(n_1641),
.Y(n_1715)
);

CKINVDCx20_ASAP7_75t_R g1716 ( 
.A(n_1673),
.Y(n_1716)
);

OR2x6_ASAP7_75t_L g1717 ( 
.A(n_1692),
.B(n_1693),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1644),
.B(n_1648),
.Y(n_1718)
);

AOI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1583),
.A2(n_1693),
.B(n_1692),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1694),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1579),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1582),
.A2(n_1661),
.B1(n_1667),
.B2(n_1574),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1634),
.Y(n_1723)
);

AO21x2_ASAP7_75t_L g1724 ( 
.A1(n_1630),
.A2(n_1653),
.B(n_1614),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1671),
.B(n_1584),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1576),
.B(n_1676),
.Y(n_1726)
);

AO21x2_ASAP7_75t_L g1727 ( 
.A1(n_1653),
.A2(n_1654),
.B(n_1650),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1684),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1646),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1646),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1600),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1609),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1613),
.Y(n_1733)
);

AOI221xp5_ASAP7_75t_L g1734 ( 
.A1(n_1668),
.A2(n_1685),
.B1(n_1696),
.B2(n_1672),
.C(n_1674),
.Y(n_1734)
);

OR2x6_ASAP7_75t_L g1735 ( 
.A(n_1660),
.B(n_1602),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1657),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1575),
.B(n_1663),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1665),
.B(n_1677),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1682),
.B(n_1683),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1628),
.B(n_1608),
.Y(n_1740)
);

OR2x6_ASAP7_75t_L g1741 ( 
.A(n_1604),
.B(n_1662),
.Y(n_1741)
);

INVxp67_ASAP7_75t_SL g1742 ( 
.A(n_1631),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1687),
.B(n_1695),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1688),
.B(n_1690),
.Y(n_1744)
);

OA21x2_ASAP7_75t_L g1745 ( 
.A1(n_1652),
.A2(n_1603),
.B(n_1592),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1659),
.A2(n_1572),
.B1(n_1594),
.B2(n_1595),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1572),
.B(n_1587),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1599),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1621),
.B(n_1622),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1603),
.B(n_1675),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1601),
.Y(n_1751)
);

CKINVDCx14_ASAP7_75t_R g1752 ( 
.A(n_1697),
.Y(n_1752)
);

OR2x6_ASAP7_75t_L g1753 ( 
.A(n_1604),
.B(n_1675),
.Y(n_1753)
);

AO21x2_ASAP7_75t_L g1754 ( 
.A1(n_1668),
.A2(n_1674),
.B(n_1696),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1577),
.Y(n_1755)
);

INVxp67_ASAP7_75t_SL g1756 ( 
.A(n_1589),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1623),
.Y(n_1757)
);

AO21x2_ASAP7_75t_L g1758 ( 
.A1(n_1672),
.A2(n_1680),
.B(n_1685),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1588),
.B(n_1593),
.Y(n_1759)
);

OA21x2_ASAP7_75t_L g1760 ( 
.A1(n_1626),
.A2(n_1645),
.B(n_1606),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_SL g1761 ( 
.A(n_1643),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1700),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1700),
.Y(n_1763)
);

INVxp67_ASAP7_75t_L g1764 ( 
.A(n_1742),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1703),
.Y(n_1765)
);

AOI221xp5_ASAP7_75t_L g1766 ( 
.A1(n_1722),
.A2(n_1680),
.B1(n_1580),
.B2(n_1686),
.C(n_1678),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1715),
.B(n_1625),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1715),
.B(n_1625),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1704),
.B(n_1620),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1703),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1746),
.A2(n_1722),
.B1(n_1734),
.B2(n_1712),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1699),
.B(n_1691),
.Y(n_1772)
);

BUFx6f_ASAP7_75t_L g1773 ( 
.A(n_1698),
.Y(n_1773)
);

OR2x6_ASAP7_75t_L g1774 ( 
.A(n_1698),
.B(n_1617),
.Y(n_1774)
);

NAND2x1_ASAP7_75t_L g1775 ( 
.A(n_1698),
.B(n_1627),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1709),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1699),
.B(n_1664),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1750),
.B(n_1610),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1755),
.B(n_1596),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1718),
.B(n_1649),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1717),
.B(n_1640),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1714),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1718),
.B(n_1612),
.Y(n_1783)
);

BUFx3_ASAP7_75t_L g1784 ( 
.A(n_1714),
.Y(n_1784)
);

INVxp67_ASAP7_75t_SL g1785 ( 
.A(n_1706),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1717),
.B(n_1615),
.Y(n_1786)
);

NOR2x1_ASAP7_75t_L g1787 ( 
.A(n_1698),
.B(n_1658),
.Y(n_1787)
);

AOI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1734),
.A2(n_1754),
.B1(n_1758),
.B2(n_1712),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1750),
.B(n_1629),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1725),
.B(n_1720),
.Y(n_1790)
);

INVxp67_ASAP7_75t_L g1791 ( 
.A(n_1707),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1720),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1754),
.A2(n_1578),
.B1(n_1669),
.B2(n_1633),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1723),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1747),
.B(n_1616),
.Y(n_1795)
);

OAI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1737),
.A2(n_1638),
.B1(n_1578),
.B2(n_1619),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1747),
.B(n_1702),
.Y(n_1797)
);

NOR2x1p5_ASAP7_75t_L g1798 ( 
.A(n_1710),
.B(n_1618),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1749),
.B(n_1635),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1725),
.B(n_1639),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1705),
.B(n_1731),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1723),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1797),
.B(n_1729),
.Y(n_1803)
);

BUFx3_ASAP7_75t_L g1804 ( 
.A(n_1784),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1766),
.A2(n_1758),
.B1(n_1754),
.B2(n_1717),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1790),
.B(n_1801),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1797),
.B(n_1729),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1789),
.B(n_1778),
.Y(n_1808)
);

OA21x2_ASAP7_75t_L g1809 ( 
.A1(n_1785),
.A2(n_1708),
.B(n_1728),
.Y(n_1809)
);

INVx4_ASAP7_75t_L g1810 ( 
.A(n_1774),
.Y(n_1810)
);

OAI33xp33_ASAP7_75t_L g1811 ( 
.A1(n_1771),
.A2(n_1755),
.A3(n_1705),
.B1(n_1738),
.B2(n_1737),
.B3(n_1744),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1788),
.A2(n_1761),
.B1(n_1735),
.B2(n_1753),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1789),
.B(n_1729),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1794),
.Y(n_1814)
);

OAI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1766),
.A2(n_1717),
.B1(n_1744),
.B2(n_1738),
.C(n_1698),
.Y(n_1815)
);

OAI211xp5_ASAP7_75t_L g1816 ( 
.A1(n_1771),
.A2(n_1745),
.B(n_1760),
.C(n_1751),
.Y(n_1816)
);

AOI31xp33_ASAP7_75t_L g1817 ( 
.A1(n_1787),
.A2(n_1752),
.A3(n_1701),
.B(n_1756),
.Y(n_1817)
);

AO221x1_ASAP7_75t_L g1818 ( 
.A1(n_1796),
.A2(n_1711),
.B1(n_1757),
.B2(n_1751),
.C(n_1730),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1793),
.A2(n_1761),
.B1(n_1735),
.B2(n_1741),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1790),
.B(n_1731),
.Y(n_1820)
);

NAND2xp33_ASAP7_75t_R g1821 ( 
.A(n_1777),
.B(n_1759),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_1800),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1779),
.B(n_1740),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1787),
.A2(n_1758),
.B1(n_1754),
.B2(n_1717),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1794),
.Y(n_1825)
);

AOI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1796),
.A2(n_1758),
.B1(n_1735),
.B2(n_1701),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1778),
.B(n_1781),
.Y(n_1827)
);

AOI21x1_ASAP7_75t_L g1828 ( 
.A1(n_1775),
.A2(n_1748),
.B(n_1736),
.Y(n_1828)
);

INVx5_ASAP7_75t_SL g1829 ( 
.A(n_1774),
.Y(n_1829)
);

OAI211xp5_ASAP7_75t_L g1830 ( 
.A1(n_1764),
.A2(n_1745),
.B(n_1760),
.C(n_1719),
.Y(n_1830)
);

NAND2xp33_ASAP7_75t_R g1831 ( 
.A(n_1777),
.B(n_1759),
.Y(n_1831)
);

INVxp67_ASAP7_75t_L g1832 ( 
.A(n_1779),
.Y(n_1832)
);

AOI221xp5_ASAP7_75t_L g1833 ( 
.A1(n_1764),
.A2(n_1732),
.B1(n_1726),
.B2(n_1739),
.C(n_1743),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1802),
.Y(n_1834)
);

OAI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1774),
.A2(n_1735),
.B1(n_1741),
.B2(n_1753),
.Y(n_1835)
);

BUFx2_ASAP7_75t_L g1836 ( 
.A(n_1784),
.Y(n_1836)
);

OAI221xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1780),
.A2(n_1735),
.B1(n_1753),
.B2(n_1741),
.C(n_1656),
.Y(n_1837)
);

NAND2xp33_ASAP7_75t_R g1838 ( 
.A(n_1772),
.B(n_1760),
.Y(n_1838)
);

INVx1_ASAP7_75t_SL g1839 ( 
.A(n_1800),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1781),
.B(n_1767),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1802),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1801),
.B(n_1727),
.Y(n_1842)
);

AOI221xp5_ASAP7_75t_L g1843 ( 
.A1(n_1791),
.A2(n_1732),
.B1(n_1739),
.B2(n_1726),
.C(n_1743),
.Y(n_1843)
);

AOI222xp33_ASAP7_75t_L g1844 ( 
.A1(n_1791),
.A2(n_1711),
.B1(n_1772),
.B2(n_1716),
.C1(n_1786),
.C2(n_1733),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1792),
.Y(n_1845)
);

INVxp67_ASAP7_75t_L g1846 ( 
.A(n_1799),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1781),
.B(n_1730),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1827),
.B(n_1840),
.Y(n_1848)
);

OAI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1805),
.A2(n_1745),
.B(n_1760),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1814),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1814),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1809),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1825),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1827),
.B(n_1767),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1825),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1834),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1817),
.B(n_1773),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1834),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1844),
.B(n_1773),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1841),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1832),
.B(n_1792),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1841),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1845),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1840),
.B(n_1768),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1808),
.B(n_1768),
.Y(n_1865)
);

BUFx3_ASAP7_75t_L g1866 ( 
.A(n_1836),
.Y(n_1866)
);

NOR2x1_ASAP7_75t_SL g1867 ( 
.A(n_1816),
.B(n_1774),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1811),
.B(n_1823),
.Y(n_1868)
);

INVx5_ASAP7_75t_L g1869 ( 
.A(n_1829),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1808),
.B(n_1786),
.Y(n_1870)
);

BUFx2_ASAP7_75t_L g1871 ( 
.A(n_1810),
.Y(n_1871)
);

INVx4_ASAP7_75t_SL g1872 ( 
.A(n_1804),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1845),
.Y(n_1873)
);

NAND2x1p5_ASAP7_75t_SL g1874 ( 
.A(n_1837),
.B(n_1786),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1826),
.B(n_1773),
.Y(n_1875)
);

OA21x2_ASAP7_75t_L g1876 ( 
.A1(n_1830),
.A2(n_1721),
.B(n_1728),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1828),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1847),
.B(n_1769),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1842),
.B(n_1782),
.Y(n_1879)
);

NOR2x1p5_ASAP7_75t_L g1880 ( 
.A(n_1810),
.B(n_1775),
.Y(n_1880)
);

INVx4_ASAP7_75t_SL g1881 ( 
.A(n_1804),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1868),
.B(n_1833),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1853),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1866),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1868),
.B(n_1843),
.Y(n_1885)
);

NAND2x1p5_ASAP7_75t_L g1886 ( 
.A(n_1869),
.B(n_1810),
.Y(n_1886)
);

NAND4xp75_ASAP7_75t_L g1887 ( 
.A(n_1859),
.B(n_1745),
.C(n_1636),
.D(n_1713),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1859),
.A2(n_1812),
.B1(n_1815),
.B2(n_1819),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1870),
.B(n_1848),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1870),
.B(n_1848),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1853),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1853),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1870),
.B(n_1847),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1848),
.B(n_1813),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1861),
.B(n_1795),
.Y(n_1895)
);

HB1xp67_ASAP7_75t_L g1896 ( 
.A(n_1866),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1855),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1861),
.B(n_1795),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1871),
.B(n_1637),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1877),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1871),
.B(n_1822),
.Y(n_1901)
);

INVx4_ASAP7_75t_L g1902 ( 
.A(n_1869),
.Y(n_1902)
);

AOI22xp5_ASAP7_75t_L g1903 ( 
.A1(n_1849),
.A2(n_1838),
.B1(n_1824),
.B2(n_1724),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1872),
.B(n_1813),
.Y(n_1904)
);

OAI322xp33_ASAP7_75t_L g1905 ( 
.A1(n_1875),
.A2(n_1842),
.A3(n_1821),
.B1(n_1831),
.B2(n_1783),
.C1(n_1780),
.C2(n_1806),
.Y(n_1905)
);

A2O1A1Ixp33_ASAP7_75t_L g1906 ( 
.A1(n_1857),
.A2(n_1783),
.B(n_1773),
.C(n_1701),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1871),
.B(n_1839),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1855),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1855),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1875),
.B(n_1806),
.Y(n_1910)
);

AOI221xp5_ASAP7_75t_L g1911 ( 
.A1(n_1849),
.A2(n_1818),
.B1(n_1835),
.B2(n_1846),
.C(n_1836),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1872),
.B(n_1803),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1878),
.B(n_1820),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1858),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1852),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1878),
.B(n_1820),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1858),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1872),
.B(n_1803),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1872),
.B(n_1807),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1878),
.B(n_1807),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1872),
.B(n_1818),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1852),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1869),
.B(n_1773),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1880),
.B(n_1798),
.Y(n_1924)
);

OAI33xp33_ASAP7_75t_L g1925 ( 
.A1(n_1858),
.A2(n_1770),
.A3(n_1765),
.B1(n_1763),
.B2(n_1762),
.B3(n_1776),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1879),
.B(n_1782),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1863),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1883),
.Y(n_1928)
);

INVx3_ASAP7_75t_SL g1929 ( 
.A(n_1902),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1885),
.B(n_1854),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1889),
.Y(n_1931)
);

NOR2x1p5_ASAP7_75t_SL g1932 ( 
.A(n_1887),
.B(n_1852),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1882),
.B(n_1854),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1924),
.B(n_1921),
.Y(n_1934)
);

AOI222xp33_ASAP7_75t_L g1935 ( 
.A1(n_1888),
.A2(n_1867),
.B1(n_1857),
.B2(n_1881),
.C1(n_1872),
.C2(n_1866),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1884),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1889),
.Y(n_1937)
);

INVxp67_ASAP7_75t_L g1938 ( 
.A(n_1899),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1883),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1924),
.B(n_1872),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1891),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1924),
.B(n_1881),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1924),
.B(n_1881),
.Y(n_1943)
);

AOI211xp5_ASAP7_75t_L g1944 ( 
.A1(n_1905),
.A2(n_1874),
.B(n_1866),
.C(n_1867),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1903),
.B(n_1854),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1891),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1903),
.B(n_1864),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1901),
.B(n_1864),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1890),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1905),
.B(n_1666),
.Y(n_1950)
);

AOI21xp33_ASAP7_75t_L g1951 ( 
.A1(n_1923),
.A2(n_1869),
.B(n_1876),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1892),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1892),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1890),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1910),
.B(n_1879),
.Y(n_1955)
);

OR2x2_ASAP7_75t_L g1956 ( 
.A(n_1913),
.B(n_1879),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1907),
.B(n_1864),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1896),
.B(n_1865),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1897),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1895),
.B(n_1898),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1916),
.B(n_1863),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1926),
.B(n_1863),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1921),
.B(n_1881),
.Y(n_1963)
);

NAND3xp33_ASAP7_75t_L g1964 ( 
.A(n_1911),
.B(n_1869),
.C(n_1876),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1936),
.Y(n_1965)
);

BUFx3_ASAP7_75t_L g1966 ( 
.A(n_1936),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1928),
.Y(n_1967)
);

INVx1_ASAP7_75t_SL g1968 ( 
.A(n_1940),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1928),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1931),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1939),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1938),
.B(n_1894),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1930),
.B(n_1894),
.Y(n_1973)
);

INVx1_ASAP7_75t_SL g1974 ( 
.A(n_1940),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1931),
.Y(n_1975)
);

OR2x6_ASAP7_75t_L g1976 ( 
.A(n_1932),
.B(n_1902),
.Y(n_1976)
);

INVx2_ASAP7_75t_SL g1977 ( 
.A(n_1929),
.Y(n_1977)
);

OAI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1944),
.A2(n_1887),
.B1(n_1906),
.B2(n_1869),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1937),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1933),
.B(n_1893),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1939),
.Y(n_1981)
);

INVx1_ASAP7_75t_SL g1982 ( 
.A(n_1942),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1950),
.B(n_1902),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1937),
.Y(n_1984)
);

INVx1_ASAP7_75t_SL g1985 ( 
.A(n_1942),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1941),
.Y(n_1986)
);

INVxp67_ASAP7_75t_L g1987 ( 
.A(n_1934),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1964),
.A2(n_1869),
.B1(n_1886),
.B2(n_1902),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1960),
.B(n_1893),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1941),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1946),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1946),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1949),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1966),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1987),
.B(n_1934),
.Y(n_1995)
);

AOI21xp5_ASAP7_75t_L g1996 ( 
.A1(n_1978),
.A2(n_1935),
.B(n_1951),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1966),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1988),
.A2(n_1947),
.B(n_1945),
.Y(n_1998)
);

OA21x2_ASAP7_75t_L g1999 ( 
.A1(n_1965),
.A2(n_1969),
.B(n_1967),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1968),
.B(n_1949),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1976),
.Y(n_2001)
);

O2A1O1Ixp33_ASAP7_75t_L g2002 ( 
.A1(n_1976),
.A2(n_1929),
.B(n_1932),
.C(n_1886),
.Y(n_2002)
);

OAI221xp5_ASAP7_75t_SL g2003 ( 
.A1(n_1976),
.A2(n_1943),
.B1(n_1954),
.B2(n_1955),
.C(n_1963),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1967),
.Y(n_2004)
);

OAI221xp5_ASAP7_75t_L g2005 ( 
.A1(n_1983),
.A2(n_1886),
.B1(n_1943),
.B2(n_1963),
.C(n_1958),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1974),
.B(n_1954),
.Y(n_2006)
);

AOI31xp33_ASAP7_75t_L g2007 ( 
.A1(n_1977),
.A2(n_1982),
.A3(n_1985),
.B(n_1972),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1969),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1971),
.Y(n_2009)
);

AOI211xp5_ASAP7_75t_SL g2010 ( 
.A1(n_1970),
.A2(n_1955),
.B(n_1959),
.C(n_1953),
.Y(n_2010)
);

NAND2xp33_ASAP7_75t_L g2011 ( 
.A(n_1977),
.B(n_1880),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1989),
.B(n_1948),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1971),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1999),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1995),
.B(n_1997),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1995),
.B(n_1970),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1999),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1994),
.B(n_1973),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1999),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1997),
.Y(n_2020)
);

HB1xp67_ASAP7_75t_L g2021 ( 
.A(n_2010),
.Y(n_2021)
);

INVx1_ASAP7_75t_SL g2022 ( 
.A(n_2000),
.Y(n_2022)
);

OAI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_2007),
.A2(n_1976),
.B1(n_1980),
.B2(n_1957),
.Y(n_2023)
);

NAND3x1_ASAP7_75t_L g2024 ( 
.A(n_2004),
.B(n_2009),
.C(n_2008),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2013),
.Y(n_2025)
);

AOI322xp5_ASAP7_75t_L g2026 ( 
.A1(n_2021),
.A2(n_2012),
.A3(n_2006),
.B1(n_2011),
.B2(n_2001),
.C1(n_1991),
.C2(n_1990),
.Y(n_2026)
);

AOI21xp33_ASAP7_75t_L g2027 ( 
.A1(n_2021),
.A2(n_2002),
.B(n_2001),
.Y(n_2027)
);

NAND4xp75_ASAP7_75t_L g2028 ( 
.A(n_2017),
.B(n_1996),
.C(n_1998),
.D(n_1979),
.Y(n_2028)
);

OAI211xp5_ASAP7_75t_L g2029 ( 
.A1(n_2014),
.A2(n_2003),
.B(n_2005),
.C(n_1979),
.Y(n_2029)
);

OAI321xp33_ASAP7_75t_L g2030 ( 
.A1(n_2023),
.A2(n_1984),
.A3(n_1993),
.B1(n_1975),
.B2(n_1990),
.C(n_1992),
.Y(n_2030)
);

NOR2x1_ASAP7_75t_L g2031 ( 
.A(n_2014),
.B(n_1981),
.Y(n_2031)
);

O2A1O1Ixp33_ASAP7_75t_L g2032 ( 
.A1(n_2019),
.A2(n_2011),
.B(n_1992),
.C(n_1986),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_2022),
.B(n_1975),
.Y(n_2033)
);

OAI21xp33_ASAP7_75t_L g2034 ( 
.A1(n_2018),
.A2(n_1993),
.B(n_1984),
.Y(n_2034)
);

OAI22xp33_ASAP7_75t_L g2035 ( 
.A1(n_2019),
.A2(n_2015),
.B1(n_2016),
.B2(n_2020),
.Y(n_2035)
);

AOI211xp5_ASAP7_75t_L g2036 ( 
.A1(n_2025),
.A2(n_1986),
.B(n_1981),
.C(n_2024),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_2026),
.B(n_1961),
.Y(n_2037)
);

INVx1_ASAP7_75t_SL g2038 ( 
.A(n_2033),
.Y(n_2038)
);

AOI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_2028),
.A2(n_1912),
.B1(n_1919),
.B2(n_1918),
.Y(n_2039)
);

AOI221xp5_ASAP7_75t_L g2040 ( 
.A1(n_2035),
.A2(n_1952),
.B1(n_1953),
.B2(n_1874),
.C(n_1900),
.Y(n_2040)
);

AOI221xp5_ASAP7_75t_L g2041 ( 
.A1(n_2027),
.A2(n_1952),
.B1(n_1874),
.B2(n_1900),
.C(n_1925),
.Y(n_2041)
);

AOI32xp33_ASAP7_75t_L g2042 ( 
.A1(n_2030),
.A2(n_1904),
.A3(n_1912),
.B1(n_1918),
.B2(n_1919),
.Y(n_2042)
);

AOI31xp33_ASAP7_75t_L g2043 ( 
.A1(n_2036),
.A2(n_1956),
.A3(n_1961),
.B(n_1962),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2038),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_2039),
.B(n_2034),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_2037),
.B(n_2029),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2043),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2040),
.Y(n_2048)
);

INVxp67_ASAP7_75t_SL g2049 ( 
.A(n_2041),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_2042),
.B(n_2031),
.Y(n_2050)
);

AOI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_2046),
.A2(n_1904),
.B1(n_1881),
.B2(n_1956),
.Y(n_2051)
);

AOI322xp5_ASAP7_75t_L g2052 ( 
.A1(n_2049),
.A2(n_2032),
.A3(n_1915),
.B1(n_1922),
.B2(n_1927),
.C1(n_1897),
.C2(n_1917),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_2044),
.Y(n_2053)
);

OR2x2_ASAP7_75t_L g2054 ( 
.A(n_2047),
.B(n_1962),
.Y(n_2054)
);

OAI221xp5_ASAP7_75t_SL g2055 ( 
.A1(n_2048),
.A2(n_1922),
.B1(n_1915),
.B2(n_1926),
.C(n_1908),
.Y(n_2055)
);

INVxp67_ASAP7_75t_SL g2056 ( 
.A(n_2050),
.Y(n_2056)
);

AOI221xp5_ASAP7_75t_SL g2057 ( 
.A1(n_2056),
.A2(n_2050),
.B1(n_2045),
.B2(n_1915),
.C(n_1922),
.Y(n_2057)
);

AOI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_2053),
.A2(n_2045),
.B1(n_1881),
.B2(n_1914),
.Y(n_2058)
);

NOR2xp67_ASAP7_75t_L g2059 ( 
.A(n_2054),
.B(n_1908),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_2058),
.B(n_2051),
.Y(n_2060)
);

AOI322xp5_ASAP7_75t_L g2061 ( 
.A1(n_2060),
.A2(n_2057),
.A3(n_2055),
.B1(n_2059),
.B2(n_2052),
.C1(n_1877),
.C2(n_1927),
.Y(n_2061)
);

XNOR2x1_ASAP7_75t_L g2062 ( 
.A(n_2061),
.B(n_1666),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2061),
.Y(n_2063)
);

INVxp67_ASAP7_75t_L g2064 ( 
.A(n_2063),
.Y(n_2064)
);

OA21x2_ASAP7_75t_L g2065 ( 
.A1(n_2062),
.A2(n_1914),
.B(n_1909),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_2065),
.Y(n_2066)
);

AND2x4_ASAP7_75t_SL g2067 ( 
.A(n_2064),
.B(n_1666),
.Y(n_2067)
);

AOI22xp33_ASAP7_75t_R g2068 ( 
.A1(n_2066),
.A2(n_1860),
.B1(n_1856),
.B2(n_1851),
.Y(n_2068)
);

AOI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_2068),
.A2(n_2067),
.B(n_1917),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_2069),
.A2(n_1909),
.B(n_1920),
.Y(n_2070)
);

AO221x1_ASAP7_75t_L g2071 ( 
.A1(n_2070),
.A2(n_1874),
.B1(n_1877),
.B2(n_1850),
.C(n_1862),
.Y(n_2071)
);

AOI22xp5_ASAP7_75t_L g2072 ( 
.A1(n_2071),
.A2(n_1881),
.B1(n_1856),
.B2(n_1860),
.Y(n_2072)
);

OA22x2_ASAP7_75t_L g2073 ( 
.A1(n_2072),
.A2(n_1851),
.B1(n_1877),
.B2(n_1873),
.Y(n_2073)
);


endmodule