module fake_jpeg_12285_n_158 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_158);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_L g32 ( 
.A1(n_13),
.A2(n_0),
.B(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_32),
.B(n_35),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_12),
.B(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_38),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_23),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_37)
);

AO21x1_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_47),
.B(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_12),
.B(n_10),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_40),
.B(n_17),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_50),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g44 ( 
.A1(n_21),
.A2(n_2),
.B(n_4),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_13),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_4),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_6),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_6),
.B1(n_29),
.B2(n_27),
.Y(n_47)
);

AO22x1_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_15),
.B1(n_24),
.B2(n_16),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_72),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_59),
.B(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_25),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_17),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_76),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx24_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_74),
.B1(n_60),
.B2(n_79),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_88),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_24),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_82),
.B(n_91),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_18),
.B(n_26),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_60),
.B(n_75),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_18),
.B1(n_26),
.B2(n_45),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_87),
.B1(n_89),
.B2(n_94),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_27),
.B1(n_19),
.B2(n_33),
.Y(n_87)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_22),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_22),
.B1(n_67),
.B2(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_22),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_65),
.B1(n_70),
.B2(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_52),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_98),
.Y(n_107)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_109),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_108),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_64),
.B(n_68),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_111),
.Y(n_123)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_91),
.B(n_63),
.Y(n_113)
);

NOR2xp67_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_116),
.Y(n_118)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_95),
.C(n_97),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_120),
.C(n_125),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_95),
.C(n_97),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_95),
.C(n_81),
.Y(n_125)
);

AOI211xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_88),
.B(n_83),
.C(n_81),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_127),
.B(n_89),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_107),
.B(n_98),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_132),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_115),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_125),
.C(n_121),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_115),
.B1(n_114),
.B2(n_105),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_109),
.B(n_86),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_133),
.A2(n_123),
.B1(n_122),
.B2(n_124),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_120),
.A2(n_100),
.B(n_102),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_134),
.B(n_137),
.Y(n_139)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_130),
.C(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_129),
.B(n_133),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_146),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_130),
.C(n_131),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_147),
.A2(n_148),
.B(n_143),
.Y(n_151)
);

BUFx12f_ASAP7_75t_SL g148 ( 
.A(n_141),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_151),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_147),
.C(n_143),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_75),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_152),
.A2(n_140),
.B(n_142),
.C(n_124),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_155),
.C(n_90),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_90),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_64),
.Y(n_158)
);


endmodule