module fake_jpeg_17824_n_46 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_46);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_8),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_0),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_7),
.B(n_6),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_SL g30 ( 
.A1(n_19),
.A2(n_20),
.B(n_24),
.C(n_17),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_1),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_18),
.A2(n_3),
.B1(n_21),
.B2(n_28),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_19),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_21),
.B1(n_25),
.B2(n_16),
.Y(n_37)
);

AOI322xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_30),
.A3(n_29),
.B1(n_37),
.B2(n_24),
.C1(n_15),
.C2(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_37),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_30),
.B1(n_34),
.B2(n_27),
.Y(n_42)
);

AOI322xp5_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_43),
.A3(n_22),
.B1(n_31),
.B2(n_36),
.C1(n_39),
.C2(n_41),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_43),
.B(n_22),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_22),
.Y(n_46)
);


endmodule