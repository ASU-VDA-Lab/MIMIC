module fake_jpeg_10170_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_38),
.Y(n_48)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_2),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_1),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_20),
.Y(n_51)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_23),
.B1(n_19),
.B2(n_33),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_53),
.B1(n_60),
.B2(n_16),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_62),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_19),
.B1(n_23),
.B2(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_30),
.B1(n_28),
.B2(n_27),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_24),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_30),
.B1(n_32),
.B2(n_26),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_2),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_66),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_37),
.B(n_24),
.Y(n_64)
);

BUFx24_ASAP7_75t_SL g81 ( 
.A(n_64),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_18),
.B1(n_26),
.B2(n_22),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_67),
.Y(n_91)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_71),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_86),
.Y(n_100)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_79),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_55),
.B(n_16),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_84),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_8),
.C(n_15),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_80),
.B(n_63),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_2),
.Y(n_84)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_3),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_48),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_77),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_54),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_98),
.B(n_104),
.Y(n_127)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_83),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_63),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_58),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_47),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_110),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_56),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_84),
.C(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_47),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_78),
.C(n_87),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_118),
.C(n_120),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_114),
.B(n_119),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_121),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_74),
.C(n_69),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_84),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_75),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_124),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_83),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_69),
.B1(n_72),
.B2(n_82),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_82),
.B1(n_127),
.B2(n_116),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_100),
.B(n_107),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_139),
.B1(n_65),
.B2(n_17),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_95),
.Y(n_130)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_126),
.A2(n_102),
.B1(n_106),
.B2(n_107),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_132),
.A2(n_138),
.B1(n_111),
.B2(n_93),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_110),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_135),
.B(n_112),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_98),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_94),
.B(n_22),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_115),
.B(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_56),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_141),
.B1(n_112),
.B2(n_65),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_93),
.B(n_26),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_52),
.B(n_59),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_138),
.B1(n_141),
.B2(n_137),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_144),
.A2(n_129),
.B1(n_142),
.B2(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_151),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_146),
.B(n_22),
.CI(n_52),
.CON(n_157),
.SN(n_157)
);

NOR3xp33_ASAP7_75t_SL g158 ( 
.A(n_148),
.B(n_3),
.C(n_4),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_59),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_152),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_15),
.C2(n_151),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

BUFx12_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_155),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_144),
.A2(n_135),
.B1(n_119),
.B2(n_52),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_149),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_159),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_153),
.C(n_147),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_163),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_146),
.C(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_167),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_152),
.C(n_5),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_165),
.Y(n_168)
);

OAI211xp5_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_171),
.B(n_172),
.C(n_157),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_155),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_158),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_175),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_171),
.A2(n_156),
.B(n_157),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_170),
.B(n_4),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_159),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_177),
.Y(n_179)
);


endmodule