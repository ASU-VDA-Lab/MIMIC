module real_jpeg_21236_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_328, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_328;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx13_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_0),
.A2(n_42),
.B1(n_43),
.B2(n_53),
.Y(n_55)
);

OAI32xp33_ASAP7_75t_L g186 ( 
.A1(n_0),
.A2(n_32),
.A3(n_43),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_1),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_65),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_65),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_65),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_62),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_62),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_62),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_3),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_104),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_104),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_104),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_4),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_97),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_97),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_97),
.Y(n_177)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_6),
.Y(n_82)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_6),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_7),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_7),
.B(n_30),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_7),
.A2(n_14),
.B(n_46),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_102),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_7),
.A2(n_81),
.B1(n_82),
.B2(n_160),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_7),
.B(n_57),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g191 ( 
.A1(n_7),
.A2(n_32),
.B(n_192),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_9),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_93),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_93),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_93),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_10),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_99),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_99),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_99),
.Y(n_238)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_12),
.A2(n_35),
.B1(n_42),
.B2(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_12),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_13),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_87),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_87),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_87),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_14),
.Y(n_44)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_14),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_16),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_16),
.A2(n_24),
.B1(n_46),
.B2(n_47),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_16),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_71),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_70),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_22),
.B(n_36),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_27),
.B1(n_30),
.B2(n_34),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_23),
.A2(n_27),
.B1(n_30),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_25),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_28),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g101 ( 
.A(n_25),
.B(n_102),
.CON(n_101),
.SN(n_101)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_27),
.A2(n_30),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_27),
.A2(n_30),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_28),
.B(n_32),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_29),
.A2(n_31),
.B1(n_101),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_31),
.B(n_102),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_66),
.C(n_68),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_37),
.A2(n_38),
.B1(n_323),
.B2(n_325),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_49),
.C(n_58),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_39),
.A2(n_294),
.B1(n_295),
.B2(n_297),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_39),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_39),
.A2(n_49),
.B1(n_297),
.B2(n_310),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_45),
.B(n_48),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_40),
.A2(n_45),
.B1(n_86),
.B2(n_88),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_40),
.A2(n_45),
.B1(n_86),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_40),
.A2(n_45),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_40),
.A2(n_45),
.B1(n_156),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_40),
.A2(n_45),
.B1(n_177),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_40),
.A2(n_45),
.B1(n_92),
.B2(n_195),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_40),
.A2(n_45),
.B1(n_88),
.B2(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_40),
.A2(n_45),
.B1(n_231),
.B2(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_40),
.A2(n_45),
.B1(n_48),
.B2(n_264),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_42),
.B(n_53),
.Y(n_187)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_43),
.A2(n_44),
.B(n_102),
.C(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_45),
.B(n_102),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_46),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_47),
.B(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_49),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_56),
.B2(n_57),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_50),
.A2(n_51),
.B1(n_57),
.B2(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_56),
.B(n_57),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_51),
.A2(n_57),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_51),
.A2(n_57),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_52),
.A2(n_55),
.B1(n_96),
.B2(n_98),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_52),
.A2(n_55),
.B1(n_98),
.B2(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_52),
.A2(n_55),
.B1(n_129),
.B2(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_52),
.A2(n_55),
.B1(n_112),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_52),
.A2(n_55),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_58),
.A2(n_59),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_60),
.A2(n_63),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_60),
.A2(n_63),
.B1(n_110),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_60),
.A2(n_63),
.B1(n_238),
.B2(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_324),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_68),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_320),
.B(n_326),
.Y(n_71)
);

OAI321xp33_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_289),
.A3(n_312),
.B1(n_318),
.B2(n_319),
.C(n_328),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_268),
.B(n_288),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_244),
.B(n_267),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_135),
.B(n_220),
.C(n_243),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_120),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_77),
.B(n_120),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_105),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_89),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_79),
.B(n_89),
.C(n_105),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_80),
.B(n_85),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_83),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_81),
.A2(n_82),
.B1(n_118),
.B2(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_81),
.A2(n_145),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_81),
.A2(n_119),
.B1(n_148),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_81),
.A2(n_82),
.B1(n_134),
.B2(n_179),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_81),
.A2(n_84),
.B1(n_119),
.B2(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_81),
.A2(n_82),
.B(n_229),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_82),
.B(n_102),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.C(n_100),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_103),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_114),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_113),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_107),
.B(n_113),
.C(n_114),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_111),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_117),
.Y(n_124)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.C(n_125),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_121),
.B(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.C(n_132),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_127),
.B(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_131),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_219),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_214),
.B(n_218),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_200),
.B(n_213),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_181),
.B(n_199),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_169),
.B(n_180),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_157),
.B(n_168),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_149),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_149),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_153),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_163),
.B(n_167),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_162),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_171),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_178),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_176),
.C(n_178),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_183),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_189),
.B1(n_197),
.B2(n_198),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_184),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_186),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_188),
.Y(n_192)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_193),
.B1(n_194),
.B2(n_196),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_190),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_196),
.C(n_197),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_201),
.B(n_202),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_210),
.C(n_211),
.Y(n_215)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_209),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_210),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_215),
.B(n_216),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_221),
.B(n_222),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_242),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_223),
.Y(n_242)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_232),
.B2(n_233),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_233),
.C(n_242),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_236),
.C(n_241),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_241),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_239),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_245),
.B(n_246),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_266),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_259),
.B2(n_260),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_260),
.C(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_252),
.C(n_256),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_254),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_258),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_265),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_261),
.A2(n_262),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_263),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g303 ( 
.A1(n_262),
.A2(n_280),
.B(n_283),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_263),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_269),
.B(n_270),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_286),
.B2(n_287),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_279),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_273),
.B(n_279),
.C(n_287),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B(n_278),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_275),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_277),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_291),
.C(n_302),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_278),
.A2(n_291),
.B1(n_292),
.B2(n_317),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_278),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_286),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_304),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_290),
.B(n_304),
.Y(n_319)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_298),
.B1(n_300),
.B2(n_301),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_293),
.Y(n_300)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_297),
.C(n_298),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_298),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_298),
.A2(n_301),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_306),
.C(n_311),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_302),
.A2(n_303),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_311),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_313),
.B(n_314),
.Y(n_318)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_322),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_323),
.Y(n_325)
);


endmodule