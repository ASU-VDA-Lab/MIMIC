module fake_jpeg_10549_n_250 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_18),
.Y(n_56)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_26),
.B(n_1),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_51),
.Y(n_71)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_57),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_50),
.B(n_28),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_58),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_59),
.B1(n_32),
.B2(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_20),
.Y(n_73)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_21),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_23),
.B1(n_32),
.B2(n_26),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_63),
.Y(n_74)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_42),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_66),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_67),
.A2(n_80),
.B1(n_83),
.B2(n_28),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_45),
.B1(n_65),
.B2(n_51),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_69),
.A2(n_85),
.B1(n_28),
.B2(n_34),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_43),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_34),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_40),
.B1(n_65),
.B2(n_57),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_72),
.A2(n_92),
.B1(n_93),
.B2(n_28),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_73),
.B(n_89),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_78),
.Y(n_107)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_22),
.B1(n_31),
.B2(n_30),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_54),
.A2(n_31),
.B1(n_30),
.B2(n_42),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_48),
.A2(n_24),
.B1(n_17),
.B2(n_33),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_17),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_1),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_56),
.B(n_17),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_3),
.Y(n_114)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_95),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_52),
.A2(n_24),
.B1(n_33),
.B2(n_34),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_50),
.A2(n_24),
.B1(n_33),
.B2(n_34),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_4),
.Y(n_122)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_64),
.A2(n_24),
.A3(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_96)
);

OAI32xp33_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_34),
.A3(n_29),
.B1(n_27),
.B2(n_6),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_101),
.B(n_109),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_66),
.B1(n_77),
.B2(n_88),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_76),
.B(n_1),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_112),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_106),
.A2(n_120),
.B1(n_118),
.B2(n_110),
.Y(n_146)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_2),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_115),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_116),
.C(n_74),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_71),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

OA21x2_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_3),
.B(n_4),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_87),
.B(n_8),
.Y(n_139)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_124),
.A2(n_128),
.B(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_129),
.Y(n_157)
);

OAI22x1_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_70),
.B1(n_77),
.B2(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_140),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_139),
.B(n_146),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_87),
.C(n_78),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_144),
.C(n_123),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_4),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_86),
.B1(n_84),
.B2(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_84),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_111),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_68),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_68),
.C(n_79),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_147),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_5),
.B(n_8),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_102),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_13),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_168),
.Y(n_191)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_109),
.A3(n_118),
.B1(n_99),
.B2(n_121),
.C1(n_98),
.C2(n_104),
.Y(n_158)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_135),
.A3(n_140),
.B1(n_127),
.B2(n_126),
.C1(n_16),
.C2(n_15),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_160),
.B(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_12),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_100),
.Y(n_164)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_171),
.Y(n_175)
);

INVxp33_ASAP7_75t_SL g170 ( 
.A(n_129),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_100),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_144),
.Y(n_176)
);

NOR2x1_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_10),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_11),
.Y(n_181)
);

XOR2x2_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_146),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_174),
.A2(n_132),
.B(n_136),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_178),
.B(n_181),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_174),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_172),
.A2(n_125),
.B1(n_150),
.B2(n_148),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_167),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_14),
.Y(n_180)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_180),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_135),
.B1(n_14),
.B2(n_16),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_151),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_185),
.B(n_189),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_11),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_186),
.B(n_165),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_157),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_192),
.C(n_162),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_12),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_197),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_164),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_199),
.A2(n_200),
.B(n_201),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_187),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_191),
.A2(n_173),
.B(n_168),
.C(n_152),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_202),
.A2(n_205),
.B1(n_193),
.B2(n_184),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_166),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_192),
.C(n_163),
.Y(n_210)
);

XOR2x2_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_163),
.Y(n_205)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_183),
.C(n_156),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_188),
.A2(n_173),
.B1(n_152),
.B2(n_153),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_208),
.A2(n_159),
.B1(n_155),
.B2(n_160),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_214),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_213),
.C(n_215),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_153),
.B1(n_178),
.B2(n_191),
.Y(n_212)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_205),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_188),
.B1(n_175),
.B2(n_185),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_190),
.C(n_184),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_193),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_220),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_196),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_227),
.C(n_215),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_220),
.A2(n_207),
.B(n_216),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_226),
.B(n_196),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_210),
.Y(n_227)
);

INVxp67_ASAP7_75t_SL g228 ( 
.A(n_219),
.Y(n_228)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_231),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_202),
.B1(n_217),
.B2(n_155),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_233),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_211),
.C(n_197),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_221),
.B(n_195),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_226),
.B(n_166),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_228),
.C(n_198),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_234),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_239),
.B(n_229),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_240),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_151),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_181),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_200),
.B(n_181),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_245),
.B(n_12),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_247),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_248),
.A2(n_246),
.B(n_243),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_238),
.Y(n_250)
);


endmodule