module fake_jpeg_29629_n_142 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_142);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_51),
.A2(n_21),
.B1(n_34),
.B2(n_32),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_40),
.B1(n_55),
.B2(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_0),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_64),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_0),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_69),
.A2(n_74),
.B1(n_79),
.B2(n_4),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_70),
.B(n_73),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_45),
.C(n_53),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_5),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_44),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_46),
.B1(n_50),
.B2(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_3),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_46),
.B1(n_37),
.B2(n_54),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_47),
.B1(n_42),
.B2(n_41),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_94),
.B1(n_17),
.B2(n_18),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_1),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_77),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_24),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_1),
.B(n_2),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_88),
.B(n_85),
.Y(n_105)
);

XNOR2x2_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_22),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_90),
.Y(n_112)
);

INVx5_ASAP7_75t_SL g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_2),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_68),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_15),
.Y(n_109)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_6),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_108),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_82),
.B(n_27),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_113),
.Y(n_121)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_7),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_8),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_110),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_19),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_112),
.B1(n_108),
.B2(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_127),
.Y(n_131)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_123),
.B(n_124),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_122),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_132),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_106),
.B(n_112),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_129),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_102),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_134),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_120),
.C(n_126),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_130),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_125),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_120),
.B(n_135),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_121),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_121),
.B(n_118),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_111),
.Y(n_142)
);


endmodule