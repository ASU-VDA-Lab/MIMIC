module fake_jpeg_14304_n_189 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_189);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_40),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_80),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_72),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_53),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_71),
.B1(n_60),
.B2(n_61),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_59),
.B1(n_66),
.B2(n_62),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_51),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_94),
.B(n_102),
.Y(n_118)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_78),
.C(n_55),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_96),
.A2(n_53),
.B(n_59),
.Y(n_115)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_58),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_76),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_93),
.B(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_104),
.B(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_65),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_106),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_102),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_111),
.B(n_2),
.Y(n_139)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_74),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_117),
.Y(n_126)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_124),
.Y(n_127)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_119),
.A2(n_122),
.B1(n_3),
.B2(n_5),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_56),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_123),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_66),
.B1(n_75),
.B2(n_73),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_63),
.C(n_67),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_137),
.B(n_30),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_139),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_64),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_131),
.B(n_135),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_76),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_0),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_138),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_75),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_1),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_24),
.B1(n_27),
.B2(n_29),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_5),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_143),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_6),
.Y(n_143)
);

AO22x1_ASAP7_75t_SL g148 ( 
.A1(n_132),
.A2(n_50),
.B1(n_34),
.B2(n_37),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_33),
.B1(n_48),
.B2(n_47),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_153),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_152),
.A2(n_156),
.B1(n_130),
.B2(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_9),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_12),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_165),
.C(n_42),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_146),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_133),
.B(n_23),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_141),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_144),
.B1(n_149),
.B2(n_148),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_161),
.B(n_125),
.Y(n_170)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_145),
.B(n_38),
.CI(n_39),
.CON(n_161),
.SN(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_41),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_169),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_174),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_172),
.B(n_173),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_153),
.C(n_163),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_180),
.A2(n_154),
.B1(n_151),
.B2(n_167),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_178),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_171),
.C(n_176),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_171),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_181),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_164),
.B(n_175),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_179),
.B(n_150),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_44),
.Y(n_189)
);


endmodule