module real_jpeg_26877_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_309, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_309;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;

INVx11_ASAP7_75t_L g93 ( 
.A(n_0),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_1),
.A2(n_39),
.B1(n_57),
.B2(n_58),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_1),
.A2(n_39),
.B1(n_45),
.B2(n_47),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_2),
.A2(n_57),
.B1(n_58),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_2),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_133),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_2),
.A2(n_45),
.B1(n_47),
.B2(n_133),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_133),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_3),
.A2(n_57),
.B1(n_58),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_3),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_SL g159 ( 
.A1(n_3),
.A2(n_29),
.B(n_63),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_3),
.B(n_65),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_3),
.A2(n_32),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_3),
.B(n_32),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_3),
.B(n_74),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_3),
.A2(n_90),
.B1(n_94),
.B2(n_236),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_3),
.A2(n_28),
.B(n_252),
.Y(n_251)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_5),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_100),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_100),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_5),
.A2(n_45),
.B1(n_47),
.B2(n_100),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_7),
.A2(n_45),
.B1(n_47),
.B2(n_52),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_52),
.Y(n_109)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_9),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_9),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_60),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g150 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_60),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_9),
.A2(n_45),
.B1(n_47),
.B2(n_60),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_50),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_10),
.A2(n_45),
.B1(n_47),
.B2(n_50),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g143 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_144),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_11),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_11),
.A2(n_57),
.B1(n_58),
.B2(n_144),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_144),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_11),
.A2(n_45),
.B1(n_47),
.B2(n_144),
.Y(n_229)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_13),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_156),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_156),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_13),
.A2(n_45),
.B1(n_47),
.B2(n_156),
.Y(n_236)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_16),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_17),
.A2(n_28),
.B1(n_29),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_17),
.A2(n_37),
.B1(n_57),
.B2(n_58),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_17),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_17),
.A2(n_37),
.B1(n_45),
.B2(n_47),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_114),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_113),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_101),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_22),
.B(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_22),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_22),
.B(n_116),
.Y(n_306)
);

FAx1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.CI(n_79),
.CON(n_22),
.SN(n_22)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_23),
.A2(n_24),
.B(n_40),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_35),
.B2(n_38),
.Y(n_24)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_25),
.A2(n_31),
.B1(n_142),
.B2(n_145),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_25),
.A2(n_31),
.B1(n_145),
.B2(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_25),
.A2(n_31),
.B1(n_167),
.B2(n_251),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_28),
.Y(n_30)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

OAI32xp33_ASAP7_75t_L g260 ( 
.A1(n_26),
.A2(n_28),
.A3(n_33),
.B1(n_253),
.B2(n_261),
.Y(n_260)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AO22x1_ASAP7_75t_L g65 ( 
.A1(n_28),
.A2(n_29),
.B1(n_63),
.B2(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_29),
.B(n_153),
.Y(n_253)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_33),
.B1(n_43),
.B2(n_44),
.Y(n_48)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_32),
.A2(n_43),
.A3(n_47),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_32),
.B(n_34),
.Y(n_261)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_36),
.A2(n_72),
.B1(n_74),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_38),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_49),
.B2(n_51),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_41),
.A2(n_42),
.B(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_41),
.A2(n_42),
.B1(n_85),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_41),
.A2(n_42),
.B1(n_128),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_41),
.A2(n_42),
.B1(n_208),
.B2(n_210),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_41),
.A2(n_42),
.B1(n_210),
.B2(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_41),
.A2(n_42),
.B1(n_149),
.B2(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_48),
.Y(n_41)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_42),
.B(n_153),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_44),
.B(n_45),
.Y(n_214)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_45),
.B(n_242),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_49),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_69),
.B2(n_78),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_54),
.A2(n_55),
.B1(n_103),
.B2(n_111),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_55),
.B(n_70),
.C(n_77),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_61),
.B1(n_67),
.B2(n_68),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_61),
.B1(n_68),
.B2(n_98),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_63),
.B(n_64),
.C(n_65),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g64 ( 
.A(n_57),
.B(n_63),
.Y(n_64)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_58),
.A2(n_66),
.B(n_153),
.C(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_61),
.A2(n_68),
.B1(n_155),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_65),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_62),
.A2(n_65),
.B1(n_99),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_62),
.A2(n_65),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_62),
.A2(n_65),
.B1(n_132),
.B2(n_183),
.Y(n_197)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_72),
.A2(n_74),
.B1(n_143),
.B2(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_72),
.A2(n_74),
.B1(n_130),
.B2(n_186),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_75),
.A2(n_77),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_96),
.B(n_97),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_80),
.A2(n_81),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_89),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_82),
.A2(n_83),
.B1(n_89),
.B2(n_96),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_86),
.A2(n_88),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_86),
.A2(n_88),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_96),
.B1(n_97),
.B2(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_94),
.B(n_95),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_90),
.A2(n_94),
.B1(n_95),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_90),
.A2(n_94),
.B1(n_126),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_90),
.A2(n_94),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_90),
.A2(n_229),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_90),
.A2(n_94),
.B1(n_224),
.B2(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_91),
.A2(n_92),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_91),
.A2(n_92),
.B1(n_161),
.B2(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_91),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

INVx5_ASAP7_75t_SL g237 ( 
.A(n_92),
.Y(n_237)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_94),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_94),
.B(n_153),
.Y(n_242)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_112),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_108),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_134),
.B(n_306),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_122),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_117),
.B(n_121),
.Y(n_294)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_122),
.A2(n_123),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.C(n_131),
.Y(n_123)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_124),
.B(n_129),
.CI(n_131),
.CON(n_289),
.SN(n_289)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_125),
.B(n_127),
.Y(n_193)
);

AOI321xp33_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_287),
.A3(n_295),
.B1(n_300),
.B2(n_305),
.C(n_309),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_188),
.C(n_200),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_171),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_137),
.B(n_171),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_157),
.C(n_163),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_138),
.B(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_151),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_146),
.B2(n_147),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_147),
.C(n_151),
.Y(n_178)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_157),
.A2(n_163),
.B1(n_164),
.B2(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_157),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_160),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_162),
.Y(n_177)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_170),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_165),
.B(n_272),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_168),
.B(n_170),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_169),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_179),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_178),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_178),
.C(n_179),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_176),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_187),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_184),
.C(n_187),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_L g301 ( 
.A1(n_189),
.A2(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_190),
.B(n_191),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_199),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_193),
.B(n_194),
.C(n_199),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_195),
.B(n_197),
.C(n_198),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_281),
.B(n_286),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_267),
.B(n_280),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_246),
.B(n_266),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_225),
.B(n_245),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_215),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_205),
.B(n_215),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_206),
.A2(n_207),
.B1(n_211),
.B2(n_212),
.Y(n_232)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_209),
.Y(n_213)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_222),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_220),
.C(n_222),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_221),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_223),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_233),
.B(n_244),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_232),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_227),
.B(n_232),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_239),
.B(n_243),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_235),
.B(n_238),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_247),
.B(n_248),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_259),
.B1(n_264),
.B2(n_265),
.Y(n_248)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_254),
.B1(n_257),
.B2(n_258),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_250),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_254),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_258),
.C(n_265),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_256),
.Y(n_277)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_259),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_262),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_268),
.B(n_269),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_273),
.B2(n_274),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_276),
.C(n_278),
.Y(n_282)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_279),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_276),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_292),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_292),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.C(n_291),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_290),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_289),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_296),
.A2(n_301),
.B(n_304),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_297),
.B(n_298),
.Y(n_304)
);


endmodule