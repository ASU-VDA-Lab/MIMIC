module fake_netlist_6_694_n_1090 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1090);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1090;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_952;
wire n_725;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_1018;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_720;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_886;
wire n_448;
wire n_953;
wire n_1017;
wire n_1004;
wire n_844;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_236;
wire n_653;
wire n_887;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_964;
wire n_982;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_409;
wire n_345;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_249;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_928;
wire n_835;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx2_ASAP7_75t_SL g213 ( 
.A(n_188),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_116),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_4),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_7),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_10),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_175),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_140),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_110),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_164),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_53),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_92),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_18),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_10),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_138),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_66),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_165),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_101),
.Y(n_230)
);

BUFx8_ASAP7_75t_SL g231 ( 
.A(n_155),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_93),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_69),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_41),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_43),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_35),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_157),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_150),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_131),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_74),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_204),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_22),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_195),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_156),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_15),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_160),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_162),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_168),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_153),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_54),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_147),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_115),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_118),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_55),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_135),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_25),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_73),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_81),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_186),
.Y(n_259)
);

BUFx8_ASAP7_75t_SL g260 ( 
.A(n_119),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_171),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_44),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_8),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_177),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_114),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_90),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_14),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_63),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_58),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_56),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_2),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_24),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_77),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_19),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_128),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_109),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_30),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_148),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_61),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_130),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_19),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_39),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_181),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_225),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_227),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_228),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_227),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_256),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_228),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_233),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g292 ( 
.A(n_231),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_236),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_236),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_223),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_257),
.Y(n_297)
);

INVxp33_ASAP7_75t_SL g298 ( 
.A(n_215),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g299 ( 
.A(n_231),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_227),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_230),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_232),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_234),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_235),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_238),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_239),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_240),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_247),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_244),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_253),
.Y(n_311)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_216),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_280),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_262),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_233),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_268),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_269),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_283),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_241),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_244),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_271),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_241),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_217),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_226),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_242),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_263),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_267),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_274),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_277),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_213),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_288),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_282),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_297),
.A2(n_279),
.B1(n_313),
.B2(n_289),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_288),
.Y(n_337)
);

OAI21x1_ASAP7_75t_L g338 ( 
.A1(n_310),
.A2(n_264),
.B(n_221),
.Y(n_338)
);

OAI21x1_ASAP7_75t_L g339 ( 
.A1(n_310),
.A2(n_264),
.B(n_221),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_286),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_289),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_286),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_295),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_286),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_295),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_314),
.B(n_270),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_291),
.A2(n_279),
.B1(n_281),
.B2(n_219),
.Y(n_347)
);

BUFx8_ASAP7_75t_L g348 ( 
.A(n_327),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_291),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_300),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_300),
.Y(n_351)
);

AND2x4_ASAP7_75t_L g352 ( 
.A(n_296),
.B(n_278),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_286),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_320),
.Y(n_354)
);

CKINVDCx6p67_ASAP7_75t_R g355 ( 
.A(n_315),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_333),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_298),
.B(n_218),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_321),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_301),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_333),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_218),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_287),
.B(n_218),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_302),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_284),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_315),
.A2(n_276),
.B1(n_275),
.B2(n_273),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_285),
.Y(n_367)
);

OAI21x1_ASAP7_75t_L g368 ( 
.A1(n_303),
.A2(n_221),
.B(n_220),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_304),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_305),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_326),
.B(n_214),
.Y(n_372)
);

CKINVDCx8_ASAP7_75t_R g373 ( 
.A(n_327),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_328),
.B(n_266),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_333),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_306),
.Y(n_377)
);

BUFx8_ASAP7_75t_SL g378 ( 
.A(n_319),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_298),
.A2(n_265),
.B1(n_261),
.B2(n_222),
.Y(n_379)
);

AND2x6_ASAP7_75t_L g380 ( 
.A(n_307),
.B(n_260),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_308),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_309),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_330),
.B(n_332),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_311),
.Y(n_384)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_290),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_331),
.B(n_224),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_316),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_293),
.B(n_229),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_378),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_343),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_R g391 ( 
.A(n_373),
.B(n_319),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_343),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_371),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_357),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_371),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_349),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_346),
.B(n_292),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_355),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_355),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_376),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_348),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_336),
.A2(n_324),
.B1(n_312),
.B2(n_292),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_376),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_348),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

NAND2xp33_ASAP7_75t_R g406 ( 
.A(n_354),
.B(n_312),
.Y(n_406)
);

BUFx10_ASAP7_75t_L g407 ( 
.A(n_362),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_348),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_382),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_382),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_350),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_350),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_340),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_373),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_384),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_366),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_366),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_340),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_341),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_346),
.B(n_299),
.Y(n_420)
);

AOI21x1_ASAP7_75t_L g421 ( 
.A1(n_335),
.A2(n_318),
.B(n_317),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_379),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_379),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_383),
.B(n_294),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_386),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_384),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_354),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_372),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_374),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_334),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_365),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_365),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_367),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_336),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_347),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_388),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_388),
.Y(n_437)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_340),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_358),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_380),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_SL g441 ( 
.A(n_363),
.B(n_299),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_R g442 ( 
.A(n_346),
.B(n_322),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_334),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_380),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_346),
.B(n_237),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_380),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_367),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_380),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_340),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_380),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_377),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_352),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_352),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_352),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_363),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_R g456 ( 
.A(n_387),
.B(n_324),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_340),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_352),
.B(n_243),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_428),
.B(n_385),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_396),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_409),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_410),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_429),
.B(n_385),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_415),
.Y(n_464)
);

AND2x6_ASAP7_75t_L g465 ( 
.A(n_397),
.B(n_323),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_426),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_431),
.B(n_385),
.Y(n_467)
);

BUFx10_ASAP7_75t_L g468 ( 
.A(n_389),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_390),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_390),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_425),
.B(n_246),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_436),
.B(n_377),
.Y(n_472)
);

NAND2x1p5_ASAP7_75t_L g473 ( 
.A(n_432),
.B(n_338),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_424),
.B(n_387),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_433),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_391),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_447),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_430),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_427),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_R g480 ( 
.A(n_414),
.B(n_442),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_399),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_424),
.B(n_387),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_430),
.B(n_368),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_392),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_443),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_407),
.B(n_260),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_413),
.Y(n_487)
);

AO22x2_ASAP7_75t_L g488 ( 
.A1(n_420),
.A2(n_368),
.B1(n_360),
.B2(n_364),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_437),
.B(n_360),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_452),
.B(n_249),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_443),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_456),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_442),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_421),
.B(n_364),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_456),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_411),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_453),
.B(n_250),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_454),
.B(n_369),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_411),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_407),
.B(n_381),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_455),
.A2(n_439),
.B1(n_445),
.B2(n_458),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_412),
.B(n_337),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_422),
.B(n_381),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_451),
.B(n_337),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_419),
.B(n_369),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_393),
.B(n_370),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_395),
.B(n_370),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_423),
.B(n_251),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_400),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_403),
.Y(n_510)
);

NAND3xp33_ASAP7_75t_L g511 ( 
.A(n_405),
.B(n_351),
.C(n_345),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_418),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_441),
.B(n_252),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_418),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_394),
.B(n_359),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_449),
.B(n_359),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_398),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_402),
.B(n_338),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_401),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_449),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_391),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_406),
.A2(n_254),
.B1(n_255),
.B2(n_258),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_434),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_416),
.B(n_417),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_457),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_413),
.B(n_345),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_435),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_438),
.B(n_351),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_440),
.B(n_377),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_444),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_446),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_448),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_450),
.B(n_377),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_493),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_493),
.B(n_404),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_478),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_485),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_491),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_508),
.B(n_408),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_461),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_503),
.B(n_406),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_469),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_462),
.Y(n_544)
);

A2O1A1Ixp33_ASAP7_75t_L g545 ( 
.A1(n_474),
.A2(n_339),
.B(n_259),
.C(n_377),
.Y(n_545)
);

NAND3xp33_ASAP7_75t_L g546 ( 
.A(n_474),
.B(n_361),
.C(n_357),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_466),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_482),
.B(n_353),
.Y(n_548)
);

NOR3xp33_ASAP7_75t_L g549 ( 
.A(n_525),
.B(n_356),
.C(n_342),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_480),
.B(n_357),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_464),
.B(n_36),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_482),
.B(n_472),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_475),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_477),
.Y(n_554)
);

BUFx8_ASAP7_75t_L g555 ( 
.A(n_524),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_506),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_505),
.B(n_357),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_489),
.B(n_357),
.Y(n_558)
);

INVx8_ASAP7_75t_L g559 ( 
.A(n_465),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_506),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_507),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_472),
.B(n_353),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_507),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_504),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_517),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_504),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_533),
.B(n_361),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_460),
.Y(n_568)
);

OAI221xp5_ASAP7_75t_L g569 ( 
.A1(n_519),
.A2(n_356),
.B1(n_342),
.B2(n_375),
.C(n_361),
.Y(n_569)
);

AO22x2_ASAP7_75t_L g570 ( 
.A1(n_492),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_498),
.B(n_37),
.Y(n_571)
);

AND2x4_ASAP7_75t_SL g572 ( 
.A(n_468),
.B(n_498),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_500),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_467),
.B(n_38),
.Y(n_574)
);

BUFx8_ASAP7_75t_L g575 ( 
.A(n_479),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_528),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_576)
);

BUFx8_ASAP7_75t_L g577 ( 
.A(n_520),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_467),
.B(n_361),
.Y(n_578)
);

NAND2x1p5_ASAP7_75t_L g579 ( 
.A(n_532),
.B(n_375),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_484),
.Y(n_580)
);

OAI221xp5_ASAP7_75t_L g581 ( 
.A1(n_501),
.A2(n_356),
.B1(n_375),
.B2(n_344),
.C(n_6),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_494),
.A2(n_375),
.B1(n_344),
.B2(n_5),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_470),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_516),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_502),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_496),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_R g587 ( 
.A(n_476),
.B(n_40),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_499),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_522),
.B(n_42),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_494),
.A2(n_344),
.B1(n_4),
.B2(n_5),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_488),
.A2(n_344),
.B1(n_6),
.B2(n_7),
.Y(n_591)
);

OR2x2_ASAP7_75t_SL g592 ( 
.A(n_528),
.B(n_3),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_487),
.B(n_344),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_502),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_592),
.A2(n_495),
.B1(n_486),
.B2(n_481),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_552),
.A2(n_534),
.B(n_530),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_552),
.A2(n_534),
.B(n_530),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_542),
.B(n_573),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_568),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_565),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_535),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_573),
.B(n_495),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_564),
.B(n_465),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_535),
.B(n_471),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_548),
.A2(n_545),
.B(n_585),
.Y(n_605)
);

AOI22x1_ASAP7_75t_L g606 ( 
.A1(n_594),
.A2(n_488),
.B1(n_473),
.B2(n_531),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_566),
.B(n_465),
.Y(n_607)
);

AND2x4_ASAP7_75t_SL g608 ( 
.A(n_571),
.B(n_468),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_562),
.A2(n_515),
.B(n_532),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_558),
.B(n_465),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_571),
.B(n_551),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_565),
.Y(n_612)
);

O2A1O1Ixp33_ASAP7_75t_L g613 ( 
.A1(n_581),
.A2(n_459),
.B(n_463),
.C(n_513),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_557),
.B(n_515),
.Y(n_614)
);

AND2x2_ASAP7_75t_SL g615 ( 
.A(n_540),
.B(n_532),
.Y(n_615)
);

BUFx4f_ASAP7_75t_L g616 ( 
.A(n_572),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_543),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_565),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_574),
.A2(n_497),
.B1(n_490),
.B2(n_523),
.Y(n_619)
);

OAI321xp33_ASAP7_75t_L g620 ( 
.A1(n_576),
.A2(n_483),
.A3(n_473),
.B1(n_510),
.B2(n_509),
.C(n_511),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_536),
.B(n_518),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_575),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_593),
.A2(n_548),
.B(n_578),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_541),
.B(n_488),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_544),
.B(n_512),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_575),
.Y(n_626)
);

NOR3xp33_ASAP7_75t_L g627 ( 
.A(n_556),
.B(n_511),
.C(n_512),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_569),
.A2(n_527),
.B(n_521),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_569),
.A2(n_527),
.B(n_526),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_547),
.B(n_514),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_551),
.B(n_529),
.Y(n_631)
);

O2A1O1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_553),
.A2(n_8),
.B(n_9),
.C(n_11),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_546),
.A2(n_550),
.B(n_559),
.Y(n_633)
);

O2A1O1Ixp33_ASAP7_75t_L g634 ( 
.A1(n_554),
.A2(n_9),
.B(n_11),
.C(n_12),
.Y(n_634)
);

AOI21x1_ASAP7_75t_L g635 ( 
.A1(n_537),
.A2(n_46),
.B(n_45),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_538),
.B(n_12),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_539),
.B(n_583),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_559),
.A2(n_48),
.B(n_47),
.Y(n_638)
);

AO22x1_ASAP7_75t_L g639 ( 
.A1(n_589),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_579),
.A2(n_50),
.B(n_49),
.Y(n_640)
);

INVx1_ASAP7_75t_SL g641 ( 
.A(n_587),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_582),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_559),
.A2(n_52),
.B(n_51),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_586),
.B(n_57),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_560),
.B(n_16),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_588),
.B(n_59),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_598),
.B(n_602),
.Y(n_647)
);

A2O1A1Ixp33_ASAP7_75t_SL g648 ( 
.A1(n_605),
.A2(n_549),
.B(n_591),
.C(n_590),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_615),
.B(n_611),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_619),
.B(n_589),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_601),
.Y(n_651)
);

OAI21xp33_ASAP7_75t_SL g652 ( 
.A1(n_603),
.A2(n_584),
.B(n_563),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_604),
.B(n_561),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_637),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_642),
.A2(n_549),
.B1(n_570),
.B2(n_580),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_637),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_616),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_621),
.B(n_614),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_617),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_645),
.B(n_570),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_597),
.A2(n_609),
.B(n_605),
.Y(n_661)
);

OA21x2_ASAP7_75t_L g662 ( 
.A1(n_606),
.A2(n_623),
.B(n_628),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_608),
.B(n_567),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_625),
.Y(n_664)
);

A2O1A1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_613),
.A2(n_567),
.B(n_577),
.C(n_555),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_618),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_631),
.A2(n_62),
.B(n_60),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_599),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_630),
.Y(n_669)
);

AO31x2_ASAP7_75t_L g670 ( 
.A1(n_624),
.A2(n_17),
.A3(n_18),
.B(n_20),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_633),
.A2(n_127),
.B(n_212),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_641),
.B(n_555),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_636),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_618),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_600),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_644),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_616),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_600),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_644),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_607),
.B(n_627),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_610),
.A2(n_577),
.B1(n_21),
.B2(n_22),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_629),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_612),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_646),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_646),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_612),
.Y(n_686)
);

BUFx12f_ASAP7_75t_L g687 ( 
.A(n_622),
.Y(n_687)
);

OAI321xp33_ASAP7_75t_L g688 ( 
.A1(n_632),
.A2(n_23),
.A3(n_24),
.B1(n_25),
.B2(n_26),
.C(n_27),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_638),
.A2(n_132),
.B(n_210),
.Y(n_689)
);

BUFx2_ASAP7_75t_L g690 ( 
.A(n_595),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_639),
.Y(n_691)
);

A2O1A1Ixp33_ASAP7_75t_SL g692 ( 
.A1(n_620),
.A2(n_129),
.B(n_209),
.C(n_208),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_634),
.B(n_643),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_640),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_SL g695 ( 
.A(n_626),
.B(n_64),
.Y(n_695)
);

OAI21xp33_ASAP7_75t_SL g696 ( 
.A1(n_635),
.A2(n_26),
.B(n_27),
.Y(n_696)
);

INVxp67_ASAP7_75t_L g697 ( 
.A(n_601),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_596),
.A2(n_133),
.B(n_207),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_599),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_616),
.Y(n_700)
);

O2A1O1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_613),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_647),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_657),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_668),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_659),
.Y(n_705)
);

BUFx2_ASAP7_75t_SL g706 ( 
.A(n_699),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_651),
.Y(n_707)
);

INVxp67_ASAP7_75t_SL g708 ( 
.A(n_654),
.Y(n_708)
);

BUFx5_ASAP7_75t_L g709 ( 
.A(n_694),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_657),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_658),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_656),
.B(n_28),
.Y(n_712)
);

BUFx12f_ASAP7_75t_L g713 ( 
.A(n_657),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_687),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_677),
.Y(n_715)
);

BUFx12f_ASAP7_75t_L g716 ( 
.A(n_677),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_677),
.Y(n_717)
);

BUFx2_ASAP7_75t_SL g718 ( 
.A(n_700),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_700),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_700),
.B(n_65),
.Y(n_720)
);

INVx6_ASAP7_75t_SL g721 ( 
.A(n_663),
.Y(n_721)
);

BUFx4f_ASAP7_75t_SL g722 ( 
.A(n_678),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_672),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_678),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_678),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_674),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_653),
.B(n_29),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_650),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_675),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_664),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_690),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_666),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_686),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_683),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_650),
.B(n_31),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_663),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_649),
.Y(n_737)
);

NAND2x1p5_ASAP7_75t_L g738 ( 
.A(n_691),
.B(n_67),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_650),
.B(n_32),
.Y(n_739)
);

BUFx6f_ASAP7_75t_SL g740 ( 
.A(n_669),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_673),
.Y(n_741)
);

BUFx8_ASAP7_75t_SL g742 ( 
.A(n_660),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_650),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_676),
.B(n_33),
.Y(n_744)
);

INVx6_ASAP7_75t_SL g745 ( 
.A(n_697),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_679),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_680),
.Y(n_747)
);

BUFx2_ASAP7_75t_SL g748 ( 
.A(n_681),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_670),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_684),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_670),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_665),
.B(n_68),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_693),
.Y(n_753)
);

INVx6_ASAP7_75t_L g754 ( 
.A(n_695),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_655),
.B(n_34),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_682),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_685),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_652),
.A2(n_34),
.B1(n_70),
.B2(n_71),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_696),
.Y(n_759)
);

AO21x2_ASAP7_75t_L g760 ( 
.A1(n_661),
.A2(n_72),
.B(n_75),
.Y(n_760)
);

INVx5_ASAP7_75t_L g761 ( 
.A(n_692),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_662),
.Y(n_762)
);

BUFx24_ASAP7_75t_L g763 ( 
.A(n_688),
.Y(n_763)
);

INVx5_ASAP7_75t_SL g764 ( 
.A(n_689),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_667),
.B(n_76),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_701),
.Y(n_766)
);

BUFx2_ASAP7_75t_SL g767 ( 
.A(n_671),
.Y(n_767)
);

INVx4_ASAP7_75t_L g768 ( 
.A(n_698),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_747),
.B(n_648),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_746),
.A2(n_78),
.B(n_79),
.Y(n_770)
);

OAI222xp33_ASAP7_75t_L g771 ( 
.A1(n_728),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.C1(n_84),
.C2(n_85),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_736),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_728),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_773)
);

OAI21x1_ASAP7_75t_L g774 ( 
.A1(n_746),
.A2(n_89),
.B(n_91),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_711),
.B(n_94),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_750),
.A2(n_95),
.B(n_96),
.Y(n_776)
);

OAI21x1_ASAP7_75t_L g777 ( 
.A1(n_735),
.A2(n_97),
.B(n_98),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_748),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_778)
);

NAND2xp33_ASAP7_75t_L g779 ( 
.A(n_747),
.B(n_103),
.Y(n_779)
);

O2A1O1Ixp33_ASAP7_75t_SL g780 ( 
.A1(n_735),
.A2(n_104),
.B(n_105),
.C(n_106),
.Y(n_780)
);

O2A1O1Ixp33_ASAP7_75t_SL g781 ( 
.A1(n_766),
.A2(n_107),
.B(n_108),
.C(n_111),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_708),
.B(n_112),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_737),
.B(n_113),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_713),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_708),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_755),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_711),
.B(n_122),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_732),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_758),
.A2(n_753),
.B(n_756),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_SL g790 ( 
.A1(n_731),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_705),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_743),
.B(n_126),
.Y(n_792)
);

OAI21x1_ASAP7_75t_L g793 ( 
.A1(n_739),
.A2(n_134),
.B(n_136),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_736),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_730),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_739),
.A2(n_137),
.B(n_139),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_737),
.B(n_141),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_706),
.Y(n_798)
);

AO21x2_ASAP7_75t_L g799 ( 
.A1(n_760),
.A2(n_142),
.B(n_143),
.Y(n_799)
);

OA21x2_ASAP7_75t_L g800 ( 
.A1(n_759),
.A2(n_144),
.B(n_145),
.Y(n_800)
);

XOR2xp5_ASAP7_75t_L g801 ( 
.A(n_704),
.B(n_146),
.Y(n_801)
);

O2A1O1Ixp33_ASAP7_75t_SL g802 ( 
.A1(n_744),
.A2(n_149),
.B(n_151),
.C(n_152),
.Y(n_802)
);

O2A1O1Ixp33_ASAP7_75t_SL g803 ( 
.A1(n_744),
.A2(n_154),
.B(n_158),
.C(n_159),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_716),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_702),
.B(n_161),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_757),
.Y(n_806)
);

AO31x2_ASAP7_75t_L g807 ( 
.A1(n_768),
.A2(n_163),
.A3(n_166),
.B(n_167),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_741),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_702),
.B(n_169),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_749),
.Y(n_810)
);

INVx4_ASAP7_75t_L g811 ( 
.A(n_722),
.Y(n_811)
);

OAI21x1_ASAP7_75t_L g812 ( 
.A1(n_738),
.A2(n_170),
.B(n_172),
.Y(n_812)
);

OAI21x1_ASAP7_75t_L g813 ( 
.A1(n_712),
.A2(n_173),
.B(n_174),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_729),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_752),
.A2(n_176),
.B(n_178),
.C(n_179),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_761),
.A2(n_180),
.B(n_182),
.Y(n_816)
);

OAI21x1_ASAP7_75t_SL g817 ( 
.A1(n_712),
.A2(n_183),
.B(n_184),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_752),
.B(n_185),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_751),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_754),
.A2(n_727),
.B1(n_763),
.B2(n_740),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_754),
.B(n_187),
.Y(n_821)
);

AO21x2_ASAP7_75t_L g822 ( 
.A1(n_760),
.A2(n_189),
.B(n_190),
.Y(n_822)
);

O2A1O1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_726),
.A2(n_191),
.B(n_192),
.C(n_193),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_733),
.Y(n_824)
);

OAI21x1_ASAP7_75t_L g825 ( 
.A1(n_767),
.A2(n_194),
.B(n_196),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_795),
.Y(n_826)
);

INVxp67_ASAP7_75t_SL g827 ( 
.A(n_785),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_SL g828 ( 
.A1(n_820),
.A2(n_754),
.B1(n_763),
.B2(n_740),
.Y(n_828)
);

AOI21x1_ASAP7_75t_L g829 ( 
.A1(n_769),
.A2(n_765),
.B(n_720),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_810),
.Y(n_830)
);

OAI22xp33_ASAP7_75t_L g831 ( 
.A1(n_820),
.A2(n_723),
.B1(n_761),
.B2(n_768),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_808),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_819),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_791),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_788),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_769),
.Y(n_836)
);

INVx1_ASAP7_75t_SL g837 ( 
.A(n_782),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_807),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_807),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_806),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_807),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_799),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_782),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_799),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_822),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_822),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_813),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_800),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_816),
.A2(n_761),
.B(n_707),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_806),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_772),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_800),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_789),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_789),
.B(n_816),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_777),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_793),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_770),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_796),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_814),
.B(n_709),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_774),
.Y(n_860)
);

OAI21x1_ASAP7_75t_L g861 ( 
.A1(n_776),
.A2(n_762),
.B(n_764),
.Y(n_861)
);

OAI21x1_ASAP7_75t_L g862 ( 
.A1(n_825),
.A2(n_764),
.B(n_761),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_787),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_787),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_809),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_824),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_809),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_817),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_854),
.A2(n_818),
.B1(n_790),
.B2(n_773),
.Y(n_869)
);

BUFx10_ASAP7_75t_L g870 ( 
.A(n_836),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_832),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_840),
.Y(n_872)
);

CKINVDCx6p67_ASAP7_75t_R g873 ( 
.A(n_851),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_852),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_850),
.B(n_798),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_830),
.B(n_804),
.Y(n_876)
);

OR2x2_ASAP7_75t_L g877 ( 
.A(n_837),
.B(n_805),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_859),
.B(n_784),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_854),
.A2(n_773),
.B1(n_818),
.B2(n_786),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_R g880 ( 
.A(n_829),
.B(n_779),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_826),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_R g882 ( 
.A(n_829),
.B(n_722),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_R g883 ( 
.A(n_836),
.B(n_714),
.Y(n_883)
);

OR2x6_ASAP7_75t_L g884 ( 
.A(n_854),
.B(n_812),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_851),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_837),
.B(n_783),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_832),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_843),
.B(n_797),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_826),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_859),
.B(n_775),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_851),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_832),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_834),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_865),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_854),
.A2(n_821),
.B1(n_786),
.B2(n_792),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_830),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_R g897 ( 
.A(n_853),
.B(n_772),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_866),
.Y(n_898)
);

AO32x2_ASAP7_75t_L g899 ( 
.A1(n_827),
.A2(n_811),
.A3(n_715),
.B1(n_742),
.B2(n_771),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_830),
.B(n_794),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_866),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_833),
.Y(n_902)
);

AO31x2_ASAP7_75t_L g903 ( 
.A1(n_839),
.A2(n_841),
.A3(n_845),
.B(n_842),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_834),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_843),
.B(n_783),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_854),
.A2(n_815),
.B1(n_778),
.B2(n_821),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_874),
.B(n_900),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_903),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_886),
.B(n_877),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_874),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_894),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_881),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_870),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_889),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_903),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_871),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_903),
.Y(n_917)
);

INVx4_ASAP7_75t_L g918 ( 
.A(n_885),
.Y(n_918)
);

INVxp67_ASAP7_75t_SL g919 ( 
.A(n_886),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_887),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_902),
.B(n_848),
.Y(n_921)
);

INVxp67_ASAP7_75t_SL g922 ( 
.A(n_872),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_892),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_898),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_878),
.B(n_848),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_876),
.B(n_865),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_905),
.B(n_863),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_901),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_893),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_904),
.B(n_853),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_897),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_930),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_931),
.A2(n_854),
.B1(n_906),
.B2(n_879),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_931),
.A2(n_906),
.B1(n_879),
.B2(n_849),
.Y(n_934)
);

AOI221xp5_ASAP7_75t_L g935 ( 
.A1(n_919),
.A2(n_849),
.B1(n_867),
.B2(n_864),
.C(n_863),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_913),
.B(n_900),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_930),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_918),
.A2(n_869),
.B1(n_895),
.B2(n_828),
.Y(n_938)
);

OAI21xp33_ASAP7_75t_L g939 ( 
.A1(n_909),
.A2(n_880),
.B(n_828),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_922),
.A2(n_771),
.B(n_823),
.Y(n_940)
);

NAND4xp25_ASAP7_75t_SL g941 ( 
.A(n_927),
.B(n_875),
.C(n_823),
.D(n_852),
.Y(n_941)
);

OAI22xp33_ASAP7_75t_L g942 ( 
.A1(n_918),
.A2(n_884),
.B1(n_868),
.B2(n_831),
.Y(n_942)
);

NAND3xp33_ASAP7_75t_L g943 ( 
.A(n_926),
.B(n_867),
.C(n_864),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_912),
.Y(n_944)
);

NAND4xp25_ASAP7_75t_L g945 ( 
.A(n_918),
.B(n_888),
.C(n_868),
.D(n_910),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_907),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_913),
.A2(n_868),
.B(n_848),
.C(n_876),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_912),
.Y(n_948)
);

OAI221xp5_ASAP7_75t_L g949 ( 
.A1(n_934),
.A2(n_939),
.B1(n_933),
.B2(n_938),
.C(n_940),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_932),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_944),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_941),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_948),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_936),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_937),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_946),
.B(n_907),
.Y(n_956)
);

INVx4_ASAP7_75t_L g957 ( 
.A(n_936),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_947),
.B(n_907),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_943),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_940),
.A2(n_884),
.B1(n_880),
.B2(n_882),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_950),
.B(n_945),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_955),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_951),
.Y(n_963)
);

AND2x4_ASAP7_75t_SL g964 ( 
.A(n_957),
.B(n_918),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_SL g965 ( 
.A1(n_952),
.A2(n_942),
.B(n_801),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_955),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_959),
.B(n_911),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_953),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_962),
.B(n_959),
.Y(n_969)
);

OAI31xp33_ASAP7_75t_L g970 ( 
.A1(n_965),
.A2(n_949),
.A3(n_960),
.B(n_954),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_966),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_967),
.B(n_954),
.Y(n_972)
);

NAND3xp33_ASAP7_75t_L g973 ( 
.A(n_965),
.B(n_935),
.C(n_957),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_964),
.A2(n_957),
.B1(n_958),
.B2(n_956),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_961),
.B(n_953),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_971),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_975),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_974),
.B(n_956),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_969),
.B(n_972),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_973),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_970),
.B(n_963),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_971),
.B(n_968),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_971),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_972),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_974),
.B(n_958),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_971),
.B(n_910),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_980),
.A2(n_891),
.B1(n_913),
.B2(n_873),
.Y(n_987)
);

NOR2x1_ASAP7_75t_L g988 ( 
.A(n_981),
.B(n_811),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_984),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_979),
.B(n_914),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_977),
.Y(n_991)
);

INVxp67_ASAP7_75t_SL g992 ( 
.A(n_981),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_978),
.B(n_907),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_976),
.B(n_914),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_992),
.A2(n_985),
.B1(n_983),
.B2(n_982),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_988),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_989),
.B(n_982),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_991),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_993),
.B(n_987),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_990),
.B(n_986),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_994),
.B(n_986),
.Y(n_1001)
);

OAI21xp33_ASAP7_75t_L g1002 ( 
.A1(n_999),
.A2(n_883),
.B(n_882),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_995),
.B(n_925),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_997),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_996),
.B(n_925),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_1000),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_1004),
.B(n_998),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_1006),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_1005),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_1003),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_1002),
.B(n_1001),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_1004),
.B(n_929),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_1009),
.B(n_929),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1008),
.B(n_916),
.Y(n_1014)
);

NOR4xp25_ASAP7_75t_L g1015 ( 
.A(n_1011),
.B(n_780),
.C(n_802),
.D(n_803),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_1010),
.B(n_1007),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_1012),
.A2(n_780),
.B(n_803),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1009),
.B(n_916),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_1016),
.B(n_883),
.Y(n_1019)
);

AOI221xp5_ASAP7_75t_L g1020 ( 
.A1(n_1018),
.A2(n_802),
.B1(n_781),
.B2(n_710),
.C(n_703),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_1013),
.A2(n_745),
.B1(n_917),
.B2(n_908),
.Y(n_1021)
);

AOI221xp5_ASAP7_75t_L g1022 ( 
.A1(n_1014),
.A2(n_719),
.B1(n_717),
.B2(n_703),
.C(n_720),
.Y(n_1022)
);

NAND3xp33_ASAP7_75t_SL g1023 ( 
.A(n_1019),
.B(n_1022),
.C(n_1017),
.Y(n_1023)
);

AOI222xp33_ASAP7_75t_L g1024 ( 
.A1(n_1021),
.A2(n_1015),
.B1(n_792),
.B2(n_844),
.C1(n_717),
.C2(n_719),
.Y(n_1024)
);

NOR3xp33_ASAP7_75t_L g1025 ( 
.A(n_1020),
.B(n_745),
.C(n_724),
.Y(n_1025)
);

NAND4xp25_ASAP7_75t_L g1026 ( 
.A(n_1019),
.B(n_718),
.C(n_855),
.D(n_856),
.Y(n_1026)
);

AOI211xp5_ASAP7_75t_L g1027 ( 
.A1(n_1019),
.A2(n_717),
.B(n_703),
.C(n_719),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_1019),
.Y(n_1028)
);

OAI211xp5_ASAP7_75t_L g1029 ( 
.A1(n_1019),
.A2(n_734),
.B(n_725),
.C(n_897),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_1019),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_1028),
.A2(n_921),
.B(n_858),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1030),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_1023),
.B(n_921),
.Y(n_1033)
);

AOI221xp5_ASAP7_75t_L g1034 ( 
.A1(n_1025),
.A2(n_734),
.B1(n_725),
.B2(n_855),
.C(n_858),
.Y(n_1034)
);

OAI322xp33_ASAP7_75t_L g1035 ( 
.A1(n_1024),
.A2(n_917),
.A3(n_915),
.B1(n_908),
.B2(n_734),
.C1(n_725),
.C2(n_856),
.Y(n_1035)
);

AOI21xp33_ASAP7_75t_SL g1036 ( 
.A1(n_1029),
.A2(n_197),
.B(n_198),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1027),
.B(n_1026),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1028),
.B(n_896),
.Y(n_1038)
);

NOR3xp33_ASAP7_75t_L g1039 ( 
.A(n_1028),
.B(n_847),
.C(n_860),
.Y(n_1039)
);

NOR2x1_ASAP7_75t_L g1040 ( 
.A(n_1030),
.B(n_917),
.Y(n_1040)
);

NAND3x2_ASAP7_75t_L g1041 ( 
.A(n_1033),
.B(n_920),
.C(n_838),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1032),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1038),
.Y(n_1043)
);

AOI211xp5_ASAP7_75t_L g1044 ( 
.A1(n_1036),
.A2(n_866),
.B(n_896),
.C(n_847),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1037),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1034),
.A2(n_847),
.B(n_884),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_1031),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1040),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_1039),
.B(n_794),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_SL g1050 ( 
.A(n_1035),
.B(n_721),
.C(n_915),
.Y(n_1050)
);

NOR3xp33_ASAP7_75t_L g1051 ( 
.A(n_1032),
.B(n_857),
.C(n_860),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_SL g1052 ( 
.A(n_1032),
.B(n_721),
.C(n_890),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1033),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1042),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_1043),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_1045),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_1053),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1047),
.B(n_920),
.Y(n_1058)
);

NAND2xp33_ASAP7_75t_R g1059 ( 
.A(n_1048),
.B(n_199),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1044),
.B(n_1049),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_1049),
.Y(n_1061)
);

NOR2xp67_ASAP7_75t_L g1062 ( 
.A(n_1050),
.B(n_200),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_1059),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1055),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1056),
.A2(n_1052),
.B1(n_1051),
.B2(n_1041),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_1057),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1054),
.A2(n_1046),
.B1(n_896),
.B2(n_870),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1062),
.A2(n_928),
.B1(n_924),
.B2(n_923),
.Y(n_1068)
);

OA21x2_ASAP7_75t_L g1069 ( 
.A1(n_1060),
.A2(n_862),
.B(n_924),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_1063),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1066),
.Y(n_1071)
);

OAI22x1_ASAP7_75t_L g1072 ( 
.A1(n_1065),
.A2(n_1061),
.B1(n_1058),
.B2(n_928),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_1071),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_SL g1074 ( 
.A1(n_1073),
.A2(n_1064),
.B1(n_1070),
.B2(n_1072),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_1074),
.B(n_1067),
.Y(n_1075)
);

OAI222xp33_ASAP7_75t_L g1076 ( 
.A1(n_1075),
.A2(n_1068),
.B1(n_1069),
.B2(n_838),
.C1(n_923),
.C2(n_844),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1075),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1075),
.A2(n_833),
.B1(n_844),
.B2(n_857),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_1077),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1078),
.A2(n_833),
.B1(n_844),
.B2(n_857),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_1076),
.A2(n_857),
.B1(n_860),
.B2(n_845),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1077),
.A2(n_201),
.B(n_203),
.Y(n_1082)
);

AOI222xp33_ASAP7_75t_L g1083 ( 
.A1(n_1079),
.A2(n_846),
.B1(n_845),
.B2(n_842),
.C1(n_205),
.C2(n_206),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_1082),
.A2(n_860),
.B1(n_842),
.B2(n_846),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_SL g1085 ( 
.A1(n_1081),
.A2(n_1080),
.B1(n_211),
.B2(n_899),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1079),
.A2(n_846),
.B1(n_764),
.B2(n_839),
.Y(n_1086)
);

NOR2x1p5_ASAP7_75t_L g1087 ( 
.A(n_1083),
.B(n_835),
.Y(n_1087)
);

OA21x2_ASAP7_75t_L g1088 ( 
.A1(n_1084),
.A2(n_862),
.B(n_861),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1087),
.A2(n_1086),
.B1(n_1085),
.B2(n_839),
.Y(n_1089)
);

AOI211xp5_ASAP7_75t_L g1090 ( 
.A1(n_1089),
.A2(n_1088),
.B(n_862),
.C(n_841),
.Y(n_1090)
);


endmodule