module fake_netlist_5_468_n_6187 (n_924, n_1263, n_977, n_1378, n_611, n_1126, n_1423, n_1729, n_1166, n_1751, n_469, n_1508, n_82, n_785, n_549, n_532, n_1161, n_1677, n_1150, n_226, n_1780, n_1488, n_667, n_790, n_1055, n_1501, n_111, n_880, n_544, n_1007, n_155, n_552, n_1528, n_1370, n_1292, n_1198, n_1360, n_1099, n_956, n_564, n_423, n_1738, n_21, n_105, n_1021, n_4, n_551, n_1323, n_1466, n_688, n_1695, n_1353, n_800, n_1347, n_1535, n_1789, n_1666, n_671, n_819, n_1451, n_1022, n_915, n_1545, n_864, n_173, n_859, n_951, n_1264, n_447, n_247, n_1494, n_292, n_625, n_854, n_1462, n_1580, n_674, n_417, n_516, n_933, n_1152, n_497, n_1607, n_1563, n_606, n_275, n_26, n_877, n_2, n_1696, n_755, n_1118, n_6, n_1686, n_947, n_1285, n_373, n_307, n_1359, n_530, n_87, n_150, n_1107, n_1728, n_556, n_1230, n_668, n_375, n_301, n_929, n_1124, n_902, n_1576, n_191, n_1104, n_1294, n_659, n_51, n_1705, n_1257, n_171, n_1182, n_579, n_1698, n_1261, n_938, n_1098, n_320, n_1154, n_1242, n_1135, n_24, n_406, n_519, n_1016, n_1243, n_546, n_101, n_1280, n_281, n_240, n_291, n_231, n_257, n_731, n_371, n_1483, n_1314, n_1512, n_709, n_1490, n_317, n_1236, n_1633, n_569, n_1778, n_227, n_920, n_1289, n_1517, n_94, n_335, n_1669, n_370, n_976, n_343, n_1449, n_308, n_1566, n_297, n_156, n_1078, n_1670, n_775, n_219, n_157, n_600, n_1484, n_1374, n_1328, n_223, n_264, n_1598, n_1723, n_955, n_163, n_339, n_1146, n_882, n_183, n_243, n_1036, n_1097, n_1749, n_347, n_59, n_550, n_696, n_897, n_215, n_350, n_196, n_798, n_646, n_1428, n_436, n_1394, n_1414, n_1216, n_290, n_580, n_1040, n_578, n_926, n_344, n_1218, n_422, n_475, n_777, n_1070, n_1547, n_1030, n_72, n_1755, n_415, n_1071, n_485, n_1165, n_1267, n_1561, n_496, n_1391, n_958, n_1034, n_670, n_1513, n_1600, n_48, n_521, n_663, n_845, n_673, n_837, n_1239, n_528, n_1796, n_680, n_1473, n_1587, n_395, n_164, n_553, n_901, n_813, n_1521, n_1284, n_1590, n_214, n_1748, n_1672, n_675, n_888, n_1167, n_1626, n_637, n_1384, n_1556, n_184, n_446, n_1064, n_144, n_858, n_114, n_96, n_923, n_691, n_1151, n_881, n_1405, n_1706, n_468, n_213, n_129, n_342, n_464, n_363, n_1582, n_197, n_1069, n_1784, n_1075, n_1450, n_1322, n_1471, n_1750, n_1459, n_460, n_889, n_973, n_1700, n_477, n_571, n_1585, n_461, n_1599, n_1211, n_1197, n_1523, n_907, n_1447, n_1377, n_190, n_989, n_1039, n_34, n_228, n_283, n_1403, n_488, n_736, n_892, n_1000, n_1202, n_1278, n_1002, n_1463, n_1581, n_49, n_310, n_54, n_593, n_12, n_748, n_586, n_1058, n_1667, n_838, n_332, n_1053, n_1224, n_349, n_1248, n_230, n_1331, n_953, n_279, n_1014, n_1241, n_70, n_289, n_963, n_1052, n_954, n_627, n_1385, n_440, n_793, n_478, n_476, n_1527, n_534, n_884, n_345, n_944, n_1754, n_1623, n_91, n_1565, n_182, n_143, n_647, n_237, n_407, n_1072, n_832, n_857, n_207, n_561, n_1319, n_1712, n_1387, n_1532, n_18, n_1027, n_971, n_1156, n_117, n_326, n_794, n_404, n_686, n_847, n_1393, n_596, n_1775, n_1368, n_558, n_702, n_1276, n_822, n_1412, n_1709, n_728, n_266, n_1162, n_272, n_1538, n_1199, n_1779, n_352, n_53, n_1038, n_520, n_1369, n_409, n_1660, n_887, n_154, n_71, n_300, n_809, n_870, n_931, n_599, n_1711, n_1662, n_1481, n_434, n_1544, n_868, n_639, n_914, n_411, n_414, n_1629, n_1293, n_965, n_1743, n_935, n_121, n_1175, n_817, n_360, n_36, n_1479, n_64, n_759, n_28, n_806, n_1766, n_1477, n_324, n_1635, n_1571, n_187, n_1189, n_103, n_97, n_11, n_7, n_1259, n_1690, n_706, n_746, n_1649, n_747, n_52, n_784, n_110, n_1733, n_1244, n_431, n_1194, n_615, n_851, n_1759, n_843, n_1788, n_523, n_913, n_1537, n_705, n_865, n_61, n_678, n_697, n_127, n_1222, n_75, n_1679, n_776, n_1790, n_1415, n_367, n_452, n_525, n_1260, n_1746, n_1647, n_1464, n_649, n_547, n_43, n_1444, n_1191, n_1674, n_116, n_1710, n_284, n_1128, n_139, n_1734, n_744, n_590, n_629, n_1308, n_1767, n_254, n_1680, n_1233, n_23, n_1615, n_1529, n_526, n_293, n_372, n_677, n_244, n_47, n_1333, n_1121, n_314, n_368, n_433, n_604, n_8, n_949, n_100, n_1443, n_1008, n_946, n_1539, n_1001, n_1503, n_498, n_1468, n_1559, n_1765, n_689, n_738, n_1624, n_640, n_1510, n_252, n_624, n_1380, n_1744, n_1617, n_295, n_133, n_1010, n_1231, n_739, n_1279, n_1406, n_1195, n_610, n_1760, n_936, n_568, n_1500, n_39, n_1090, n_757, n_633, n_439, n_106, n_259, n_448, n_758, n_999, n_93, n_1656, n_1158, n_1509, n_563, n_1145, n_878, n_524, n_204, n_394, n_1678, n_1049, n_1153, n_741, n_1639, n_1306, n_1068, n_122, n_331, n_10, n_906, n_1163, n_1207, n_919, n_908, n_90, n_724, n_1781, n_658, n_1740, n_1362, n_1586, n_456, n_959, n_535, n_152, n_940, n_1445, n_9, n_1492, n_1773, n_592, n_1169, n_45, n_1596, n_1692, n_1017, n_123, n_978, n_1434, n_1054, n_1474, n_1665, n_1269, n_1095, n_1614, n_267, n_514, n_457, n_1079, n_1045, n_1208, n_603, n_1431, n_484, n_1593, n_1033, n_442, n_131, n_636, n_660, n_1640, n_1732, n_1009, n_1148, n_109, n_742, n_750, n_995, n_454, n_1609, n_374, n_185, n_396, n_1383, n_1073, n_255, n_662, n_459, n_218, n_962, n_1215, n_1171, n_1578, n_723, n_1065, n_1592, n_1336, n_1721, n_1758, n_1574, n_473, n_1309, n_1426, n_1043, n_355, n_486, n_1548, n_614, n_337, n_1421, n_88, n_1286, n_1177, n_1355, n_168, n_974, n_727, n_1159, n_957, n_773, n_208, n_142, n_743, n_299, n_303, n_296, n_613, n_1119, n_1240, n_65, n_829, n_1612, n_1416, n_1724, n_361, n_700, n_1237, n_573, n_69, n_1420, n_1132, n_388, n_1366, n_1300, n_1127, n_761, n_1785, n_1568, n_1006, n_329, n_274, n_1270, n_1664, n_1486, n_582, n_1332, n_1390, n_73, n_19, n_309, n_30, n_512, n_1591, n_84, n_130, n_322, n_1682, n_1249, n_652, n_1111, n_1365, n_25, n_1349, n_1093, n_288, n_1031, n_263, n_609, n_1041, n_1265, n_44, n_224, n_1562, n_383, n_834, n_112, n_765, n_893, n_1015, n_1140, n_891, n_1651, n_239, n_630, n_55, n_504, n_511, n_874, n_358, n_1101, n_77, n_102, n_1106, n_1456, n_1304, n_1324, n_987, n_261, n_174, n_1455, n_767, n_993, n_1407, n_1551, n_545, n_441, n_860, n_450, n_429, n_948, n_1217, n_628, n_365, n_729, n_1131, n_1084, n_970, n_911, n_1430, n_83, n_513, n_1094, n_1354, n_560, n_1534, n_340, n_1351, n_1044, n_1205, n_346, n_1209, n_1552, n_495, n_602, n_574, n_1435, n_879, n_16, n_58, n_623, n_405, n_824, n_359, n_1645, n_490, n_1327, n_996, n_921, n_1684, n_233, n_1717, n_572, n_366, n_815, n_1795, n_128, n_120, n_327, n_135, n_1381, n_1611, n_1037, n_1080, n_1274, n_1316, n_1708, n_426, n_1438, n_1082, n_589, n_716, n_1630, n_562, n_1436, n_62, n_1691, n_952, n_1229, n_391, n_701, n_1437, n_1023, n_645, n_539, n_803, n_1092, n_238, n_1776, n_531, n_1757, n_890, n_764, n_1056, n_1424, n_162, n_960, n_222, n_1290, n_1123, n_1467, n_1047, n_634, n_199, n_32, n_1252, n_348, n_1382, n_1029, n_925, n_1206, n_424, n_1311, n_1519, n_256, n_950, n_1553, n_380, n_419, n_1346, n_444, n_1299, n_1060, n_1141, n_316, n_389, n_418, n_248, n_136, n_86, n_146, n_912, n_315, n_968, n_451, n_619, n_408, n_1386, n_1699, n_376, n_967, n_1442, n_74, n_1139, n_515, n_57, n_351, n_885, n_397, n_1432, n_1357, n_483, n_683, n_1632, n_1057, n_1051, n_1085, n_1066, n_721, n_1157, n_841, n_1050, n_22, n_802, n_46, n_1608, n_983, n_38, n_280, n_1305, n_873, n_378, n_1112, n_762, n_1283, n_1644, n_17, n_690, n_33, n_583, n_302, n_1343, n_1203, n_1631, n_821, n_1763, n_1768, n_321, n_1179, n_621, n_753, n_455, n_1048, n_1719, n_1288, n_212, n_385, n_507, n_1560, n_1605, n_330, n_1228, n_972, n_692, n_820, n_1200, n_1301, n_1363, n_1668, n_1185, n_991, n_828, n_779, n_576, n_1143, n_1579, n_1329, n_1312, n_1439, n_804, n_537, n_1688, n_945, n_492, n_153, n_1504, n_943, n_341, n_250, n_992, n_543, n_260, n_842, n_650, n_984, n_694, n_286, n_1643, n_883, n_470, n_325, n_449, n_1594, n_132, n_1214, n_1342, n_1400, n_900, n_856, n_1793, n_918, n_942, n_189, n_1147, n_1557, n_1610, n_13, n_1077, n_1422, n_540, n_618, n_896, n_323, n_195, n_356, n_894, n_1636, n_1730, n_831, n_964, n_1373, n_1350, n_1511, n_1470, n_1096, n_234, n_1575, n_1697, n_1735, n_833, n_5, n_1646, n_225, n_1307, n_988, n_814, n_192, n_1549, n_1201, n_1114, n_655, n_1616, n_1446, n_669, n_472, n_1458, n_1176, n_1472, n_387, n_1149, n_398, n_1671, n_635, n_763, n_1020, n_1062, n_211, n_1219, n_3, n_1204, n_178, n_1035, n_287, n_555, n_783, n_1188, n_1722, n_661, n_41, n_849, n_15, n_336, n_584, n_681, n_1638, n_1786, n_50, n_430, n_510, n_216, n_311, n_830, n_1296, n_1413, n_801, n_241, n_875, n_357, n_1110, n_1655, n_445, n_749, n_1134, n_1358, n_717, n_165, n_939, n_482, n_1088, n_588, n_1173, n_789, n_1232, n_1603, n_734, n_638, n_866, n_107, n_969, n_1401, n_1019, n_1105, n_249, n_304, n_1338, n_577, n_1522, n_1687, n_1637, n_1419, n_338, n_149, n_1653, n_693, n_1506, n_14, n_836, n_990, n_1389, n_975, n_1256, n_1702, n_567, n_1465, n_778, n_1122, n_151, n_306, n_458, n_770, n_1375, n_1102, n_711, n_1499, n_85, n_1187, n_1441, n_1392, n_1597, n_1164, n_1659, n_489, n_1174, n_1371, n_617, n_1303, n_1572, n_876, n_1516, n_1190, n_1736, n_1685, n_118, n_601, n_917, n_1714, n_966, n_253, n_1116, n_1661, n_1212, n_1541, n_172, n_206, n_217, n_726, n_982, n_1573, n_1453, n_1731, n_818, n_861, n_1713, n_1183, n_1658, n_899, n_1253, n_210, n_1737, n_774, n_1628, n_1335, n_1514, n_1777, n_1059, n_1345, n_176, n_1133, n_1771, n_557, n_1410, n_1005, n_607, n_1003, n_679, n_710, n_527, n_1168, n_707, n_937, n_1427, n_393, n_108, n_487, n_1584, n_665, n_1726, n_66, n_1440, n_177, n_421, n_1356, n_1787, n_910, n_1657, n_768, n_1475, n_1302, n_1774, n_1725, n_205, n_1136, n_1313, n_1491, n_754, n_1496, n_179, n_1125, n_125, n_410, n_708, n_529, n_735, n_232, n_1109, n_126, n_895, n_1310, n_202, n_427, n_1399, n_1543, n_791, n_732, n_1533, n_193, n_808, n_797, n_1025, n_500, n_1067, n_1720, n_148, n_435, n_159, n_766, n_1457, n_541, n_538, n_1117, n_799, n_687, n_715, n_1742, n_1480, n_1482, n_1213, n_1266, n_536, n_872, n_594, n_200, n_1291, n_1297, n_1753, n_1782, n_1155, n_1418, n_89, n_1524, n_1689, n_1485, n_115, n_1011, n_1184, n_985, n_869, n_810, n_416, n_827, n_401, n_1703, n_1352, n_626, n_1650, n_1144, n_1137, n_1570, n_1170, n_305, n_137, n_676, n_294, n_318, n_653, n_642, n_1602, n_194, n_855, n_1178, n_1461, n_850, n_684, n_124, n_268, n_664, n_503, n_235, n_1372, n_605, n_1273, n_353, n_620, n_643, n_916, n_1081, n_493, n_1235, n_703, n_698, n_980, n_1115, n_1282, n_1318, n_1783, n_780, n_998, n_1454, n_467, n_1227, n_1531, n_840, n_1334, n_501, n_823, n_245, n_725, n_1388, n_1417, n_1295, n_672, n_581, n_382, n_554, n_1625, n_898, n_1762, n_1013, n_1452, n_718, n_265, n_1120, n_719, n_443, n_1791, n_198, n_1747, n_714, n_1683, n_909, n_1497, n_1530, n_997, n_932, n_612, n_1409, n_788, n_1326, n_119, n_1268, n_559, n_825, n_508, n_506, n_1320, n_1663, n_737, n_1718, n_986, n_509, n_1317, n_147, n_1518, n_1715, n_1281, n_67, n_1192, n_1024, n_1063, n_209, n_1792, n_1564, n_1613, n_733, n_1489, n_1376, n_941, n_981, n_1569, n_68, n_867, n_186, n_134, n_587, n_63, n_792, n_756, n_1429, n_399, n_1238, n_548, n_812, n_298, n_518, n_505, n_1772, n_282, n_752, n_905, n_1476, n_1108, n_782, n_1100, n_1395, n_862, n_1425, n_760, n_1620, n_381, n_220, n_390, n_1330, n_31, n_481, n_1675, n_1727, n_1554, n_1745, n_769, n_42, n_1046, n_271, n_934, n_1618, n_826, n_886, n_1221, n_654, n_1172, n_167, n_379, n_428, n_1341, n_570, n_1641, n_1361, n_1707, n_853, n_377, n_751, n_786, n_1083, n_1142, n_1129, n_392, n_158, n_704, n_787, n_1770, n_138, n_961, n_1756, n_771, n_276, n_95, n_1716, n_1225, n_1520, n_169, n_522, n_1287, n_1262, n_400, n_930, n_181, n_1411, n_221, n_622, n_1577, n_1087, n_386, n_994, n_1701, n_848, n_1550, n_1498, n_1223, n_1272, n_104, n_682, n_1567, n_56, n_141, n_1247, n_922, n_816, n_1648, n_591, n_145, n_1536, n_1344, n_313, n_631, n_479, n_1246, n_1339, n_1478, n_432, n_1769, n_839, n_1210, n_1364, n_328, n_140, n_1250, n_369, n_871, n_598, n_685, n_928, n_608, n_1367, n_78, n_1460, n_772, n_1555, n_499, n_1589, n_517, n_98, n_402, n_413, n_1086, n_796, n_1619, n_236, n_1502, n_1469, n_1012, n_1, n_1396, n_1348, n_903, n_1525, n_1752, n_740, n_203, n_384, n_1404, n_80, n_1794, n_35, n_1315, n_277, n_1061, n_92, n_333, n_1298, n_1652, n_462, n_1193, n_1676, n_1255, n_258, n_1113, n_29, n_79, n_1226, n_722, n_1277, n_188, n_844, n_201, n_471, n_852, n_1487, n_40, n_1028, n_1601, n_781, n_474, n_542, n_463, n_1546, n_595, n_502, n_466, n_420, n_1337, n_1495, n_632, n_699, n_979, n_1515, n_1627, n_1245, n_846, n_1673, n_465, n_76, n_362, n_1321, n_170, n_27, n_161, n_273, n_585, n_1739, n_270, n_616, n_81, n_745, n_1654, n_1103, n_648, n_1379, n_312, n_1076, n_1091, n_1408, n_494, n_1761, n_641, n_730, n_1325, n_1595, n_354, n_575, n_480, n_425, n_795, n_695, n_180, n_656, n_1606, n_1220, n_37, n_1694, n_1540, n_229, n_437, n_1642, n_60, n_403, n_453, n_1130, n_720, n_0, n_1526, n_863, n_805, n_1604, n_1275, n_1764, n_113, n_712, n_246, n_1583, n_1042, n_1402, n_269, n_285, n_412, n_1493, n_657, n_644, n_1741, n_1160, n_1397, n_491, n_1258, n_1074, n_1621, n_251, n_160, n_566, n_565, n_1448, n_1507, n_1398, n_597, n_1181, n_1505, n_1634, n_1196, n_651, n_1340, n_334, n_811, n_1558, n_807, n_835, n_175, n_666, n_262, n_1433, n_1704, n_99, n_1254, n_1026, n_1234, n_319, n_364, n_1138, n_927, n_20, n_1089, n_1004, n_1186, n_1032, n_242, n_1681, n_1018, n_1693, n_438, n_713, n_904, n_1588, n_1622, n_166, n_1180, n_1271, n_533, n_1542, n_1251, n_278, n_6187);

input n_924;
input n_1263;
input n_977;
input n_1378;
input n_611;
input n_1126;
input n_1423;
input n_1729;
input n_1166;
input n_1751;
input n_469;
input n_1508;
input n_82;
input n_785;
input n_549;
input n_532;
input n_1161;
input n_1677;
input n_1150;
input n_226;
input n_1780;
input n_1488;
input n_667;
input n_790;
input n_1055;
input n_1501;
input n_111;
input n_880;
input n_544;
input n_1007;
input n_155;
input n_552;
input n_1528;
input n_1370;
input n_1292;
input n_1198;
input n_1360;
input n_1099;
input n_956;
input n_564;
input n_423;
input n_1738;
input n_21;
input n_105;
input n_1021;
input n_4;
input n_551;
input n_1323;
input n_1466;
input n_688;
input n_1695;
input n_1353;
input n_800;
input n_1347;
input n_1535;
input n_1789;
input n_1666;
input n_671;
input n_819;
input n_1451;
input n_1022;
input n_915;
input n_1545;
input n_864;
input n_173;
input n_859;
input n_951;
input n_1264;
input n_447;
input n_247;
input n_1494;
input n_292;
input n_625;
input n_854;
input n_1462;
input n_1580;
input n_674;
input n_417;
input n_516;
input n_933;
input n_1152;
input n_497;
input n_1607;
input n_1563;
input n_606;
input n_275;
input n_26;
input n_877;
input n_2;
input n_1696;
input n_755;
input n_1118;
input n_6;
input n_1686;
input n_947;
input n_1285;
input n_373;
input n_307;
input n_1359;
input n_530;
input n_87;
input n_150;
input n_1107;
input n_1728;
input n_556;
input n_1230;
input n_668;
input n_375;
input n_301;
input n_929;
input n_1124;
input n_902;
input n_1576;
input n_191;
input n_1104;
input n_1294;
input n_659;
input n_51;
input n_1705;
input n_1257;
input n_171;
input n_1182;
input n_579;
input n_1698;
input n_1261;
input n_938;
input n_1098;
input n_320;
input n_1154;
input n_1242;
input n_1135;
input n_24;
input n_406;
input n_519;
input n_1016;
input n_1243;
input n_546;
input n_101;
input n_1280;
input n_281;
input n_240;
input n_291;
input n_231;
input n_257;
input n_731;
input n_371;
input n_1483;
input n_1314;
input n_1512;
input n_709;
input n_1490;
input n_317;
input n_1236;
input n_1633;
input n_569;
input n_1778;
input n_227;
input n_920;
input n_1289;
input n_1517;
input n_94;
input n_335;
input n_1669;
input n_370;
input n_976;
input n_343;
input n_1449;
input n_308;
input n_1566;
input n_297;
input n_156;
input n_1078;
input n_1670;
input n_775;
input n_219;
input n_157;
input n_600;
input n_1484;
input n_1374;
input n_1328;
input n_223;
input n_264;
input n_1598;
input n_1723;
input n_955;
input n_163;
input n_339;
input n_1146;
input n_882;
input n_183;
input n_243;
input n_1036;
input n_1097;
input n_1749;
input n_347;
input n_59;
input n_550;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_646;
input n_1428;
input n_436;
input n_1394;
input n_1414;
input n_1216;
input n_290;
input n_580;
input n_1040;
input n_578;
input n_926;
input n_344;
input n_1218;
input n_422;
input n_475;
input n_777;
input n_1070;
input n_1547;
input n_1030;
input n_72;
input n_1755;
input n_415;
input n_1071;
input n_485;
input n_1165;
input n_1267;
input n_1561;
input n_496;
input n_1391;
input n_958;
input n_1034;
input n_670;
input n_1513;
input n_1600;
input n_48;
input n_521;
input n_663;
input n_845;
input n_673;
input n_837;
input n_1239;
input n_528;
input n_1796;
input n_680;
input n_1473;
input n_1587;
input n_395;
input n_164;
input n_553;
input n_901;
input n_813;
input n_1521;
input n_1284;
input n_1590;
input n_214;
input n_1748;
input n_1672;
input n_675;
input n_888;
input n_1167;
input n_1626;
input n_637;
input n_1384;
input n_1556;
input n_184;
input n_446;
input n_1064;
input n_144;
input n_858;
input n_114;
input n_96;
input n_923;
input n_691;
input n_1151;
input n_881;
input n_1405;
input n_1706;
input n_468;
input n_213;
input n_129;
input n_342;
input n_464;
input n_363;
input n_1582;
input n_197;
input n_1069;
input n_1784;
input n_1075;
input n_1450;
input n_1322;
input n_1471;
input n_1750;
input n_1459;
input n_460;
input n_889;
input n_973;
input n_1700;
input n_477;
input n_571;
input n_1585;
input n_461;
input n_1599;
input n_1211;
input n_1197;
input n_1523;
input n_907;
input n_1447;
input n_1377;
input n_190;
input n_989;
input n_1039;
input n_34;
input n_228;
input n_283;
input n_1403;
input n_488;
input n_736;
input n_892;
input n_1000;
input n_1202;
input n_1278;
input n_1002;
input n_1463;
input n_1581;
input n_49;
input n_310;
input n_54;
input n_593;
input n_12;
input n_748;
input n_586;
input n_1058;
input n_1667;
input n_838;
input n_332;
input n_1053;
input n_1224;
input n_349;
input n_1248;
input n_230;
input n_1331;
input n_953;
input n_279;
input n_1014;
input n_1241;
input n_70;
input n_289;
input n_963;
input n_1052;
input n_954;
input n_627;
input n_1385;
input n_440;
input n_793;
input n_478;
input n_476;
input n_1527;
input n_534;
input n_884;
input n_345;
input n_944;
input n_1754;
input n_1623;
input n_91;
input n_1565;
input n_182;
input n_143;
input n_647;
input n_237;
input n_407;
input n_1072;
input n_832;
input n_857;
input n_207;
input n_561;
input n_1319;
input n_1712;
input n_1387;
input n_1532;
input n_18;
input n_1027;
input n_971;
input n_1156;
input n_117;
input n_326;
input n_794;
input n_404;
input n_686;
input n_847;
input n_1393;
input n_596;
input n_1775;
input n_1368;
input n_558;
input n_702;
input n_1276;
input n_822;
input n_1412;
input n_1709;
input n_728;
input n_266;
input n_1162;
input n_272;
input n_1538;
input n_1199;
input n_1779;
input n_352;
input n_53;
input n_1038;
input n_520;
input n_1369;
input n_409;
input n_1660;
input n_887;
input n_154;
input n_71;
input n_300;
input n_809;
input n_870;
input n_931;
input n_599;
input n_1711;
input n_1662;
input n_1481;
input n_434;
input n_1544;
input n_868;
input n_639;
input n_914;
input n_411;
input n_414;
input n_1629;
input n_1293;
input n_965;
input n_1743;
input n_935;
input n_121;
input n_1175;
input n_817;
input n_360;
input n_36;
input n_1479;
input n_64;
input n_759;
input n_28;
input n_806;
input n_1766;
input n_1477;
input n_324;
input n_1635;
input n_1571;
input n_187;
input n_1189;
input n_103;
input n_97;
input n_11;
input n_7;
input n_1259;
input n_1690;
input n_706;
input n_746;
input n_1649;
input n_747;
input n_52;
input n_784;
input n_110;
input n_1733;
input n_1244;
input n_431;
input n_1194;
input n_615;
input n_851;
input n_1759;
input n_843;
input n_1788;
input n_523;
input n_913;
input n_1537;
input n_705;
input n_865;
input n_61;
input n_678;
input n_697;
input n_127;
input n_1222;
input n_75;
input n_1679;
input n_776;
input n_1790;
input n_1415;
input n_367;
input n_452;
input n_525;
input n_1260;
input n_1746;
input n_1647;
input n_1464;
input n_649;
input n_547;
input n_43;
input n_1444;
input n_1191;
input n_1674;
input n_116;
input n_1710;
input n_284;
input n_1128;
input n_139;
input n_1734;
input n_744;
input n_590;
input n_629;
input n_1308;
input n_1767;
input n_254;
input n_1680;
input n_1233;
input n_23;
input n_1615;
input n_1529;
input n_526;
input n_293;
input n_372;
input n_677;
input n_244;
input n_47;
input n_1333;
input n_1121;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_949;
input n_100;
input n_1443;
input n_1008;
input n_946;
input n_1539;
input n_1001;
input n_1503;
input n_498;
input n_1468;
input n_1559;
input n_1765;
input n_689;
input n_738;
input n_1624;
input n_640;
input n_1510;
input n_252;
input n_624;
input n_1380;
input n_1744;
input n_1617;
input n_295;
input n_133;
input n_1010;
input n_1231;
input n_739;
input n_1279;
input n_1406;
input n_1195;
input n_610;
input n_1760;
input n_936;
input n_568;
input n_1500;
input n_39;
input n_1090;
input n_757;
input n_633;
input n_439;
input n_106;
input n_259;
input n_448;
input n_758;
input n_999;
input n_93;
input n_1656;
input n_1158;
input n_1509;
input n_563;
input n_1145;
input n_878;
input n_524;
input n_204;
input n_394;
input n_1678;
input n_1049;
input n_1153;
input n_741;
input n_1639;
input n_1306;
input n_1068;
input n_122;
input n_331;
input n_10;
input n_906;
input n_1163;
input n_1207;
input n_919;
input n_908;
input n_90;
input n_724;
input n_1781;
input n_658;
input n_1740;
input n_1362;
input n_1586;
input n_456;
input n_959;
input n_535;
input n_152;
input n_940;
input n_1445;
input n_9;
input n_1492;
input n_1773;
input n_592;
input n_1169;
input n_45;
input n_1596;
input n_1692;
input n_1017;
input n_123;
input n_978;
input n_1434;
input n_1054;
input n_1474;
input n_1665;
input n_1269;
input n_1095;
input n_1614;
input n_267;
input n_514;
input n_457;
input n_1079;
input n_1045;
input n_1208;
input n_603;
input n_1431;
input n_484;
input n_1593;
input n_1033;
input n_442;
input n_131;
input n_636;
input n_660;
input n_1640;
input n_1732;
input n_1009;
input n_1148;
input n_109;
input n_742;
input n_750;
input n_995;
input n_454;
input n_1609;
input n_374;
input n_185;
input n_396;
input n_1383;
input n_1073;
input n_255;
input n_662;
input n_459;
input n_218;
input n_962;
input n_1215;
input n_1171;
input n_1578;
input n_723;
input n_1065;
input n_1592;
input n_1336;
input n_1721;
input n_1758;
input n_1574;
input n_473;
input n_1309;
input n_1426;
input n_1043;
input n_355;
input n_486;
input n_1548;
input n_614;
input n_337;
input n_1421;
input n_88;
input n_1286;
input n_1177;
input n_1355;
input n_168;
input n_974;
input n_727;
input n_1159;
input n_957;
input n_773;
input n_208;
input n_142;
input n_743;
input n_299;
input n_303;
input n_296;
input n_613;
input n_1119;
input n_1240;
input n_65;
input n_829;
input n_1612;
input n_1416;
input n_1724;
input n_361;
input n_700;
input n_1237;
input n_573;
input n_69;
input n_1420;
input n_1132;
input n_388;
input n_1366;
input n_1300;
input n_1127;
input n_761;
input n_1785;
input n_1568;
input n_1006;
input n_329;
input n_274;
input n_1270;
input n_1664;
input n_1486;
input n_582;
input n_1332;
input n_1390;
input n_73;
input n_19;
input n_309;
input n_30;
input n_512;
input n_1591;
input n_84;
input n_130;
input n_322;
input n_1682;
input n_1249;
input n_652;
input n_1111;
input n_1365;
input n_25;
input n_1349;
input n_1093;
input n_288;
input n_1031;
input n_263;
input n_609;
input n_1041;
input n_1265;
input n_44;
input n_224;
input n_1562;
input n_383;
input n_834;
input n_112;
input n_765;
input n_893;
input n_1015;
input n_1140;
input n_891;
input n_1651;
input n_239;
input n_630;
input n_55;
input n_504;
input n_511;
input n_874;
input n_358;
input n_1101;
input n_77;
input n_102;
input n_1106;
input n_1456;
input n_1304;
input n_1324;
input n_987;
input n_261;
input n_174;
input n_1455;
input n_767;
input n_993;
input n_1407;
input n_1551;
input n_545;
input n_441;
input n_860;
input n_450;
input n_429;
input n_948;
input n_1217;
input n_628;
input n_365;
input n_729;
input n_1131;
input n_1084;
input n_970;
input n_911;
input n_1430;
input n_83;
input n_513;
input n_1094;
input n_1354;
input n_560;
input n_1534;
input n_340;
input n_1351;
input n_1044;
input n_1205;
input n_346;
input n_1209;
input n_1552;
input n_495;
input n_602;
input n_574;
input n_1435;
input n_879;
input n_16;
input n_58;
input n_623;
input n_405;
input n_824;
input n_359;
input n_1645;
input n_490;
input n_1327;
input n_996;
input n_921;
input n_1684;
input n_233;
input n_1717;
input n_572;
input n_366;
input n_815;
input n_1795;
input n_128;
input n_120;
input n_327;
input n_135;
input n_1381;
input n_1611;
input n_1037;
input n_1080;
input n_1274;
input n_1316;
input n_1708;
input n_426;
input n_1438;
input n_1082;
input n_589;
input n_716;
input n_1630;
input n_562;
input n_1436;
input n_62;
input n_1691;
input n_952;
input n_1229;
input n_391;
input n_701;
input n_1437;
input n_1023;
input n_645;
input n_539;
input n_803;
input n_1092;
input n_238;
input n_1776;
input n_531;
input n_1757;
input n_890;
input n_764;
input n_1056;
input n_1424;
input n_162;
input n_960;
input n_222;
input n_1290;
input n_1123;
input n_1467;
input n_1047;
input n_634;
input n_199;
input n_32;
input n_1252;
input n_348;
input n_1382;
input n_1029;
input n_925;
input n_1206;
input n_424;
input n_1311;
input n_1519;
input n_256;
input n_950;
input n_1553;
input n_380;
input n_419;
input n_1346;
input n_444;
input n_1299;
input n_1060;
input n_1141;
input n_316;
input n_389;
input n_418;
input n_248;
input n_136;
input n_86;
input n_146;
input n_912;
input n_315;
input n_968;
input n_451;
input n_619;
input n_408;
input n_1386;
input n_1699;
input n_376;
input n_967;
input n_1442;
input n_74;
input n_1139;
input n_515;
input n_57;
input n_351;
input n_885;
input n_397;
input n_1432;
input n_1357;
input n_483;
input n_683;
input n_1632;
input n_1057;
input n_1051;
input n_1085;
input n_1066;
input n_721;
input n_1157;
input n_841;
input n_1050;
input n_22;
input n_802;
input n_46;
input n_1608;
input n_983;
input n_38;
input n_280;
input n_1305;
input n_873;
input n_378;
input n_1112;
input n_762;
input n_1283;
input n_1644;
input n_17;
input n_690;
input n_33;
input n_583;
input n_302;
input n_1343;
input n_1203;
input n_1631;
input n_821;
input n_1763;
input n_1768;
input n_321;
input n_1179;
input n_621;
input n_753;
input n_455;
input n_1048;
input n_1719;
input n_1288;
input n_212;
input n_385;
input n_507;
input n_1560;
input n_1605;
input n_330;
input n_1228;
input n_972;
input n_692;
input n_820;
input n_1200;
input n_1301;
input n_1363;
input n_1668;
input n_1185;
input n_991;
input n_828;
input n_779;
input n_576;
input n_1143;
input n_1579;
input n_1329;
input n_1312;
input n_1439;
input n_804;
input n_537;
input n_1688;
input n_945;
input n_492;
input n_153;
input n_1504;
input n_943;
input n_341;
input n_250;
input n_992;
input n_543;
input n_260;
input n_842;
input n_650;
input n_984;
input n_694;
input n_286;
input n_1643;
input n_883;
input n_470;
input n_325;
input n_449;
input n_1594;
input n_132;
input n_1214;
input n_1342;
input n_1400;
input n_900;
input n_856;
input n_1793;
input n_918;
input n_942;
input n_189;
input n_1147;
input n_1557;
input n_1610;
input n_13;
input n_1077;
input n_1422;
input n_540;
input n_618;
input n_896;
input n_323;
input n_195;
input n_356;
input n_894;
input n_1636;
input n_1730;
input n_831;
input n_964;
input n_1373;
input n_1350;
input n_1511;
input n_1470;
input n_1096;
input n_234;
input n_1575;
input n_1697;
input n_1735;
input n_833;
input n_5;
input n_1646;
input n_225;
input n_1307;
input n_988;
input n_814;
input n_192;
input n_1549;
input n_1201;
input n_1114;
input n_655;
input n_1616;
input n_1446;
input n_669;
input n_472;
input n_1458;
input n_1176;
input n_1472;
input n_387;
input n_1149;
input n_398;
input n_1671;
input n_635;
input n_763;
input n_1020;
input n_1062;
input n_211;
input n_1219;
input n_3;
input n_1204;
input n_178;
input n_1035;
input n_287;
input n_555;
input n_783;
input n_1188;
input n_1722;
input n_661;
input n_41;
input n_849;
input n_15;
input n_336;
input n_584;
input n_681;
input n_1638;
input n_1786;
input n_50;
input n_430;
input n_510;
input n_216;
input n_311;
input n_830;
input n_1296;
input n_1413;
input n_801;
input n_241;
input n_875;
input n_357;
input n_1110;
input n_1655;
input n_445;
input n_749;
input n_1134;
input n_1358;
input n_717;
input n_165;
input n_939;
input n_482;
input n_1088;
input n_588;
input n_1173;
input n_789;
input n_1232;
input n_1603;
input n_734;
input n_638;
input n_866;
input n_107;
input n_969;
input n_1401;
input n_1019;
input n_1105;
input n_249;
input n_304;
input n_1338;
input n_577;
input n_1522;
input n_1687;
input n_1637;
input n_1419;
input n_338;
input n_149;
input n_1653;
input n_693;
input n_1506;
input n_14;
input n_836;
input n_990;
input n_1389;
input n_975;
input n_1256;
input n_1702;
input n_567;
input n_1465;
input n_778;
input n_1122;
input n_151;
input n_306;
input n_458;
input n_770;
input n_1375;
input n_1102;
input n_711;
input n_1499;
input n_85;
input n_1187;
input n_1441;
input n_1392;
input n_1597;
input n_1164;
input n_1659;
input n_489;
input n_1174;
input n_1371;
input n_617;
input n_1303;
input n_1572;
input n_876;
input n_1516;
input n_1190;
input n_1736;
input n_1685;
input n_118;
input n_601;
input n_917;
input n_1714;
input n_966;
input n_253;
input n_1116;
input n_1661;
input n_1212;
input n_1541;
input n_172;
input n_206;
input n_217;
input n_726;
input n_982;
input n_1573;
input n_1453;
input n_1731;
input n_818;
input n_861;
input n_1713;
input n_1183;
input n_1658;
input n_899;
input n_1253;
input n_210;
input n_1737;
input n_774;
input n_1628;
input n_1335;
input n_1514;
input n_1777;
input n_1059;
input n_1345;
input n_176;
input n_1133;
input n_1771;
input n_557;
input n_1410;
input n_1005;
input n_607;
input n_1003;
input n_679;
input n_710;
input n_527;
input n_1168;
input n_707;
input n_937;
input n_1427;
input n_393;
input n_108;
input n_487;
input n_1584;
input n_665;
input n_1726;
input n_66;
input n_1440;
input n_177;
input n_421;
input n_1356;
input n_1787;
input n_910;
input n_1657;
input n_768;
input n_1475;
input n_1302;
input n_1774;
input n_1725;
input n_205;
input n_1136;
input n_1313;
input n_1491;
input n_754;
input n_1496;
input n_179;
input n_1125;
input n_125;
input n_410;
input n_708;
input n_529;
input n_735;
input n_232;
input n_1109;
input n_126;
input n_895;
input n_1310;
input n_202;
input n_427;
input n_1399;
input n_1543;
input n_791;
input n_732;
input n_1533;
input n_193;
input n_808;
input n_797;
input n_1025;
input n_500;
input n_1067;
input n_1720;
input n_148;
input n_435;
input n_159;
input n_766;
input n_1457;
input n_541;
input n_538;
input n_1117;
input n_799;
input n_687;
input n_715;
input n_1742;
input n_1480;
input n_1482;
input n_1213;
input n_1266;
input n_536;
input n_872;
input n_594;
input n_200;
input n_1291;
input n_1297;
input n_1753;
input n_1782;
input n_1155;
input n_1418;
input n_89;
input n_1524;
input n_1689;
input n_1485;
input n_115;
input n_1011;
input n_1184;
input n_985;
input n_869;
input n_810;
input n_416;
input n_827;
input n_401;
input n_1703;
input n_1352;
input n_626;
input n_1650;
input n_1144;
input n_1137;
input n_1570;
input n_1170;
input n_305;
input n_137;
input n_676;
input n_294;
input n_318;
input n_653;
input n_642;
input n_1602;
input n_194;
input n_855;
input n_1178;
input n_1461;
input n_850;
input n_684;
input n_124;
input n_268;
input n_664;
input n_503;
input n_235;
input n_1372;
input n_605;
input n_1273;
input n_353;
input n_620;
input n_643;
input n_916;
input n_1081;
input n_493;
input n_1235;
input n_703;
input n_698;
input n_980;
input n_1115;
input n_1282;
input n_1318;
input n_1783;
input n_780;
input n_998;
input n_1454;
input n_467;
input n_1227;
input n_1531;
input n_840;
input n_1334;
input n_501;
input n_823;
input n_245;
input n_725;
input n_1388;
input n_1417;
input n_1295;
input n_672;
input n_581;
input n_382;
input n_554;
input n_1625;
input n_898;
input n_1762;
input n_1013;
input n_1452;
input n_718;
input n_265;
input n_1120;
input n_719;
input n_443;
input n_1791;
input n_198;
input n_1747;
input n_714;
input n_1683;
input n_909;
input n_1497;
input n_1530;
input n_997;
input n_932;
input n_612;
input n_1409;
input n_788;
input n_1326;
input n_119;
input n_1268;
input n_559;
input n_825;
input n_508;
input n_506;
input n_1320;
input n_1663;
input n_737;
input n_1718;
input n_986;
input n_509;
input n_1317;
input n_147;
input n_1518;
input n_1715;
input n_1281;
input n_67;
input n_1192;
input n_1024;
input n_1063;
input n_209;
input n_1792;
input n_1564;
input n_1613;
input n_733;
input n_1489;
input n_1376;
input n_941;
input n_981;
input n_1569;
input n_68;
input n_867;
input n_186;
input n_134;
input n_587;
input n_63;
input n_792;
input n_756;
input n_1429;
input n_399;
input n_1238;
input n_548;
input n_812;
input n_298;
input n_518;
input n_505;
input n_1772;
input n_282;
input n_752;
input n_905;
input n_1476;
input n_1108;
input n_782;
input n_1100;
input n_1395;
input n_862;
input n_1425;
input n_760;
input n_1620;
input n_381;
input n_220;
input n_390;
input n_1330;
input n_31;
input n_481;
input n_1675;
input n_1727;
input n_1554;
input n_1745;
input n_769;
input n_42;
input n_1046;
input n_271;
input n_934;
input n_1618;
input n_826;
input n_886;
input n_1221;
input n_654;
input n_1172;
input n_167;
input n_379;
input n_428;
input n_1341;
input n_570;
input n_1641;
input n_1361;
input n_1707;
input n_853;
input n_377;
input n_751;
input n_786;
input n_1083;
input n_1142;
input n_1129;
input n_392;
input n_158;
input n_704;
input n_787;
input n_1770;
input n_138;
input n_961;
input n_1756;
input n_771;
input n_276;
input n_95;
input n_1716;
input n_1225;
input n_1520;
input n_169;
input n_522;
input n_1287;
input n_1262;
input n_400;
input n_930;
input n_181;
input n_1411;
input n_221;
input n_622;
input n_1577;
input n_1087;
input n_386;
input n_994;
input n_1701;
input n_848;
input n_1550;
input n_1498;
input n_1223;
input n_1272;
input n_104;
input n_682;
input n_1567;
input n_56;
input n_141;
input n_1247;
input n_922;
input n_816;
input n_1648;
input n_591;
input n_145;
input n_1536;
input n_1344;
input n_313;
input n_631;
input n_479;
input n_1246;
input n_1339;
input n_1478;
input n_432;
input n_1769;
input n_839;
input n_1210;
input n_1364;
input n_328;
input n_140;
input n_1250;
input n_369;
input n_871;
input n_598;
input n_685;
input n_928;
input n_608;
input n_1367;
input n_78;
input n_1460;
input n_772;
input n_1555;
input n_499;
input n_1589;
input n_517;
input n_98;
input n_402;
input n_413;
input n_1086;
input n_796;
input n_1619;
input n_236;
input n_1502;
input n_1469;
input n_1012;
input n_1;
input n_1396;
input n_1348;
input n_903;
input n_1525;
input n_1752;
input n_740;
input n_203;
input n_384;
input n_1404;
input n_80;
input n_1794;
input n_35;
input n_1315;
input n_277;
input n_1061;
input n_92;
input n_333;
input n_1298;
input n_1652;
input n_462;
input n_1193;
input n_1676;
input n_1255;
input n_258;
input n_1113;
input n_29;
input n_79;
input n_1226;
input n_722;
input n_1277;
input n_188;
input n_844;
input n_201;
input n_471;
input n_852;
input n_1487;
input n_40;
input n_1028;
input n_1601;
input n_781;
input n_474;
input n_542;
input n_463;
input n_1546;
input n_595;
input n_502;
input n_466;
input n_420;
input n_1337;
input n_1495;
input n_632;
input n_699;
input n_979;
input n_1515;
input n_1627;
input n_1245;
input n_846;
input n_1673;
input n_465;
input n_76;
input n_362;
input n_1321;
input n_170;
input n_27;
input n_161;
input n_273;
input n_585;
input n_1739;
input n_270;
input n_616;
input n_81;
input n_745;
input n_1654;
input n_1103;
input n_648;
input n_1379;
input n_312;
input n_1076;
input n_1091;
input n_1408;
input n_494;
input n_1761;
input n_641;
input n_730;
input n_1325;
input n_1595;
input n_354;
input n_575;
input n_480;
input n_425;
input n_795;
input n_695;
input n_180;
input n_656;
input n_1606;
input n_1220;
input n_37;
input n_1694;
input n_1540;
input n_229;
input n_437;
input n_1642;
input n_60;
input n_403;
input n_453;
input n_1130;
input n_720;
input n_0;
input n_1526;
input n_863;
input n_805;
input n_1604;
input n_1275;
input n_1764;
input n_113;
input n_712;
input n_246;
input n_1583;
input n_1042;
input n_1402;
input n_269;
input n_285;
input n_412;
input n_1493;
input n_657;
input n_644;
input n_1741;
input n_1160;
input n_1397;
input n_491;
input n_1258;
input n_1074;
input n_1621;
input n_251;
input n_160;
input n_566;
input n_565;
input n_1448;
input n_1507;
input n_1398;
input n_597;
input n_1181;
input n_1505;
input n_1634;
input n_1196;
input n_651;
input n_1340;
input n_334;
input n_811;
input n_1558;
input n_807;
input n_835;
input n_175;
input n_666;
input n_262;
input n_1433;
input n_1704;
input n_99;
input n_1254;
input n_1026;
input n_1234;
input n_319;
input n_364;
input n_1138;
input n_927;
input n_20;
input n_1089;
input n_1004;
input n_1186;
input n_1032;
input n_242;
input n_1681;
input n_1018;
input n_1693;
input n_438;
input n_713;
input n_904;
input n_1588;
input n_1622;
input n_166;
input n_1180;
input n_1271;
input n_533;
input n_1542;
input n_1251;
input n_278;

output n_6187;

wire n_6122;
wire n_2253;
wire n_2756;
wire n_2417;
wire n_4706;
wire n_5567;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_5287;
wire n_2327;
wire n_2899;
wire n_5484;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_5978;
wire n_2395;
wire n_5161;
wire n_5776;
wire n_5512;
wire n_5207;
wire n_2347;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_5035;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_3615;
wire n_2059;
wire n_2487;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_6072;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_4211;
wire n_3448;
wire n_3019;
wire n_2096;
wire n_3776;
wire n_2530;
wire n_4517;
wire n_2483;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1860;
wire n_4615;
wire n_2076;
wire n_6090;
wire n_5480;
wire n_2147;
wire n_3010;
wire n_2770;
wire n_4131;
wire n_5402;
wire n_2584;
wire n_5851;
wire n_3188;
wire n_5509;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_3283;
wire n_5469;
wire n_2323;
wire n_5744;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_5453;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_5202;
wire n_5648;
wire n_3214;
wire n_2091;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_5922;
wire n_4678;
wire n_2032;
wire n_2587;
wire n_5848;
wire n_5406;
wire n_6085;
wire n_3947;
wire n_3490;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_2384;
wire n_3156;
wire n_3376;
wire n_5037;
wire n_4468;
wire n_5661;
wire n_3653;
wire n_5562;
wire n_3702;
wire n_4976;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_5398;
wire n_6096;
wire n_2276;
wire n_5852;
wire n_2089;
wire n_3420;
wire n_5144;
wire n_3361;
wire n_4758;
wire n_4255;
wire n_5577;
wire n_4484;
wire n_3668;
wire n_4237;
wire n_2934;
wire n_1880;
wire n_3550;
wire n_5689;
wire n_5894;
wire n_2079;
wire n_2238;
wire n_3418;
wire n_4901;
wire n_2859;
wire n_3395;
wire n_4917;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_5825;
wire n_2968;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_4421;
wire n_6098;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_4469;
wire n_4414;
wire n_5184;
wire n_4532;
wire n_3339;
wire n_3735;
wire n_3349;
wire n_2248;
wire n_3007;
wire n_5686;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_5463;
wire n_2100;
wire n_5236;
wire n_3310;
wire n_3487;
wire n_6062;
wire n_2258;
wire n_3983;
wire n_4405;
wire n_5433;
wire n_1926;
wire n_4195;
wire n_4969;
wire n_4504;
wire n_5909;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_6043;
wire n_2987;
wire n_4567;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_2175;
wire n_5055;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_5397;
wire n_4471;
wire n_5031;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_5709;
wire n_3208;
wire n_6021;
wire n_3331;
wire n_2379;
wire n_4983;
wire n_5695;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_5860;
wire n_3649;
wire n_4302;
wire n_2514;
wire n_5862;
wire n_5189;
wire n_5381;
wire n_4786;
wire n_3257;
wire n_4160;
wire n_2293;
wire n_5854;
wire n_5516;
wire n_4051;
wire n_2028;
wire n_3009;
wire n_3981;
wire n_5936;
wire n_6126;
wire n_1841;
wire n_6027;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_1891;
wire n_5254;
wire n_3526;
wire n_2546;
wire n_3790;
wire n_3491;
wire n_4613;
wire n_4649;
wire n_1888;
wire n_5615;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_5902;
wire n_4028;
wire n_5479;
wire n_3819;
wire n_6013;
wire n_2449;
wire n_5083;
wire n_5888;
wire n_2297;
wire n_4186;
wire n_4731;
wire n_2177;
wire n_3747;
wire n_5698;
wire n_5592;
wire n_2227;
wire n_4618;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_2876;
wire n_4099;
wire n_3484;
wire n_3620;
wire n_2479;
wire n_5870;
wire n_4295;
wire n_5303;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_5807;
wire n_5863;
wire n_5943;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_4697;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_4810;
wire n_3317;
wire n_4391;
wire n_5954;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_4638;
wire n_3455;
wire n_6097;
wire n_5047;
wire n_3452;
wire n_5346;
wire n_1994;
wire n_5517;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_2796;
wire n_2342;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_6008;
wire n_3095;
wire n_2805;
wire n_5624;
wire n_4918;
wire n_5714;
wire n_5806;
wire n_3856;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_6185;
wire n_5010;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_2857;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_6004;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_2947;
wire n_5580;
wire n_4299;
wire n_5937;
wire n_4801;
wire n_3515;
wire n_2886;
wire n_2093;
wire n_2473;
wire n_3287;
wire n_3378;
wire n_5435;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_5373;
wire n_5745;
wire n_4294;
wire n_5279;
wire n_4125;
wire n_4232;
wire n_4949;
wire n_2941;
wire n_2457;
wire n_5493;
wire n_4790;
wire n_2536;
wire n_2952;
wire n_4847;
wire n_6179;
wire n_5321;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_6019;
wire n_3505;
wire n_4610;
wire n_3730;
wire n_4489;
wire n_5210;
wire n_4967;
wire n_5657;
wire n_6083;
wire n_4992;
wire n_3001;
wire n_3945;
wire n_4542;
wire n_2729;
wire n_2261;
wire n_3597;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_5857;
wire n_4534;
wire n_4500;
wire n_5014;
wire n_3185;
wire n_6087;
wire n_3523;
wire n_2829;
wire n_4597;
wire n_4329;
wire n_4087;
wire n_3811;
wire n_3200;
wire n_5756;
wire n_2231;
wire n_6041;
wire n_2017;
wire n_2604;
wire n_4257;
wire n_3453;
wire n_2390;
wire n_5708;
wire n_3213;
wire n_3077;
wire n_3474;
wire n_3984;
wire n_5927;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_1823;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_5638;
wire n_4189;
wire n_5670;
wire n_1875;
wire n_2803;
wire n_3707;
wire n_1846;
wire n_5584;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_5965;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_4687;
wire n_5751;
wire n_5664;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_5641;
wire n_4037;
wire n_2922;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2727;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_3618;
wire n_2593;
wire n_5262;
wire n_3683;
wire n_6037;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_5963;
wire n_5980;
wire n_4763;
wire n_3590;
wire n_5310;
wire n_4594;
wire n_6153;
wire n_3424;
wire n_5970;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_3171;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_5441;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_5690;
wire n_2163;
wire n_5885;
wire n_2254;
wire n_3546;
wire n_2647;
wire n_4443;
wire n_5461;
wire n_4507;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_3244;
wire n_6028;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_5629;
wire n_4452;
wire n_4348;
wire n_5634;
wire n_5430;
wire n_5362;
wire n_4355;
wire n_3494;
wire n_5702;
wire n_5050;
wire n_5063;
wire n_5229;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_3110;
wire n_4572;
wire n_3073;
wire n_5527;
wire n_5609;
wire n_5416;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_5266;
wire n_3178;
wire n_5355;
wire n_2334;
wire n_4521;
wire n_4488;
wire n_5977;
wire n_2289;
wire n_3051;
wire n_2783;
wire n_2263;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_4519;
wire n_5551;
wire n_3715;
wire n_6073;
wire n_5767;
wire n_3040;
wire n_1938;
wire n_5640;
wire n_2499;
wire n_3568;
wire n_5655;
wire n_5475;
wire n_3737;
wire n_6138;
wire n_1967;
wire n_3255;
wire n_5692;
wire n_4856;
wire n_2997;
wire n_5921;
wire n_4400;
wire n_5168;
wire n_3326;
wire n_3734;
wire n_4778;
wire n_2429;
wire n_6159;
wire n_5322;
wire n_4352;
wire n_4441;
wire n_4761;
wire n_6173;
wire n_1804;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_2364;
wire n_2533;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_5371;
wire n_2291;
wire n_4043;
wire n_3601;
wire n_5418;
wire n_1865;
wire n_2973;
wire n_2094;
wire n_2393;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_2043;
wire n_2751;
wire n_6131;
wire n_4893;
wire n_5032;
wire n_1934;
wire n_5933;
wire n_4948;
wire n_4000;
wire n_3240;
wire n_2025;
wire n_4406;
wire n_2758;
wire n_1807;
wire n_2618;
wire n_5112;
wire n_5386;
wire n_2559;
wire n_4748;
wire n_2295;
wire n_3931;
wire n_4010;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_2795;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_3380;
wire n_5644;
wire n_2098;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_5424;
wire n_3198;
wire n_2641;
wire n_1895;
wire n_4728;
wire n_4247;
wire n_4933;
wire n_4018;
wire n_3900;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_3872;
wire n_4336;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_3877;
wire n_2995;
wire n_5496;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_4052;
wire n_5864;
wire n_3459;
wire n_4398;
wire n_3155;
wire n_2633;
wire n_4954;
wire n_2435;
wire n_2097;
wire n_5460;
wire n_4304;
wire n_3911;
wire n_5333;
wire n_4431;
wire n_4192;
wire n_5570;
wire n_3736;
wire n_4805;
wire n_4885;
wire n_5983;
wire n_5804;
wire n_3565;
wire n_6167;
wire n_4701;
wire n_2575;
wire n_5910;
wire n_5040;
wire n_1904;
wire n_1899;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_4631;
wire n_3035;
wire n_5194;
wire n_5717;
wire n_5464;
wire n_5886;
wire n_3639;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_1915;
wire n_5610;
wire n_5239;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_1979;
wire n_2924;
wire n_4111;
wire n_2484;
wire n_5785;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_5305;
wire n_5994;
wire n_4538;
wire n_6093;
wire n_6010;
wire n_2754;
wire n_5376;
wire n_2489;
wire n_5204;
wire n_2012;
wire n_4094;
wire n_3503;
wire n_2866;
wire n_3561;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_4878;
wire n_3934;
wire n_4985;
wire n_5788;
wire n_3922;
wire n_3846;
wire n_5897;
wire n_2103;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_3074;
wire n_1999;
wire n_2372;
wire n_3673;
wire n_3768;
wire n_2861;
wire n_2630;
wire n_3943;
wire n_2430;
wire n_2433;
wire n_3293;
wire n_5795;
wire n_5508;
wire n_5582;
wire n_4022;
wire n_4852;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_3415;
wire n_2284;
wire n_5746;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_4601;
wire n_2687;
wire n_1890;
wire n_4220;
wire n_1944;
wire n_5630;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_5504;
wire n_4223;
wire n_1889;
wire n_5025;
wire n_2966;
wire n_2326;
wire n_2188;
wire n_6032;
wire n_4644;
wire n_4456;
wire n_5060;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_5775;
wire n_2748;
wire n_3311;
wire n_3272;
wire n_2898;
wire n_2717;
wire n_1861;
wire n_5731;
wire n_5581;
wire n_3628;
wire n_3691;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_5831;
wire n_2573;
wire n_4435;
wire n_2939;
wire n_6039;
wire n_3807;
wire n_5884;
wire n_2447;
wire n_4764;
wire n_5653;
wire n_5394;
wire n_2774;
wire n_4655;
wire n_3161;
wire n_4581;
wire n_6084;
wire n_4827;
wire n_2488;
wire n_3477;
wire n_5421;
wire n_2476;
wire n_4399;
wire n_2781;
wire n_5309;
wire n_2778;
wire n_4782;
wire n_4363;
wire n_2887;
wire n_4864;
wire n_2691;
wire n_3054;
wire n_4335;
wire n_5889;
wire n_2526;
wire n_2703;
wire n_2167;
wire n_5764;
wire n_5428;
wire n_3391;
wire n_6102;
wire n_4259;
wire n_5541;
wire n_2709;
wire n_5543;
wire n_5678;
wire n_5935;
wire n_4865;
wire n_4056;
wire n_4564;
wire n_3840;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_5950;
wire n_2173;
wire n_1842;
wire n_3738;
wire n_5995;
wire n_6162;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_6006;
wire n_3245;
wire n_4417;
wire n_6109;
wire n_4899;
wire n_2119;
wire n_2157;
wire n_2552;
wire n_5411;
wire n_2453;
wire n_4798;
wire n_3509;
wire n_3352;
wire n_5671;
wire n_3076;
wire n_3535;
wire n_2182;
wire n_3251;
wire n_2931;
wire n_5185;
wire n_3118;
wire n_3511;
wire n_3443;
wire n_2146;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_3521;
wire n_5379;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_2918;
wire n_3232;
wire n_5945;
wire n_2112;
wire n_2958;
wire n_4981;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_5811;
wire n_4430;
wire n_5565;
wire n_4081;
wire n_3132;
wire n_4407;
wire n_3951;
wire n_4894;
wire n_5780;
wire n_5643;
wire n_3238;
wire n_3210;
wire n_5846;
wire n_2036;
wire n_3267;
wire n_4995;
wire n_5524;
wire n_3964;
wire n_3772;
wire n_1956;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_6104;
wire n_3884;
wire n_3726;
wire n_2525;
wire n_2892;
wire n_2907;
wire n_6145;
wire n_3577;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_4057;
wire n_4332;
wire n_4314;
wire n_3347;
wire n_3216;
wire n_3809;
wire n_2113;
wire n_4288;
wire n_6076;
wire n_3567;
wire n_5066;
wire n_3939;
wire n_6092;
wire n_5401;
wire n_5843;
wire n_4241;
wire n_3321;
wire n_3212;
wire n_2256;
wire n_3152;
wire n_5106;
wire n_5468;
wire n_2920;
wire n_4265;
wire n_5883;
wire n_5319;
wire n_2247;
wire n_3705;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_5455;
wire n_2268;
wire n_3778;
wire n_5706;
wire n_5337;
wire n_3304;
wire n_3912;
wire n_2739;
wire n_2771;
wire n_4604;
wire n_5223;
wire n_5962;
wire n_3795;
wire n_5020;
wire n_4419;
wire n_4477;
wire n_3179;
wire n_3256;
wire n_2386;
wire n_3086;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_2568;
wire n_5364;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_5895;
wire n_4639;
wire n_3713;
wire n_3663;
wire n_5649;
wire n_5046;
wire n_5166;
wire n_3246;
wire n_2495;
wire n_5088;
wire n_2302;
wire n_5457;
wire n_5532;
wire n_2069;
wire n_3434;
wire n_1806;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_4243;
wire n_4982;
wire n_3695;
wire n_4330;
wire n_2482;
wire n_2677;
wire n_5544;
wire n_3832;
wire n_3987;
wire n_5987;
wire n_6180;
wire n_5352;
wire n_5824;
wire n_4991;
wire n_5538;
wire n_5919;
wire n_2329;
wire n_2142;
wire n_6176;
wire n_5410;
wire n_3332;
wire n_3048;
wire n_3937;
wire n_6124;
wire n_2203;
wire n_4525;
wire n_3782;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_3786;
wire n_2888;
wire n_5742;
wire n_3638;
wire n_5992;
wire n_5503;
wire n_4177;
wire n_3763;
wire n_2669;
wire n_2306;
wire n_5958;
wire n_3022;
wire n_4264;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_5129;
wire n_2149;
wire n_5500;
wire n_3060;
wire n_4276;
wire n_5219;
wire n_5605;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_5654;
wire n_2408;
wire n_5320;
wire n_1877;
wire n_3049;
wire n_5107;
wire n_5999;
wire n_4485;
wire n_4626;
wire n_6100;
wire n_2659;
wire n_4975;
wire n_1852;
wire n_5602;
wire n_3089;
wire n_6050;
wire n_2470;
wire n_5405;
wire n_3985;
wire n_5253;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_2551;
wire n_2682;
wire n_5903;
wire n_3440;
wire n_6171;
wire n_4569;
wire n_2699;
wire n_4897;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_5491;
wire n_2615;
wire n_3940;
wire n_5842;
wire n_2985;
wire n_5722;
wire n_5636;
wire n_5065;
wire n_2753;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_5492;
wire n_3141;
wire n_5084;
wire n_5667;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_4919;
wire n_4025;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_5918;
wire n_4503;
wire n_3507;
wire n_3821;
wire n_2700;
wire n_3367;
wire n_4464;
wire n_5877;
wire n_3096;
wire n_3496;
wire n_4114;
wire n_2544;
wire n_2356;
wire n_4556;
wire n_5454;
wire n_2620;
wire n_4089;
wire n_6156;
wire n_5913;
wire n_5621;
wire n_2919;
wire n_4327;
wire n_4218;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_2757;
wire n_5573;
wire n_4353;
wire n_2042;
wire n_2921;
wire n_2720;
wire n_1854;
wire n_4990;
wire n_6088;
wire n_5529;
wire n_1856;
wire n_4959;
wire n_4161;
wire n_5800;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_4466;
wire n_2262;
wire n_2462;
wire n_3625;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2837;
wire n_4844;
wire n_2979;
wire n_5257;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_2548;
wire n_5645;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_5779;
wire n_4388;
wire n_4206;
wire n_6140;
wire n_4738;
wire n_3909;
wire n_6164;
wire n_3207;
wire n_3944;
wire n_4434;
wire n_4837;
wire n_3042;
wire n_1942;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_5012;
wire n_1876;
wire n_4620;
wire n_5697;
wire n_1810;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_2222;
wire n_3510;
wire n_6147;
wire n_3218;
wire n_2667;
wire n_6011;
wire n_3150;
wire n_4325;
wire n_2413;
wire n_3775;
wire n_4133;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_4481;
wire n_3416;
wire n_4379;
wire n_2181;
wire n_1829;
wire n_6183;
wire n_5882;
wire n_4030;
wire n_4490;
wire n_3138;
wire n_4397;
wire n_2928;
wire n_4820;
wire n_3770;
wire n_5094;
wire n_4938;
wire n_4179;
wire n_3469;
wire n_5336;
wire n_2723;
wire n_5672;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_5548;
wire n_5601;
wire n_3855;
wire n_2054;
wire n_5339;
wire n_4931;
wire n_6099;
wire n_3158;
wire n_5693;
wire n_2623;
wire n_3113;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_3288;
wire n_5514;
wire n_4404;
wire n_5091;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_5486;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_5599;
wire n_6116;
wire n_4356;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_4291;
wire n_5403;
wire n_4386;
wire n_4149;
wire n_2982;
wire n_2481;
wire n_3545;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_2339;
wire n_5782;
wire n_4637;
wire n_4935;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_5608;
wire n_3741;
wire n_3410;
wire n_2029;
wire n_5298;
wire n_5596;
wire n_1887;
wire n_4413;
wire n_5728;
wire n_2346;
wire n_3990;
wire n_4493;
wire n_3475;
wire n_2882;
wire n_2338;
wire n_5726;
wire n_3672;
wire n_5290;
wire n_3197;
wire n_3109;
wire n_2721;
wire n_5095;
wire n_3002;
wire n_5324;
wire n_3897;
wire n_5928;
wire n_3845;
wire n_2081;
wire n_4570;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_5911;
wire n_2418;
wire n_5589;
wire n_5841;
wire n_2179;
wire n_2521;
wire n_3458;
wire n_5712;
wire n_3330;
wire n_4606;
wire n_6166;
wire n_4774;
wire n_2477;
wire n_3887;
wire n_4093;
wire n_4672;
wire n_3519;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_4766;
wire n_5633;
wire n_2896;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_5583;
wire n_4460;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_6064;
wire n_6110;
wire n_2255;
wire n_2272;
wire n_1965;
wire n_1902;
wire n_1941;
wire n_5501;
wire n_3938;
wire n_5377;
wire n_2878;
wire n_5652;
wire n_6135;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_3189;
wire n_2066;
wire n_3154;
wire n_6141;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_2220;
wire n_4349;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1935;
wire n_6036;
wire n_3366;
wire n_2696;
wire n_4863;
wire n_3242;
wire n_6071;
wire n_3525;
wire n_3486;
wire n_2405;
wire n_3995;
wire n_2953;
wire n_2088;
wire n_4036;
wire n_5100;
wire n_5849;
wire n_2578;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_5367;
wire n_2656;
wire n_3524;
wire n_5616;
wire n_5034;
wire n_5988;
wire n_6035;
wire n_3549;
wire n_2092;
wire n_5959;
wire n_2075;
wire n_3658;
wire n_4807;
wire n_6150;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1919;
wire n_4230;
wire n_3419;
wire n_2053;
wire n_1958;
wire n_5917;
wire n_5754;
wire n_6016;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_5628;
wire n_1808;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_5003;
wire n_5252;
wire n_2731;
wire n_6143;
wire n_5614;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_3979;
wire n_4582;
wire n_2998;
wire n_4684;
wire n_5981;
wire n_6095;
wire n_4840;
wire n_3162;
wire n_2760;
wire n_3377;
wire n_3749;
wire n_5720;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_5325;
wire n_5696;
wire n_2637;
wire n_5375;
wire n_4384;
wire n_4423;
wire n_4096;
wire n_2881;
wire n_3282;
wire n_3231;
wire n_1966;
wire n_4996;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_5759;
wire n_4478;
wire n_5753;
wire n_2646;
wire n_5536;
wire n_5173;
wire n_3920;
wire n_4890;
wire n_5691;
wire n_5794;
wire n_5027;
wire n_5647;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_4106;
wire n_3717;
wire n_5738;
wire n_2743;
wire n_2675;
wire n_3052;
wire n_5215;
wire n_3743;
wire n_1932;
wire n_4721;
wire n_5597;
wire n_5635;
wire n_1983;
wire n_5975;
wire n_4029;
wire n_3870;
wire n_4496;
wire n_3529;
wire n_1977;
wire n_2153;
wire n_4338;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_2318;
wire n_2502;
wire n_2504;
wire n_4495;
wire n_4762;
wire n_5942;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_5940;
wire n_5121;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_5555;
wire n_2446;
wire n_3488;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_5784;
wire n_5576;
wire n_4668;
wire n_4953;
wire n_5466;
wire n_3898;
wire n_5284;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_4759;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_3552;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_5578;
wire n_2361;
wire n_4113;
wire n_1998;
wire n_4686;
wire n_5530;
wire n_3759;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_5741;
wire n_5991;
wire n_3933;
wire n_3206;
wire n_5506;
wire n_3966;
wire n_5243;
wire n_5449;
wire n_5221;
wire n_4183;
wire n_4068;
wire n_4872;
wire n_6000;
wire n_4233;
wire n_3192;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_2649;
wire n_5792;
wire n_1929;
wire n_5575;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_3324;
wire n_3914;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_3742;
wire n_2252;
wire n_6113;
wire n_4819;
wire n_2576;
wire n_4900;
wire n_3390;
wire n_3746;
wire n_2373;
wire n_3817;
wire n_2745;
wire n_2493;
wire n_4930;
wire n_5276;
wire n_5078;
wire n_4537;
wire n_2885;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_4282;
wire n_3485;
wire n_4180;
wire n_3839;
wire n_5205;
wire n_3333;
wire n_5651;
wire n_2845;
wire n_6144;
wire n_4143;
wire n_4659;
wire n_2602;
wire n_5819;
wire n_4579;
wire n_4616;
wire n_3014;
wire n_2547;
wire n_5998;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_5721;
wire n_5673;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_3135;
wire n_2401;
wire n_5476;
wire n_2003;
wire n_5856;
wire n_5446;
wire n_4895;
wire n_3573;
wire n_3148;
wire n_5944;
wire n_2264;
wire n_3534;
wire n_4275;
wire n_3970;
wire n_3438;
wire n_4098;
wire n_5684;
wire n_5861;
wire n_5976;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_2184;
wire n_5312;
wire n_5850;
wire n_3217;
wire n_3425;
wire n_3404;
wire n_5111;
wire n_5890;
wire n_4055;
wire n_2926;
wire n_3540;
wire n_3670;
wire n_3973;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_5687;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_2065;
wire n_4017;
wire n_5839;
wire n_3397;
wire n_3740;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_2977;
wire n_6182;
wire n_3723;
wire n_5674;
wire n_3600;
wire n_4134;
wire n_6053;
wire n_2836;
wire n_5682;
wire n_2130;
wire n_5167;
wire n_3239;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_5612;
wire n_6125;
wire n_2850;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_4740;
wire n_5301;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_5898;
wire n_2221;
wire n_3576;
wire n_1868;
wire n_4049;
wire n_5214;
wire n_3862;
wire n_5487;
wire n_5563;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_5497;
wire n_4724;
wire n_5832;
wire n_5526;
wire n_2818;
wire n_3646;
wire n_2129;
wire n_3345;
wire n_4546;
wire n_3584;
wire n_3756;
wire n_2889;
wire n_5593;
wire n_5021;
wire n_2772;
wire n_5444;
wire n_1924;
wire n_4382;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_2260;
wire n_5389;
wire n_1813;
wire n_4833;
wire n_3056;
wire n_2345;
wire n_5110;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_5425;
wire n_3289;
wire n_1973;
wire n_5737;
wire n_2579;
wire n_4228;
wire n_4401;
wire n_6112;
wire n_2788;
wire n_2984;
wire n_3364;
wire n_5560;
wire n_1873;
wire n_3201;
wire n_5666;
wire n_3472;
wire n_6151;
wire n_2874;
wire n_5179;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_4968;
wire n_5030;
wire n_3949;
wire n_5961;
wire n_3543;
wire n_3050;
wire n_3903;
wire n_4834;
wire n_5272;
wire n_2742;
wire n_3314;
wire n_2183;
wire n_4158;
wire n_2360;
wire n_6015;
wire n_3254;
wire n_5361;
wire n_5683;
wire n_4171;
wire n_5847;
wire n_4045;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_5740;
wire n_2834;
wire n_2531;
wire n_5015;
wire n_2702;
wire n_5729;
wire n_2030;
wire n_3115;
wire n_4749;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_2234;
wire n_4804;
wire n_5545;
wire n_2209;
wire n_4270;
wire n_2797;
wire n_5152;
wire n_2321;
wire n_3680;
wire n_5905;
wire n_3497;
wire n_5409;
wire n_2940;
wire n_5688;
wire n_2612;
wire n_5128;
wire n_4566;
wire n_2841;
wire n_3322;
wire n_4576;
wire n_2505;
wire n_2427;
wire n_4061;
wire n_2070;
wire n_3250;
wire n_2594;
wire n_5798;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_5986;
wire n_3112;
wire n_2349;
wire n_3874;
wire n_5415;
wire n_4676;
wire n_5770;
wire n_5892;
wire n_4544;
wire n_2170;
wire n_5676;
wire n_5802;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_4591;
wire n_3266;
wire n_4646;
wire n_5769;
wire n_6065;
wire n_4563;
wire n_4725;
wire n_2210;
wire n_4169;
wire n_5331;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_2426;
wire n_4320;
wire n_5341;
wire n_5930;
wire n_5814;
wire n_4881;
wire n_5979;
wire n_5271;
wire n_5089;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_4012;
wire n_5518;
wire n_4636;
wire n_5637;
wire n_4584;
wire n_5622;
wire n_3910;
wire n_4711;
wire n_3319;
wire n_5240;
wire n_3335;
wire n_5813;
wire n_3413;
wire n_5495;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_5546;
wire n_2689;
wire n_3259;
wire n_5482;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_3688;
wire n_3016;
wire n_5393;
wire n_2599;
wire n_3338;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_5966;
wire n_5041;
wire n_5431;
wire n_2200;
wire n_3261;
wire n_5026;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_5059;
wire n_5505;
wire n_3127;
wire n_3732;
wire n_4250;
wire n_5329;
wire n_3596;
wire n_4699;
wire n_3906;
wire n_4127;
wire n_3297;
wire n_2683;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_5908;
wire n_6018;
wire n_4202;
wire n_5212;
wire n_5000;
wire n_2853;
wire n_5939;
wire n_3766;
wire n_2880;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_5931;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_5420;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_3621;
wire n_5234;
wire n_5835;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_6029;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_5440;
wire n_5679;
wire n_3710;
wire n_5938;
wire n_4155;
wire n_2031;
wire n_3891;
wire n_5891;
wire n_4144;
wire n_5724;
wire n_5774;
wire n_2165;
wire n_3379;
wire n_4374;
wire n_3532;
wire n_5131;
wire n_1818;
wire n_2127;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_4548;
wire n_5923;
wire n_5790;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_1845;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_4816;
wire n_2983;
wire n_3810;
wire n_2715;
wire n_6132;
wire n_5598;
wire n_2085;
wire n_5306;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_2672;
wire n_2651;
wire n_4358;
wire n_5147;
wire n_3656;
wire n_2071;
wire n_2643;
wire n_2561;
wire n_4793;
wire n_5677;
wire n_4168;
wire n_3446;
wire n_5997;
wire n_5511;
wire n_5680;
wire n_3028;
wire n_4806;
wire n_4350;
wire n_5533;
wire n_5838;
wire n_6058;
wire n_5280;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_6170;
wire n_1931;
wire n_4187;
wire n_4166;
wire n_5206;
wire n_3222;
wire n_1801;
wire n_5419;
wire n_6130;
wire n_2970;
wire n_2235;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_3755;
wire n_5803;
wire n_4258;
wire n_6014;
wire n_4498;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_4064;
wire n_4936;
wire n_5387;
wire n_1863;
wire n_3841;
wire n_2118;
wire n_4770;
wire n_5985;
wire n_2944;
wire n_2407;
wire n_4907;
wire n_5058;
wire n_6158;
wire n_3262;
wire n_6119;
wire n_5018;
wire n_4006;
wire n_5896;
wire n_4861;
wire n_3690;
wire n_2358;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_2833;
wire n_4712;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_1950;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_5097;
wire n_2750;
wire n_5730;
wire n_3899;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_5816;
wire n_4069;
wire n_2784;
wire n_3718;
wire n_3092;
wire n_3470;
wire n_4862;
wire n_2557;
wire n_5300;
wire n_4850;
wire n_3781;
wire n_4813;
wire n_4912;
wire n_2590;
wire n_2330;
wire n_5748;
wire n_2942;
wire n_5525;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_3889;
wire n_6139;
wire n_4256;
wire n_4224;
wire n_3508;
wire n_4024;
wire n_2267;
wire n_2218;
wire n_5650;
wire n_2636;
wire n_1825;
wire n_1951;
wire n_5400;
wire n_1883;
wire n_2759;
wire n_4415;
wire n_5552;
wire n_4702;
wire n_4252;
wire n_4457;
wire n_6063;
wire n_5139;
wire n_2319;
wire n_3481;
wire n_5481;
wire n_2808;
wire n_6070;
wire n_2679;
wire n_2676;
wire n_5821;
wire n_4491;
wire n_2930;
wire n_5733;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_5871;
wire n_2611;
wire n_4261;
wire n_6184;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_2698;
wire n_5043;
wire n_5707;
wire n_4001;
wire n_3047;
wire n_2454;
wire n_4371;
wire n_5836;
wire n_5281;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_4268;
wire n_5048;
wire n_5521;
wire n_5028;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_4194;
wire n_5585;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_2990;
wire n_6121;
wire n_3119;
wire n_4142;
wire n_4082;
wire n_5561;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_3279;
wire n_2621;
wire n_5799;
wire n_5073;
wire n_5024;
wire n_5875;
wire n_4262;
wire n_2671;
wire n_1798;
wire n_4720;
wire n_4685;
wire n_6101;
wire n_5968;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_5812;
wire n_6148;
wire n_5515;
wire n_6106;
wire n_4014;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_2913;
wire n_2336;
wire n_5607;
wire n_4175;
wire n_2005;
wire n_1916;
wire n_4648;
wire n_5006;
wire n_5734;
wire n_6081;
wire n_4892;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_4970;
wire n_3816;
wire n_5404;
wire n_4108;
wire n_4486;
wire n_6047;
wire n_2960;
wire n_5438;
wire n_4627;
wire n_2290;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_2145;
wire n_5725;
wire n_3030;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_5163;
wire n_2039;
wire n_5768;
wire n_4961;
wire n_3753;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_3396;
wire n_4023;
wire n_4420;
wire n_5685;
wire n_1923;
wire n_5773;
wire n_6055;
wire n_5138;
wire n_5374;
wire n_6108;
wire n_2116;
wire n_6165;
wire n_1828;
wire n_2320;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_4396;
wire n_5127;
wire n_4367;
wire n_2087;
wire n_5485;
wire n_5766;
wire n_5216;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_5805;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_2355;
wire n_2133;
wire n_3830;
wire n_2585;
wire n_2725;
wire n_5175;
wire n_3883;
wire n_4152;
wire n_2565;
wire n_5948;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_5611;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_5900;
wire n_3466;
wire n_4962;
wire n_2595;
wire n_3411;
wire n_4958;
wire n_4271;
wire n_5171;
wire n_3586;
wire n_5554;
wire n_4071;
wire n_4921;
wire n_1980;
wire n_5427;
wire n_5639;
wire n_3065;
wire n_4361;
wire n_5417;
wire n_4614;
wire n_2681;
wire n_3103;
wire n_4945;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_2775;
wire n_4693;
wire n_5488;
wire n_4326;
wire n_3557;
wire n_2230;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_6127;
wire n_2851;
wire n_4305;
wire n_5781;
wire n_2490;
wire n_4213;
wire n_2849;
wire n_3692;
wire n_2204;
wire n_5747;
wire n_5969;
wire n_4929;
wire n_1961;
wire n_4964;
wire n_6079;
wire n_4802;
wire n_4139;
wire n_3029;
wire n_2508;
wire n_4031;
wire n_2416;
wire n_5437;
wire n_5826;
wire n_3881;
wire n_2461;
wire n_2243;
wire n_4583;
wire n_4210;
wire n_5245;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_2368;
wire n_2890;
wire n_2554;
wire n_3698;
wire n_3927;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_4891;
wire n_5603;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_5716;
wire n_3993;
wire n_4940;
wire n_5208;
wire n_3588;
wire n_2308;
wire n_4590;
wire n_5606;
wire n_4830;
wire n_5231;
wire n_5237;
wire n_4664;
wire n_3860;
wire n_5456;
wire n_3160;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_6040;
wire n_3847;
wire n_4946;
wire n_4906;
wire n_5727;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_5390;
wire n_5347;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_2440;
wire n_4883;
wire n_2923;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_4297;
wire n_5833;
wire n_3800;
wire n_2403;
wire n_5407;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_3991;
wire n_3134;
wire n_4172;
wire n_4791;
wire n_4536;
wire n_5149;
wire n_5967;
wire n_2463;
wire n_5151;
wire n_4773;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_2472;
wire n_4611;
wire n_4755;
wire n_5982;
wire n_2294;
wire n_4960;
wire n_2993;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2948;
wire n_2309;
wire n_5827;
wire n_5494;
wire n_4362;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2685;
wire n_2037;
wire n_1953;
wire n_4422;
wire n_6123;
wire n_2589;
wire n_3482;
wire n_6082;
wire n_2233;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_5228;
wire n_3956;
wire n_5758;
wire n_5323;
wire n_3572;
wire n_4215;
wire n_4280;
wire n_3375;
wire n_4047;
wire n_5471;
wire n_5434;
wire n_2082;
wire n_5941;
wire n_5879;
wire n_3167;
wire n_5558;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_5338;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_5669;
wire n_3854;
wire n_2468;
wire n_3078;
wire n_3253;
wire n_4027;
wire n_2280;
wire n_4599;
wire n_5830;
wire n_3363;
wire n_4812;
wire n_5760;
wire n_3689;
wire n_2020;
wire n_4628;
wire n_5668;
wire n_1881;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_5878;
wire n_5588;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_5765;
wire n_3950;
wire n_4458;
wire n_4121;
wire n_5090;
wire n_4476;
wire n_5613;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_6080;
wire n_1848;
wire n_5571;
wire n_2126;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_5513;
wire n_4803;
wire n_5972;
wire n_4079;
wire n_4091;
wire n_5916;
wire n_5984;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_6094;
wire n_2935;
wire n_5132;
wire n_5191;
wire n_3085;
wire n_5869;
wire n_5925;
wire n_5359;
wire n_2574;
wire n_5293;
wire n_4316;
wire n_3697;
wire n_2638;
wire n_4044;
wire n_4062;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_5510;
wire n_6046;
wire n_2016;
wire n_2949;
wire n_2711;
wire n_5363;
wire n_5200;
wire n_5659;
wire n_5618;
wire n_2867;
wire n_1894;
wire n_2794;
wire n_3145;
wire n_3124;
wire n_4253;
wire n_5356;
wire n_5369;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_3517;
wire n_3100;
wire n_2522;
wire n_6111;
wire n_1834;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_3506;
wire n_3605;
wire n_2409;
wire n_5858;
wire n_5817;
wire n_3402;
wire n_5723;
wire n_5295;
wire n_6137;
wire n_4679;
wire n_4115;
wire n_4998;
wire n_2988;
wire n_1970;
wire n_2766;
wire n_5627;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_2205;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_3401;
wire n_3226;
wire n_3902;
wire n_4730;
wire n_6074;
wire n_2779;
wire n_3654;
wire n_2164;
wire n_5996;
wire n_2115;
wire n_2232;
wire n_5327;
wire n_6045;
wire n_4713;
wire n_5137;
wire n_2811;
wire n_3348;
wire n_5796;
wire n_6068;
wire n_3358;
wire n_5791;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_1991;
wire n_2224;
wire n_5906;
wire n_4743;
wire n_3805;
wire n_3825;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_2692;
wire n_2008;
wire n_4654;
wire n_6157;
wire n_5423;
wire n_4733;
wire n_3792;
wire n_6017;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_2283;
wire n_3278;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_5736;
wire n_3312;
wire n_6105;
wire n_2197;
wire n_2199;
wire n_5069;
wire n_5700;
wire n_3285;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_6091;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_2480;
wire n_6034;
wire n_2363;
wire n_4072;
wire n_5579;
wire n_4781;
wire n_3606;
wire n_5004;
wire n_2550;
wire n_4424;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_5837;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_3878;
wire n_4450;
wire n_5642;
wire n_3553;
wire n_5880;
wire n_6169;
wire n_4746;
wire n_5713;
wire n_6005;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_3850;
wire n_4459;
wire n_2996;
wire n_5793;
wire n_5591;
wire n_4050;
wire n_2315;
wire n_3228;
wire n_2102;
wire n_5623;
wire n_5681;
wire n_4853;
wire n_2422;
wire n_2239;
wire n_6118;
wire n_5256;
wire n_2950;
wire n_5220;
wire n_5732;
wire n_3852;
wire n_5178;
wire n_4520;
wire n_2057;
wire n_4008;
wire n_5507;
wire n_5077;
wire n_5872;
wire n_3858;
wire n_1901;
wire n_6115;
wire n_4502;
wire n_3032;
wire n_4851;
wire n_5735;
wire n_3072;
wire n_3081;
wire n_3313;
wire n_2710;
wire n_3924;
wire n_4571;
wire n_2006;
wire n_5314;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_2535;
wire n_4205;
wire n_5953;
wire n_2726;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_5952;
wire n_4739;
wire n_5820;
wire n_2376;
wire n_5483;
wire n_3017;
wire n_5718;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_4879;
wire n_5051;
wire n_3926;
wire n_6152;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_2854;
wire n_4181;
wire n_5777;
wire n_2764;
wire n_4225;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_4153;
wire n_5156;
wire n_5926;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_4783;
wire n_2964;
wire n_3769;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_5951;
wire n_2442;
wire n_1943;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_6154;
wire n_6020;
wire n_2883;
wire n_4182;
wire n_2912;
wire n_4825;
wire n_5701;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_5120;
wire n_5470;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_5797;
wire n_4839;
wire n_5222;
wire n_5743;
wire n_4016;
wire n_5772;
wire n_3435;
wire n_3575;
wire n_5801;
wire n_6117;
wire n_4231;
wire n_3165;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_4083;
wire n_1937;
wire n_5971;
wire n_4461;
wire n_3234;
wire n_5392;
wire n_2381;
wire n_3303;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3024;
wire n_5443;
wire n_3512;
wire n_5600;
wire n_4939;
wire n_5169;
wire n_4389;
wire n_3930;
wire n_4448;
wire n_2161;
wire n_6160;
wire n_2404;
wire n_2083;
wire n_2503;
wire n_1936;
wire n_6031;
wire n_5502;
wire n_2027;
wire n_5568;
wire n_2642;
wire n_2500;
wire n_1918;
wire n_5656;
wire n_4831;
wire n_2513;
wire n_5974;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_2414;
wire n_3662;
wire n_4319;
wire n_5474;
wire n_2229;
wire n_4596;
wire n_5413;
wire n_2004;
wire n_5412;
wire n_3694;
wire n_2586;
wire n_6069;
wire n_5752;
wire n_4726;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_6030;
wire n_6077;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_5201;
wire n_4474;
wire n_5217;
wire n_5957;
wire n_2511;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_5490;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_5158;
wire n_4884;
wire n_4366;
wire n_4009;
wire n_4580;
wire n_6177;
wire n_5912;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_6033;
wire n_1859;
wire n_5557;
wire n_5472;
wire n_2955;
wire n_4112;
wire n_6002;
wire n_4337;
wire n_5711;
wire n_4138;
wire n_5396;
wire n_5335;
wire n_2520;
wire n_2134;
wire n_5960;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_5143;
wire n_4238;
wire n_6142;
wire n_2374;
wire n_5859;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_2396;
wire n_1799;
wire n_4734;
wire n_1939;
wire n_2486;
wire n_6163;
wire n_4635;
wire n_3501;
wire n_1869;
wire n_4013;
wire n_3039;
wire n_2011;
wire n_6025;
wire n_4242;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_5283;
wire n_5268;
wire n_4561;
wire n_2639;
wire n_6089;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_3186;
wire n_4955;
wire n_5556;
wire n_5462;
wire n_4501;
wire n_3696;
wire n_3650;
wire n_5840;
wire n_2761;
wire n_3157;
wire n_2537;
wire n_2144;
wire n_6049;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_6052;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_1949;
wire n_2936;
wire n_1946;
wire n_5914;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_6061;
wire n_4369;
wire n_5378;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_5542;
wire n_1831;
wire n_4394;
wire n_1850;
wire n_5519;
wire n_3101;
wire n_3669;
wire n_6009;
wire n_5278;
wire n_2663;
wire n_5586;
wire n_2693;
wire n_3798;
wire n_4065;
wire n_5187;
wire n_4944;
wire n_5675;
wire n_2249;
wire n_2180;
wire n_4135;
wire n_2632;
wire n_5771;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_6051;
wire n_4716;
wire n_4942;
wire n_5844;
wire n_2432;
wire n_3405;
wire n_4745;
wire n_6155;
wire n_2337;
wire n_3907;
wire n_5344;
wire n_4629;
wire n_2932;
wire n_2980;
wire n_5225;
wire n_3306;
wire n_5662;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1986;
wire n_4752;
wire n_5265;
wire n_3986;
wire n_4376;
wire n_5705;
wire n_4753;
wire n_4552;
wire n_3885;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_5574;
wire n_5126;
wire n_2214;
wire n_3427;
wire n_2055;
wire n_4067;
wire n_5553;
wire n_4176;
wire n_4042;
wire n_4385;
wire n_3320;
wire n_5009;
wire n_2688;
wire n_5368;
wire n_5626;
wire n_6114;
wire n_3651;
wire n_4333;
wire n_3359;
wire n_2865;
wire n_2706;
wire n_5499;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_5604;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_4815;
wire n_4246;
wire n_3580;
wire n_2139;
wire n_4609;
wire n_5291;
wire n_5876;
wire n_5114;
wire n_2674;
wire n_4088;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_4462;
wire n_4472;
wire n_3433;
wire n_5288;
wire n_2305;
wire n_5540;
wire n_5699;
wire n_2450;
wire n_3447;
wire n_5810;
wire n_3305;
wire n_4151;
wire n_4148;
wire n_3528;
wire n_4373;
wire n_5762;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_4630;
wire n_5408;
wire n_4643;
wire n_4331;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_3296;
wire n_2762;
wire n_4683;
wire n_5366;
wire n_1847;
wire n_2767;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_6146;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_5477;
wire n_5451;
wire n_3923;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_5086;
wire n_2801;
wire n_5901;
wire n_4011;
wire n_4905;
wire n_2763;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_1997;
wire n_3748;
wire n_3142;
wire n_4278;
wire n_4623;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_5053;
wire n_4553;
wire n_3978;
wire n_4809;
wire n_5226;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_5867;
wire n_6048;
wire n_2491;
wire n_5079;
wire n_5590;
wire n_3833;
wire n_5632;
wire n_4841;
wire n_2022;
wire n_3814;
wire n_2592;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_3513;
wire n_3133;
wire n_5660;
wire n_4645;
wire n_2992;
wire n_6174;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_6023;
wire n_2517;
wire n_3128;
wire n_5426;
wire n_2631;
wire n_2178;
wire n_2469;
wire n_5625;
wire n_5778;
wire n_3355;
wire n_2007;
wire n_3917;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_5531;
wire n_3000;
wire n_5429;
wire n_3108;
wire n_3111;
wire n_1839;
wire n_1837;
wire n_5818;
wire n_5646;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_2875;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_5448;
wire n_3471;
wire n_5432;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_3564;
wire n_3988;
wire n_6161;
wire n_3457;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_5445;
wire n_3630;
wire n_3271;
wire n_4771;
wire n_5719;
wire n_6128;
wire n_4086;
wire n_2412;
wire n_4814;
wire n_2084;
wire n_3648;
wire n_5749;
wire n_3075;
wire n_3173;
wire n_5332;
wire n_5108;
wire n_4692;
wire n_3031;
wire n_3701;
wire n_3243;
wire n_2666;
wire n_3385;
wire n_2171;
wire n_4708;
wire n_2768;
wire n_2314;
wire n_4826;
wire n_3343;
wire n_2420;
wire n_5489;
wire n_3767;
wire n_2873;
wire n_2299;
wire n_2540;
wire n_4589;
wire n_5057;
wire n_4578;
wire n_2162;
wire n_2847;
wire n_2051;
wire n_3221;
wire n_5436;
wire n_5907;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_6044;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_3502;
wire n_3098;
wire n_5013;
wire n_2312;
wire n_3015;
wire n_1920;
wire n_5569;
wire n_5439;
wire n_5619;
wire n_4147;
wire n_2048;
wire n_3607;
wire n_4925;
wire n_1921;
wire n_4974;
wire n_1800;
wire n_4932;
wire n_4510;
wire n_2571;
wire n_6181;
wire n_3276;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_5715;
wire n_6133;
wire n_3827;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_4285;
wire n_5887;
wire n_4651;
wire n_6038;
wire n_4818;
wire n_4514;
wire n_4800;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_2110;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_2033;
wire n_4341;
wire n_4312;
wire n_3399;
wire n_2628;
wire n_5932;
wire n_6178;
wire n_2132;
wire n_6012;
wire n_2400;
wire n_4633;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_3387;
wire n_5186;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_5828;
wire n_2831;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_4832;
wire n_4207;
wire n_4545;
wire n_3037;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_5054;
wire n_5631;
wire n_2467;
wire n_2288;
wire n_4063;
wire n_5399;
wire n_3592;
wire n_5694;
wire n_4650;
wire n_4888;
wire n_5326;
wire n_3394;
wire n_4874;
wire n_3793;
wire n_4669;
wire n_4339;
wire n_4041;
wire n_5459;
wire n_2858;
wire n_4060;
wire n_2658;
wire n_2895;
wire n_2128;
wire n_5528;
wire n_3097;
wire n_5391;
wire n_4541;
wire n_3824;
wire n_5422;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_5523;
wire n_3465;
wire n_4796;
wire n_3589;
wire n_2534;
wire n_6186;
wire n_4799;
wire n_5153;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_2789;
wire n_4775;
wire n_2216;
wire n_5044;
wire n_5809;
wire n_1897;
wire n_5365;
wire n_2933;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_2328;
wire n_4248;
wire n_5915;
wire n_5452;
wire n_4754;
wire n_4554;
wire n_5595;
wire n_4845;
wire n_3053;
wire n_3893;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_5535;
wire n_3875;
wire n_5370;
wire n_4003;
wire n_5372;
wire n_5299;
wire n_2402;
wire n_5594;
wire n_4301;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_1844;
wire n_3777;
wire n_5761;
wire n_4784;
wire n_2999;
wire n_5550;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_3537;
wire n_5209;
wire n_3080;
wire n_4199;
wire n_2701;
wire n_5929;
wire n_3362;
wire n_5559;
wire n_3105;
wire n_5478;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_6022;
wire n_4470;
wire n_2236;
wire n_2816;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_4188;
wire n_3913;
wire n_3417;
wire n_5868;
wire n_4034;
wire n_3327;
wire n_6172;
wire n_5275;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_2755;
wire n_5989;
wire n_3237;
wire n_1992;
wire n_4402;
wire n_4239;
wire n_3400;
wire n_4550;
wire n_3382;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_4201;
wire n_6168;
wire n_3316;
wire n_5242;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_3603;
wire n_4123;
wire n_2192;
wire n_5520;
wire n_3633;
wire n_4479;
wire n_2670;
wire n_5947;
wire n_4416;
wire n_3372;
wire n_4539;
wire n_2707;
wire n_5920;
wire n_2471;
wire n_6149;
wire n_3230;
wire n_5808;
wire n_3342;
wire n_6054;
wire n_4682;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_5458;
wire n_3861;
wire n_5617;
wire n_4736;
wire n_3780;
wire n_1928;
wire n_5244;
wire n_5382;
wire n_6107;
wire n_3957;
wire n_5274;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_6134;
wire n_5384;
wire n_3608;
wire n_6056;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_5587;
wire n_2619;
wire n_2444;
wire n_5789;
wire n_3123;
wire n_5787;
wire n_5056;
wire n_5249;
wire n_3393;
wire n_5198;
wire n_5360;
wire n_5233;
wire n_4887;
wire n_5829;
wire n_4617;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_5866;
wire n_4005;
wire n_4904;
wire n_5899;
wire n_4792;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_4980;
wire n_6026;
wire n_4290;
wire n_5247;
wire n_5865;
wire n_3727;
wire n_5317;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_2431;
wire n_4956;
wire n_5380;
wire n_2206;
wire n_5924;
wire n_3182;
wire n_5822;
wire n_2564;
wire n_4947;
wire n_4656;
wire n_3896;
wire n_3958;
wire n_3450;
wire n_4729;
wire n_5786;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_2000;
wire n_2074;
wire n_3174;
wire n_2217;
wire n_3398;
wire n_2307;
wire n_5658;
wire n_3408;
wire n_2722;
wire n_5388;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_3432;
wire n_3090;
wire n_2437;
wire n_3762;
wire n_5564;
wire n_2445;
wire n_1835;
wire n_1988;
wire n_6042;
wire n_1853;
wire n_6057;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_3972;
wire n_5539;
wire n_3308;
wire n_5036;
wire n_5547;
wire n_4772;
wire n_3467;
wire n_4322;
wire n_2830;
wire n_5893;
wire n_4354;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_5273;
wire n_4677;
wire n_3901;
wire n_5261;
wire n_3757;
wire n_3381;
wire n_5193;
wire n_2245;
wire n_4909;
wire n_2965;
wire n_3635;
wire n_6024;
wire n_5022;
wire n_5005;
wire n_2814;
wire n_3882;
wire n_3046;
wire n_2213;
wire n_5993;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_5703;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_5534;
wire n_3204;
wire n_2136;
wire n_5174;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_4380;
wire n_3129;
wire n_4126;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_5904;
wire n_4880;
wire n_1907;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_5620;
wire n_5061;
wire n_5750;
wire n_5572;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_2187;
wire n_3023;
wire n_5881;
wire n_5815;
wire n_4193;
wire n_5873;
wire n_4075;
wire n_3104;
wire n_4737;
wire n_3647;
wire n_5755;
wire n_2819;
wire n_5949;
wire n_5195;
wire n_3609;
wire n_4136;
wire n_1952;
wire n_4393;
wire n_3720;
wire n_4535;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_4794;
wire n_5955;
wire n_3959;
wire n_5763;
wire n_3140;
wire n_5246;
wire n_5964;
wire n_3724;
wire n_2104;
wire n_3011;
wire n_5164;
wire n_4196;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_5665;
wire n_3069;
wire n_5498;
wire n_4370;
wire n_1900;
wire n_5783;
wire n_5183;
wire n_6075;
wire n_3084;
wire n_6120;
wire n_2735;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_5549;
wire n_2411;
wire n_3761;
wire n_4889;
wire n_2014;
wire n_2986;
wire n_5442;
wire n_5739;
wire n_3184;
wire n_4828;
wire n_6003;
wire n_5385;
wire n_4558;
wire n_2172;
wire n_6066;
wire n_6086;
wire n_4722;
wire n_3626;
wire n_4768;
wire n_4100;
wire n_2250;
wire n_5845;
wire n_4092;
wire n_5990;
wire n_3908;
wire n_6175;
wire n_6060;
wire n_2423;
wire n_3671;
wire n_5663;
wire n_3344;
wire n_2194;
wire n_4465;
wire n_5973;
wire n_3302;
wire n_5537;
wire n_5304;
wire n_2680;
wire n_6059;
wire n_5130;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_6103;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_1797;
wire n_2957;
wire n_5855;
wire n_2357;
wire n_5757;
wire n_3309;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_4116;
wire n_5704;
wire n_2570;
wire n_1858;
wire n_2815;
wire n_5473;
wire n_3754;
wire n_4612;
wire n_5946;
wire n_2744;
wire n_4287;
wire n_2397;
wire n_2208;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_2591;
wire n_3384;
wire n_4602;
wire n_5172;
wire n_4449;
wire n_1864;
wire n_5710;
wire n_6067;
wire n_5070;
wire n_4445;
wire n_5566;
wire n_5414;
wire n_4870;
wire n_2438;
wire n_2832;
wire n_1975;
wire n_2296;
wire n_3181;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_6129;
wire n_2135;
wire n_5450;
wire n_3493;
wire n_5313;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_6136;
wire n_5834;
wire n_2823;
wire n_5874;
wire n_5270;
wire n_5956;
wire n_4345;
wire n_5188;
wire n_3281;
wire n_3307;
wire n_6078;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_5823;
wire n_3997;
wire n_5465;
wire n_4032;
wire n_3582;
wire n_5853;
wire n_2826;
wire n_3539;
wire n_4343;
wire n_4212;
wire n_4124;
wire n_5467;
wire n_5522;
wire n_4492;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_4364;
wire n_4245;
wire n_4928;
wire n_2225;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3853;
wire n_4216;
wire n_5934;
wire n_2019;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_3721;
wire n_2026;
wire n_2109;
wire n_2013;
wire n_1990;
wire n_2614;
wire n_2991;
wire n_6001;
wire n_6007;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_3473;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_5395;
wire n_2237;
wire n_3463;
wire n_3699;
wire n_5067;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_2728;
wire n_3857;

BUFx5_ASAP7_75t_L g1797 ( 
.A(n_1773),
.Y(n_1797)
);

CKINVDCx20_ASAP7_75t_R g1798 ( 
.A(n_1197),
.Y(n_1798)
);

INVxp67_ASAP7_75t_SL g1799 ( 
.A(n_280),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1768),
.Y(n_1800)
);

CKINVDCx16_ASAP7_75t_R g1801 ( 
.A(n_1780),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1652),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1667),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1552),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1195),
.Y(n_1805)
);

INVx1_ASAP7_75t_SL g1806 ( 
.A(n_592),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_313),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_553),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1783),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1425),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1710),
.Y(n_1811)
);

BUFx2_ASAP7_75t_L g1812 ( 
.A(n_1466),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_1620),
.Y(n_1813)
);

CKINVDCx20_ASAP7_75t_R g1814 ( 
.A(n_1681),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_248),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_97),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_785),
.Y(n_1817)
);

CKINVDCx20_ASAP7_75t_R g1818 ( 
.A(n_635),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1075),
.Y(n_1819)
);

INVx2_ASAP7_75t_SL g1820 ( 
.A(n_1608),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1389),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_281),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_427),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1337),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_L g1825 ( 
.A(n_1625),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_707),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1566),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_1621),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_197),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1075),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1451),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_409),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1609),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_835),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1604),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1527),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_693),
.Y(n_1837)
);

BUFx6f_ASAP7_75t_L g1838 ( 
.A(n_1699),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_1324),
.Y(n_1839)
);

CKINVDCx20_ASAP7_75t_R g1840 ( 
.A(n_454),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1773),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1750),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_398),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1362),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_416),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_977),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_679),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_585),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_1139),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_660),
.Y(n_1850)
);

BUFx3_ASAP7_75t_L g1851 ( 
.A(n_203),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_461),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1395),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1639),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_910),
.Y(n_1855)
);

BUFx6f_ASAP7_75t_L g1856 ( 
.A(n_1726),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_1560),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1035),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1640),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_8),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_66),
.Y(n_1861)
);

BUFx3_ASAP7_75t_L g1862 ( 
.A(n_794),
.Y(n_1862)
);

CKINVDCx20_ASAP7_75t_R g1863 ( 
.A(n_235),
.Y(n_1863)
);

INVx1_ASAP7_75t_SL g1864 ( 
.A(n_1186),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1555),
.Y(n_1865)
);

INVx1_ASAP7_75t_SL g1866 ( 
.A(n_1505),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1724),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1575),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1504),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_78),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1562),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_1101),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_427),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1613),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1573),
.Y(n_1875)
);

HB1xp67_ASAP7_75t_L g1876 ( 
.A(n_1691),
.Y(n_1876)
);

INVx2_ASAP7_75t_SL g1877 ( 
.A(n_680),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1303),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1723),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1448),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1369),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_161),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1177),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_839),
.Y(n_1884)
);

BUFx5_ASAP7_75t_L g1885 ( 
.A(n_1635),
.Y(n_1885)
);

CKINVDCx20_ASAP7_75t_R g1886 ( 
.A(n_1674),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_1549),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1271),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1614),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_452),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1754),
.Y(n_1891)
);

HB1xp67_ASAP7_75t_L g1892 ( 
.A(n_408),
.Y(n_1892)
);

CKINVDCx20_ASAP7_75t_R g1893 ( 
.A(n_1671),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1654),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1392),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1626),
.Y(n_1896)
);

BUFx2_ASAP7_75t_L g1897 ( 
.A(n_1565),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_40),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_121),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_421),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1192),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1220),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_1567),
.Y(n_1903)
);

BUFx2_ASAP7_75t_L g1904 ( 
.A(n_1256),
.Y(n_1904)
);

INVx2_ASAP7_75t_SL g1905 ( 
.A(n_186),
.Y(n_1905)
);

BUFx2_ASAP7_75t_L g1906 ( 
.A(n_1687),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1619),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1047),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_404),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_896),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_411),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_534),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_1605),
.Y(n_1913)
);

CKINVDCx16_ASAP7_75t_R g1914 ( 
.A(n_1623),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_569),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_1429),
.Y(n_1916)
);

BUFx8_ASAP7_75t_SL g1917 ( 
.A(n_884),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1789),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_1256),
.Y(n_1919)
);

BUFx6f_ASAP7_75t_L g1920 ( 
.A(n_441),
.Y(n_1920)
);

CKINVDCx20_ASAP7_75t_R g1921 ( 
.A(n_1607),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_871),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_610),
.Y(n_1923)
);

BUFx10_ASAP7_75t_L g1924 ( 
.A(n_1693),
.Y(n_1924)
);

CKINVDCx5p33_ASAP7_75t_R g1925 ( 
.A(n_563),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_930),
.Y(n_1926)
);

CKINVDCx20_ASAP7_75t_R g1927 ( 
.A(n_1708),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1704),
.Y(n_1928)
);

CKINVDCx5p33_ASAP7_75t_R g1929 ( 
.A(n_1638),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1452),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1434),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_813),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_989),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1273),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1576),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1641),
.Y(n_1936)
);

BUFx2_ASAP7_75t_SL g1937 ( 
.A(n_318),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_549),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_1483),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1720),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_769),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_741),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_96),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_135),
.Y(n_1944)
);

CKINVDCx5p33_ASAP7_75t_R g1945 ( 
.A(n_824),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1140),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1678),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1575),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_477),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_572),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1166),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_843),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_282),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1016),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_1002),
.Y(n_1955)
);

INVx2_ASAP7_75t_SL g1956 ( 
.A(n_1146),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1679),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_98),
.Y(n_1958)
);

BUFx5_ASAP7_75t_L g1959 ( 
.A(n_116),
.Y(n_1959)
);

INVx2_ASAP7_75t_SL g1960 ( 
.A(n_170),
.Y(n_1960)
);

BUFx5_ASAP7_75t_L g1961 ( 
.A(n_386),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_744),
.Y(n_1962)
);

CKINVDCx16_ASAP7_75t_R g1963 ( 
.A(n_809),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1590),
.Y(n_1964)
);

CKINVDCx20_ASAP7_75t_R g1965 ( 
.A(n_1374),
.Y(n_1965)
);

CKINVDCx5p33_ASAP7_75t_R g1966 ( 
.A(n_513),
.Y(n_1966)
);

CKINVDCx20_ASAP7_75t_R g1967 ( 
.A(n_1765),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1211),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1676),
.Y(n_1969)
);

CKINVDCx20_ASAP7_75t_R g1970 ( 
.A(n_1042),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1478),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_497),
.Y(n_1972)
);

BUFx10_ASAP7_75t_L g1973 ( 
.A(n_277),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1624),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_1785),
.Y(n_1975)
);

CKINVDCx14_ASAP7_75t_R g1976 ( 
.A(n_703),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_1467),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1710),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_990),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1228),
.Y(n_1980)
);

CKINVDCx16_ASAP7_75t_R g1981 ( 
.A(n_185),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_362),
.Y(n_1982)
);

INVx1_ASAP7_75t_SL g1983 ( 
.A(n_1627),
.Y(n_1983)
);

CKINVDCx5p33_ASAP7_75t_R g1984 ( 
.A(n_479),
.Y(n_1984)
);

INVx1_ASAP7_75t_SL g1985 ( 
.A(n_1616),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1610),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_963),
.Y(n_1987)
);

CKINVDCx5p33_ASAP7_75t_R g1988 ( 
.A(n_849),
.Y(n_1988)
);

INVx2_ASAP7_75t_SL g1989 ( 
.A(n_1548),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_1719),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_827),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1449),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_863),
.Y(n_1993)
);

INVx1_ASAP7_75t_SL g1994 ( 
.A(n_975),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1683),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1603),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_816),
.Y(n_1997)
);

CKINVDCx20_ASAP7_75t_R g1998 ( 
.A(n_81),
.Y(n_1998)
);

BUFx8_ASAP7_75t_SL g1999 ( 
.A(n_628),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1508),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_1119),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_1622),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_813),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1782),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_267),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_1412),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1342),
.Y(n_2007)
);

CKINVDCx20_ASAP7_75t_R g2008 ( 
.A(n_1597),
.Y(n_2008)
);

CKINVDCx5p33_ASAP7_75t_R g2009 ( 
.A(n_1270),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_1717),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_1694),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_1590),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1702),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_873),
.Y(n_2014)
);

INVx1_ASAP7_75t_SL g2015 ( 
.A(n_1008),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_273),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1143),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_190),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_827),
.Y(n_2019)
);

CKINVDCx5p33_ASAP7_75t_R g2020 ( 
.A(n_1522),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_1673),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_1360),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1763),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_555),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_994),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_49),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1336),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1648),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_957),
.Y(n_2029)
);

CKINVDCx20_ASAP7_75t_R g2030 ( 
.A(n_1772),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1706),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_358),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_1574),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_784),
.Y(n_2034)
);

CKINVDCx5p33_ASAP7_75t_R g2035 ( 
.A(n_1337),
.Y(n_2035)
);

BUFx6f_ASAP7_75t_L g2036 ( 
.A(n_837),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_1110),
.Y(n_2037)
);

BUFx10_ASAP7_75t_L g2038 ( 
.A(n_805),
.Y(n_2038)
);

BUFx3_ASAP7_75t_L g2039 ( 
.A(n_356),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_172),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_189),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_1711),
.Y(n_2042)
);

CKINVDCx20_ASAP7_75t_R g2043 ( 
.A(n_1249),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1486),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1244),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_1707),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_35),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_886),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_43),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1135),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_104),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_697),
.Y(n_2052)
);

CKINVDCx5p33_ASAP7_75t_R g2053 ( 
.A(n_1362),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_L g2054 ( 
.A(n_1587),
.Y(n_2054)
);

BUFx6f_ASAP7_75t_L g2055 ( 
.A(n_1524),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_229),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1197),
.Y(n_2057)
);

BUFx3_ASAP7_75t_L g2058 ( 
.A(n_1730),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1225),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1685),
.Y(n_2060)
);

INVx1_ASAP7_75t_SL g2061 ( 
.A(n_888),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_1644),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1787),
.Y(n_2063)
);

CKINVDCx5p33_ASAP7_75t_R g2064 ( 
.A(n_90),
.Y(n_2064)
);

BUFx3_ASAP7_75t_L g2065 ( 
.A(n_189),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_620),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_22),
.Y(n_2067)
);

CKINVDCx5p33_ASAP7_75t_R g2068 ( 
.A(n_1272),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_1164),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1205),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1592),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_469),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1305),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1701),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_209),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_1599),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_628),
.Y(n_2077)
);

BUFx10_ASAP7_75t_L g2078 ( 
.A(n_1727),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_866),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_945),
.Y(n_2080)
);

INVx1_ASAP7_75t_SL g2081 ( 
.A(n_106),
.Y(n_2081)
);

BUFx2_ASAP7_75t_L g2082 ( 
.A(n_1782),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_971),
.Y(n_2083)
);

CKINVDCx20_ASAP7_75t_R g2084 ( 
.A(n_682),
.Y(n_2084)
);

CKINVDCx5p33_ASAP7_75t_R g2085 ( 
.A(n_1785),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1563),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_10),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1546),
.Y(n_2088)
);

CKINVDCx20_ASAP7_75t_R g2089 ( 
.A(n_508),
.Y(n_2089)
);

CKINVDCx5p33_ASAP7_75t_R g2090 ( 
.A(n_385),
.Y(n_2090)
);

BUFx10_ASAP7_75t_L g2091 ( 
.A(n_1125),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1541),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_393),
.Y(n_2093)
);

CKINVDCx5p33_ASAP7_75t_R g2094 ( 
.A(n_1750),
.Y(n_2094)
);

BUFx6f_ASAP7_75t_L g2095 ( 
.A(n_1017),
.Y(n_2095)
);

BUFx6f_ASAP7_75t_L g2096 ( 
.A(n_1402),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_315),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_971),
.Y(n_2098)
);

CKINVDCx5p33_ASAP7_75t_R g2099 ( 
.A(n_1044),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_1489),
.Y(n_2100)
);

CKINVDCx5p33_ASAP7_75t_R g2101 ( 
.A(n_1450),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1060),
.Y(n_2102)
);

CKINVDCx5p33_ASAP7_75t_R g2103 ( 
.A(n_261),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_1658),
.Y(n_2104)
);

INVx1_ASAP7_75t_SL g2105 ( 
.A(n_1386),
.Y(n_2105)
);

CKINVDCx5p33_ASAP7_75t_R g2106 ( 
.A(n_1596),
.Y(n_2106)
);

CKINVDCx5p33_ASAP7_75t_R g2107 ( 
.A(n_1209),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_69),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_151),
.Y(n_2109)
);

BUFx5_ASAP7_75t_L g2110 ( 
.A(n_807),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1757),
.Y(n_2111)
);

CKINVDCx5p33_ASAP7_75t_R g2112 ( 
.A(n_1617),
.Y(n_2112)
);

INVx1_ASAP7_75t_SL g2113 ( 
.A(n_440),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_963),
.Y(n_2114)
);

CKINVDCx5p33_ASAP7_75t_R g2115 ( 
.A(n_1189),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_411),
.Y(n_2116)
);

CKINVDCx5p33_ASAP7_75t_R g2117 ( 
.A(n_1553),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_578),
.Y(n_2118)
);

CKINVDCx5p33_ASAP7_75t_R g2119 ( 
.A(n_1466),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1090),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1611),
.Y(n_2121)
);

CKINVDCx20_ASAP7_75t_R g2122 ( 
.A(n_400),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1613),
.Y(n_2123)
);

CKINVDCx5p33_ASAP7_75t_R g2124 ( 
.A(n_699),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1470),
.Y(n_2125)
);

CKINVDCx20_ASAP7_75t_R g2126 ( 
.A(n_1327),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_661),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1350),
.Y(n_2128)
);

CKINVDCx5p33_ASAP7_75t_R g2129 ( 
.A(n_130),
.Y(n_2129)
);

CKINVDCx5p33_ASAP7_75t_R g2130 ( 
.A(n_212),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1722),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1593),
.Y(n_2132)
);

CKINVDCx5p33_ASAP7_75t_R g2133 ( 
.A(n_612),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_737),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1561),
.Y(n_2135)
);

INVx1_ASAP7_75t_SL g2136 ( 
.A(n_237),
.Y(n_2136)
);

CKINVDCx5p33_ASAP7_75t_R g2137 ( 
.A(n_1603),
.Y(n_2137)
);

CKINVDCx5p33_ASAP7_75t_R g2138 ( 
.A(n_1675),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1260),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1748),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_592),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_967),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_1062),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_838),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_560),
.Y(n_2145)
);

CKINVDCx5p33_ASAP7_75t_R g2146 ( 
.A(n_29),
.Y(n_2146)
);

CKINVDCx5p33_ASAP7_75t_R g2147 ( 
.A(n_158),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_1667),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_566),
.Y(n_2149)
);

CKINVDCx5p33_ASAP7_75t_R g2150 ( 
.A(n_382),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1790),
.Y(n_2151)
);

CKINVDCx5p33_ASAP7_75t_R g2152 ( 
.A(n_794),
.Y(n_2152)
);

CKINVDCx5p33_ASAP7_75t_R g2153 ( 
.A(n_1349),
.Y(n_2153)
);

CKINVDCx5p33_ASAP7_75t_R g2154 ( 
.A(n_1290),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1033),
.Y(n_2155)
);

CKINVDCx5p33_ASAP7_75t_R g2156 ( 
.A(n_1054),
.Y(n_2156)
);

BUFx2_ASAP7_75t_L g2157 ( 
.A(n_725),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_775),
.Y(n_2158)
);

CKINVDCx5p33_ASAP7_75t_R g2159 ( 
.A(n_1656),
.Y(n_2159)
);

BUFx10_ASAP7_75t_L g2160 ( 
.A(n_125),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_446),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_466),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_1296),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_840),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_1596),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1478),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_161),
.Y(n_2167)
);

BUFx3_ASAP7_75t_L g2168 ( 
.A(n_1646),
.Y(n_2168)
);

CKINVDCx5p33_ASAP7_75t_R g2169 ( 
.A(n_1726),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_833),
.Y(n_2170)
);

CKINVDCx5p33_ASAP7_75t_R g2171 ( 
.A(n_324),
.Y(n_2171)
);

CKINVDCx20_ASAP7_75t_R g2172 ( 
.A(n_1155),
.Y(n_2172)
);

CKINVDCx5p33_ASAP7_75t_R g2173 ( 
.A(n_358),
.Y(n_2173)
);

CKINVDCx5p33_ASAP7_75t_R g2174 ( 
.A(n_1791),
.Y(n_2174)
);

CKINVDCx5p33_ASAP7_75t_R g2175 ( 
.A(n_912),
.Y(n_2175)
);

CKINVDCx5p33_ASAP7_75t_R g2176 ( 
.A(n_735),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_921),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_L g2178 ( 
.A(n_1456),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_191),
.Y(n_2179)
);

CKINVDCx20_ASAP7_75t_R g2180 ( 
.A(n_102),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_778),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_1308),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_1470),
.Y(n_2183)
);

BUFx6f_ASAP7_75t_L g2184 ( 
.A(n_688),
.Y(n_2184)
);

CKINVDCx20_ASAP7_75t_R g2185 ( 
.A(n_1715),
.Y(n_2185)
);

CKINVDCx5p33_ASAP7_75t_R g2186 ( 
.A(n_1284),
.Y(n_2186)
);

CKINVDCx5p33_ASAP7_75t_R g2187 ( 
.A(n_831),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_483),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_831),
.Y(n_2189)
);

BUFx6f_ASAP7_75t_L g2190 ( 
.A(n_1558),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_804),
.Y(n_2191)
);

BUFx6f_ASAP7_75t_L g2192 ( 
.A(n_1701),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_853),
.Y(n_2193)
);

INVxp33_ASAP7_75t_L g2194 ( 
.A(n_915),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_130),
.Y(n_2195)
);

CKINVDCx5p33_ASAP7_75t_R g2196 ( 
.A(n_946),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_160),
.Y(n_2197)
);

BUFx10_ASAP7_75t_L g2198 ( 
.A(n_508),
.Y(n_2198)
);

CKINVDCx20_ASAP7_75t_R g2199 ( 
.A(n_1414),
.Y(n_2199)
);

CKINVDCx20_ASAP7_75t_R g2200 ( 
.A(n_1653),
.Y(n_2200)
);

CKINVDCx5p33_ASAP7_75t_R g2201 ( 
.A(n_1629),
.Y(n_2201)
);

CKINVDCx20_ASAP7_75t_R g2202 ( 
.A(n_380),
.Y(n_2202)
);

HB1xp67_ASAP7_75t_L g2203 ( 
.A(n_175),
.Y(n_2203)
);

CKINVDCx14_ASAP7_75t_R g2204 ( 
.A(n_1081),
.Y(n_2204)
);

CKINVDCx5p33_ASAP7_75t_R g2205 ( 
.A(n_1731),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_1550),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1399),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_885),
.Y(n_2208)
);

CKINVDCx5p33_ASAP7_75t_R g2209 ( 
.A(n_1340),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_1684),
.Y(n_2210)
);

BUFx6f_ASAP7_75t_L g2211 ( 
.A(n_1346),
.Y(n_2211)
);

BUFx10_ASAP7_75t_L g2212 ( 
.A(n_373),
.Y(n_2212)
);

BUFx10_ASAP7_75t_L g2213 ( 
.A(n_894),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_1499),
.Y(n_2214)
);

BUFx2_ASAP7_75t_L g2215 ( 
.A(n_1595),
.Y(n_2215)
);

CKINVDCx5p33_ASAP7_75t_R g2216 ( 
.A(n_123),
.Y(n_2216)
);

CKINVDCx5p33_ASAP7_75t_R g2217 ( 
.A(n_395),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_1612),
.Y(n_2218)
);

CKINVDCx20_ASAP7_75t_R g2219 ( 
.A(n_1092),
.Y(n_2219)
);

CKINVDCx20_ASAP7_75t_R g2220 ( 
.A(n_1670),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_1668),
.Y(n_2221)
);

CKINVDCx5p33_ASAP7_75t_R g2222 ( 
.A(n_617),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_1342),
.Y(n_2223)
);

BUFx10_ASAP7_75t_L g2224 ( 
.A(n_187),
.Y(n_2224)
);

CKINVDCx5p33_ASAP7_75t_R g2225 ( 
.A(n_1544),
.Y(n_2225)
);

CKINVDCx5p33_ASAP7_75t_R g2226 ( 
.A(n_1150),
.Y(n_2226)
);

BUFx2_ASAP7_75t_SL g2227 ( 
.A(n_712),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_1386),
.Y(n_2228)
);

BUFx2_ASAP7_75t_L g2229 ( 
.A(n_991),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_292),
.Y(n_2230)
);

CKINVDCx5p33_ASAP7_75t_R g2231 ( 
.A(n_1324),
.Y(n_2231)
);

BUFx10_ASAP7_75t_L g2232 ( 
.A(n_1286),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_738),
.Y(n_2233)
);

INVx2_ASAP7_75t_SL g2234 ( 
.A(n_1402),
.Y(n_2234)
);

INVx1_ASAP7_75t_SL g2235 ( 
.A(n_1630),
.Y(n_2235)
);

CKINVDCx5p33_ASAP7_75t_R g2236 ( 
.A(n_1021),
.Y(n_2236)
);

BUFx10_ASAP7_75t_L g2237 ( 
.A(n_1131),
.Y(n_2237)
);

CKINVDCx5p33_ASAP7_75t_R g2238 ( 
.A(n_1686),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_470),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1754),
.Y(n_2240)
);

CKINVDCx5p33_ASAP7_75t_R g2241 ( 
.A(n_1120),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_997),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1600),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_1246),
.Y(n_2244)
);

BUFx3_ASAP7_75t_L g2245 ( 
.A(n_505),
.Y(n_2245)
);

CKINVDCx5p33_ASAP7_75t_R g2246 ( 
.A(n_563),
.Y(n_2246)
);

CKINVDCx5p33_ASAP7_75t_R g2247 ( 
.A(n_27),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_1538),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_1634),
.Y(n_2249)
);

BUFx10_ASAP7_75t_L g2250 ( 
.A(n_1238),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_1647),
.Y(n_2251)
);

CKINVDCx5p33_ASAP7_75t_R g2252 ( 
.A(n_64),
.Y(n_2252)
);

CKINVDCx5p33_ASAP7_75t_R g2253 ( 
.A(n_1554),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1709),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_404),
.Y(n_2255)
);

BUFx6f_ASAP7_75t_L g2256 ( 
.A(n_749),
.Y(n_2256)
);

CKINVDCx5p33_ASAP7_75t_R g2257 ( 
.A(n_1614),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1788),
.Y(n_2258)
);

CKINVDCx5p33_ASAP7_75t_R g2259 ( 
.A(n_1367),
.Y(n_2259)
);

BUFx3_ASAP7_75t_L g2260 ( 
.A(n_530),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_1546),
.Y(n_2261)
);

CKINVDCx5p33_ASAP7_75t_R g2262 ( 
.A(n_721),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_266),
.Y(n_2263)
);

BUFx8_ASAP7_75t_SL g2264 ( 
.A(n_748),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1089),
.Y(n_2265)
);

CKINVDCx5p33_ASAP7_75t_R g2266 ( 
.A(n_1792),
.Y(n_2266)
);

CKINVDCx16_ASAP7_75t_R g2267 ( 
.A(n_1627),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1328),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1549),
.Y(n_2269)
);

CKINVDCx5p33_ASAP7_75t_R g2270 ( 
.A(n_71),
.Y(n_2270)
);

CKINVDCx5p33_ASAP7_75t_R g2271 ( 
.A(n_741),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1735),
.Y(n_2272)
);

CKINVDCx5p33_ASAP7_75t_R g2273 ( 
.A(n_954),
.Y(n_2273)
);

INVx1_ASAP7_75t_SL g2274 ( 
.A(n_1728),
.Y(n_2274)
);

CKINVDCx5p33_ASAP7_75t_R g2275 ( 
.A(n_705),
.Y(n_2275)
);

BUFx3_ASAP7_75t_L g2276 ( 
.A(n_611),
.Y(n_2276)
);

INVx2_ASAP7_75t_SL g2277 ( 
.A(n_326),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_809),
.Y(n_2278)
);

CKINVDCx5p33_ASAP7_75t_R g2279 ( 
.A(n_651),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1695),
.Y(n_2280)
);

CKINVDCx5p33_ASAP7_75t_R g2281 ( 
.A(n_250),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_843),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_61),
.Y(n_2283)
);

CKINVDCx5p33_ASAP7_75t_R g2284 ( 
.A(n_1703),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_742),
.Y(n_2285)
);

BUFx10_ASAP7_75t_L g2286 ( 
.A(n_611),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_940),
.Y(n_2287)
);

CKINVDCx5p33_ASAP7_75t_R g2288 ( 
.A(n_603),
.Y(n_2288)
);

BUFx6f_ASAP7_75t_L g2289 ( 
.A(n_909),
.Y(n_2289)
);

INVx2_ASAP7_75t_SL g2290 ( 
.A(n_1000),
.Y(n_2290)
);

CKINVDCx5p33_ASAP7_75t_R g2291 ( 
.A(n_365),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_190),
.Y(n_2292)
);

CKINVDCx5p33_ASAP7_75t_R g2293 ( 
.A(n_955),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_526),
.Y(n_2294)
);

BUFx5_ASAP7_75t_L g2295 ( 
.A(n_855),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_1688),
.Y(n_2296)
);

CKINVDCx5p33_ASAP7_75t_R g2297 ( 
.A(n_1251),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1514),
.Y(n_2298)
);

CKINVDCx5p33_ASAP7_75t_R g2299 ( 
.A(n_1698),
.Y(n_2299)
);

CKINVDCx5p33_ASAP7_75t_R g2300 ( 
.A(n_88),
.Y(n_2300)
);

BUFx3_ASAP7_75t_L g2301 ( 
.A(n_1664),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_1666),
.Y(n_2302)
);

CKINVDCx5p33_ASAP7_75t_R g2303 ( 
.A(n_1588),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_203),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_493),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_877),
.Y(n_2306)
);

CKINVDCx5p33_ASAP7_75t_R g2307 ( 
.A(n_1660),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_1085),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1464),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_1571),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1615),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_96),
.Y(n_2312)
);

CKINVDCx5p33_ASAP7_75t_R g2313 ( 
.A(n_571),
.Y(n_2313)
);

CKINVDCx5p33_ASAP7_75t_R g2314 ( 
.A(n_481),
.Y(n_2314)
);

CKINVDCx20_ASAP7_75t_R g2315 ( 
.A(n_1275),
.Y(n_2315)
);

CKINVDCx5p33_ASAP7_75t_R g2316 ( 
.A(n_1777),
.Y(n_2316)
);

CKINVDCx5p33_ASAP7_75t_R g2317 ( 
.A(n_651),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_406),
.Y(n_2318)
);

CKINVDCx5p33_ASAP7_75t_R g2319 ( 
.A(n_872),
.Y(n_2319)
);

BUFx6f_ASAP7_75t_L g2320 ( 
.A(n_1561),
.Y(n_2320)
);

CKINVDCx5p33_ASAP7_75t_R g2321 ( 
.A(n_937),
.Y(n_2321)
);

CKINVDCx5p33_ASAP7_75t_R g2322 ( 
.A(n_521),
.Y(n_2322)
);

CKINVDCx5p33_ASAP7_75t_R g2323 ( 
.A(n_59),
.Y(n_2323)
);

CKINVDCx5p33_ASAP7_75t_R g2324 ( 
.A(n_1544),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1154),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_1422),
.Y(n_2326)
);

CKINVDCx20_ASAP7_75t_R g2327 ( 
.A(n_1010),
.Y(n_2327)
);

CKINVDCx5p33_ASAP7_75t_R g2328 ( 
.A(n_1521),
.Y(n_2328)
);

CKINVDCx16_ASAP7_75t_R g2329 ( 
.A(n_1712),
.Y(n_2329)
);

BUFx6f_ASAP7_75t_L g2330 ( 
.A(n_1682),
.Y(n_2330)
);

CKINVDCx20_ASAP7_75t_R g2331 ( 
.A(n_1602),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_778),
.Y(n_2332)
);

CKINVDCx5p33_ASAP7_75t_R g2333 ( 
.A(n_1729),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_488),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1714),
.Y(n_2335)
);

CKINVDCx5p33_ASAP7_75t_R g2336 ( 
.A(n_1713),
.Y(n_2336)
);

CKINVDCx5p33_ASAP7_75t_R g2337 ( 
.A(n_457),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1022),
.Y(n_2338)
);

BUFx6f_ASAP7_75t_L g2339 ( 
.A(n_1547),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_889),
.Y(n_2340)
);

CKINVDCx5p33_ASAP7_75t_R g2341 ( 
.A(n_528),
.Y(n_2341)
);

CKINVDCx5p33_ASAP7_75t_R g2342 ( 
.A(n_1725),
.Y(n_2342)
);

CKINVDCx20_ASAP7_75t_R g2343 ( 
.A(n_144),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_650),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_1496),
.Y(n_2345)
);

CKINVDCx16_ASAP7_75t_R g2346 ( 
.A(n_1697),
.Y(n_2346)
);

CKINVDCx5p33_ASAP7_75t_R g2347 ( 
.A(n_1692),
.Y(n_2347)
);

BUFx10_ASAP7_75t_L g2348 ( 
.A(n_1016),
.Y(n_2348)
);

CKINVDCx16_ASAP7_75t_R g2349 ( 
.A(n_1475),
.Y(n_2349)
);

CKINVDCx5p33_ASAP7_75t_R g2350 ( 
.A(n_1650),
.Y(n_2350)
);

CKINVDCx5p33_ASAP7_75t_R g2351 ( 
.A(n_1791),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_1293),
.Y(n_2352)
);

CKINVDCx5p33_ASAP7_75t_R g2353 ( 
.A(n_415),
.Y(n_2353)
);

CKINVDCx5p33_ASAP7_75t_R g2354 ( 
.A(n_1632),
.Y(n_2354)
);

CKINVDCx5p33_ASAP7_75t_R g2355 ( 
.A(n_1643),
.Y(n_2355)
);

BUFx6f_ASAP7_75t_L g2356 ( 
.A(n_668),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_1534),
.Y(n_2357)
);

BUFx10_ASAP7_75t_L g2358 ( 
.A(n_1538),
.Y(n_2358)
);

BUFx2_ASAP7_75t_L g2359 ( 
.A(n_1271),
.Y(n_2359)
);

CKINVDCx5p33_ASAP7_75t_R g2360 ( 
.A(n_990),
.Y(n_2360)
);

CKINVDCx5p33_ASAP7_75t_R g2361 ( 
.A(n_1634),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_1235),
.Y(n_2362)
);

BUFx6f_ASAP7_75t_L g2363 ( 
.A(n_459),
.Y(n_2363)
);

CKINVDCx5p33_ASAP7_75t_R g2364 ( 
.A(n_681),
.Y(n_2364)
);

CKINVDCx20_ASAP7_75t_R g2365 ( 
.A(n_610),
.Y(n_2365)
);

CKINVDCx5p33_ASAP7_75t_R g2366 ( 
.A(n_459),
.Y(n_2366)
);

CKINVDCx20_ASAP7_75t_R g2367 ( 
.A(n_287),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_742),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_465),
.Y(n_2369)
);

CKINVDCx5p33_ASAP7_75t_R g2370 ( 
.A(n_67),
.Y(n_2370)
);

CKINVDCx5p33_ASAP7_75t_R g2371 ( 
.A(n_1581),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_1416),
.Y(n_2372)
);

CKINVDCx5p33_ASAP7_75t_R g2373 ( 
.A(n_494),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_410),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_1661),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_151),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_1329),
.Y(n_2377)
);

BUFx10_ASAP7_75t_L g2378 ( 
.A(n_1035),
.Y(n_2378)
);

INVx3_ASAP7_75t_L g2379 ( 
.A(n_545),
.Y(n_2379)
);

BUFx3_ASAP7_75t_L g2380 ( 
.A(n_351),
.Y(n_2380)
);

CKINVDCx5p33_ASAP7_75t_R g2381 ( 
.A(n_594),
.Y(n_2381)
);

BUFx3_ASAP7_75t_L g2382 ( 
.A(n_1645),
.Y(n_2382)
);

CKINVDCx5p33_ASAP7_75t_R g2383 ( 
.A(n_1565),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_1323),
.Y(n_2384)
);

CKINVDCx5p33_ASAP7_75t_R g2385 ( 
.A(n_1425),
.Y(n_2385)
);

BUFx3_ASAP7_75t_L g2386 ( 
.A(n_1086),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_799),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_1573),
.Y(n_2388)
);

CKINVDCx5p33_ASAP7_75t_R g2389 ( 
.A(n_1289),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_1381),
.Y(n_2390)
);

CKINVDCx5p33_ASAP7_75t_R g2391 ( 
.A(n_1737),
.Y(n_2391)
);

BUFx5_ASAP7_75t_L g2392 ( 
.A(n_1657),
.Y(n_2392)
);

CKINVDCx5p33_ASAP7_75t_R g2393 ( 
.A(n_159),
.Y(n_2393)
);

CKINVDCx5p33_ASAP7_75t_R g2394 ( 
.A(n_80),
.Y(n_2394)
);

CKINVDCx5p33_ASAP7_75t_R g2395 ( 
.A(n_568),
.Y(n_2395)
);

CKINVDCx5p33_ASAP7_75t_R g2396 ( 
.A(n_1353),
.Y(n_2396)
);

CKINVDCx20_ASAP7_75t_R g2397 ( 
.A(n_855),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_1421),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_141),
.Y(n_2399)
);

CKINVDCx5p33_ASAP7_75t_R g2400 ( 
.A(n_489),
.Y(n_2400)
);

CKINVDCx5p33_ASAP7_75t_R g2401 ( 
.A(n_974),
.Y(n_2401)
);

CKINVDCx5p33_ASAP7_75t_R g2402 ( 
.A(n_363),
.Y(n_2402)
);

CKINVDCx5p33_ASAP7_75t_R g2403 ( 
.A(n_1661),
.Y(n_2403)
);

CKINVDCx5p33_ASAP7_75t_R g2404 ( 
.A(n_1665),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_737),
.Y(n_2405)
);

BUFx6f_ASAP7_75t_L g2406 ( 
.A(n_1244),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_384),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_64),
.Y(n_2408)
);

BUFx6f_ASAP7_75t_L g2409 ( 
.A(n_815),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_879),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_1674),
.Y(n_2411)
);

BUFx10_ASAP7_75t_L g2412 ( 
.A(n_487),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_1657),
.Y(n_2413)
);

BUFx10_ASAP7_75t_L g2414 ( 
.A(n_523),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_595),
.Y(n_2415)
);

CKINVDCx5p33_ASAP7_75t_R g2416 ( 
.A(n_1086),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_938),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_1671),
.Y(n_2418)
);

BUFx6f_ASAP7_75t_L g2419 ( 
.A(n_679),
.Y(n_2419)
);

CKINVDCx5p33_ASAP7_75t_R g2420 ( 
.A(n_453),
.Y(n_2420)
);

CKINVDCx5p33_ASAP7_75t_R g2421 ( 
.A(n_1332),
.Y(n_2421)
);

CKINVDCx5p33_ASAP7_75t_R g2422 ( 
.A(n_1675),
.Y(n_2422)
);

BUFx3_ASAP7_75t_L g2423 ( 
.A(n_1387),
.Y(n_2423)
);

CKINVDCx20_ASAP7_75t_R g2424 ( 
.A(n_82),
.Y(n_2424)
);

CKINVDCx5p33_ASAP7_75t_R g2425 ( 
.A(n_1705),
.Y(n_2425)
);

CKINVDCx5p33_ASAP7_75t_R g2426 ( 
.A(n_1277),
.Y(n_2426)
);

CKINVDCx5p33_ASAP7_75t_R g2427 ( 
.A(n_945),
.Y(n_2427)
);

CKINVDCx20_ASAP7_75t_R g2428 ( 
.A(n_640),
.Y(n_2428)
);

BUFx3_ASAP7_75t_L g2429 ( 
.A(n_1137),
.Y(n_2429)
);

CKINVDCx5p33_ASAP7_75t_R g2430 ( 
.A(n_1689),
.Y(n_2430)
);

CKINVDCx5p33_ASAP7_75t_R g2431 ( 
.A(n_1633),
.Y(n_2431)
);

CKINVDCx5p33_ASAP7_75t_R g2432 ( 
.A(n_1490),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_115),
.Y(n_2433)
);

CKINVDCx5p33_ASAP7_75t_R g2434 ( 
.A(n_898),
.Y(n_2434)
);

BUFx3_ASAP7_75t_L g2435 ( 
.A(n_988),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_857),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_137),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_1577),
.Y(n_2438)
);

CKINVDCx5p33_ASAP7_75t_R g2439 ( 
.A(n_282),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_57),
.Y(n_2440)
);

CKINVDCx20_ASAP7_75t_R g2441 ( 
.A(n_1161),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_574),
.Y(n_2442)
);

CKINVDCx5p33_ASAP7_75t_R g2443 ( 
.A(n_1253),
.Y(n_2443)
);

CKINVDCx5p33_ASAP7_75t_R g2444 ( 
.A(n_1480),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_1200),
.Y(n_2445)
);

CKINVDCx14_ASAP7_75t_R g2446 ( 
.A(n_143),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_1606),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_22),
.Y(n_2448)
);

BUFx10_ASAP7_75t_L g2449 ( 
.A(n_356),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_606),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_907),
.Y(n_2451)
);

CKINVDCx5p33_ASAP7_75t_R g2452 ( 
.A(n_739),
.Y(n_2452)
);

CKINVDCx20_ASAP7_75t_R g2453 ( 
.A(n_635),
.Y(n_2453)
);

BUFx3_ASAP7_75t_L g2454 ( 
.A(n_1585),
.Y(n_2454)
);

CKINVDCx5p33_ASAP7_75t_R g2455 ( 
.A(n_1516),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_1672),
.Y(n_2456)
);

BUFx10_ASAP7_75t_L g2457 ( 
.A(n_450),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_108),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_1559),
.Y(n_2459)
);

CKINVDCx5p33_ASAP7_75t_R g2460 ( 
.A(n_729),
.Y(n_2460)
);

CKINVDCx5p33_ASAP7_75t_R g2461 ( 
.A(n_1360),
.Y(n_2461)
);

CKINVDCx5p33_ASAP7_75t_R g2462 ( 
.A(n_1618),
.Y(n_2462)
);

CKINVDCx5p33_ASAP7_75t_R g2463 ( 
.A(n_703),
.Y(n_2463)
);

CKINVDCx5p33_ASAP7_75t_R g2464 ( 
.A(n_1564),
.Y(n_2464)
);

CKINVDCx20_ASAP7_75t_R g2465 ( 
.A(n_1168),
.Y(n_2465)
);

CKINVDCx20_ASAP7_75t_R g2466 ( 
.A(n_1677),
.Y(n_2466)
);

CKINVDCx5p33_ASAP7_75t_R g2467 ( 
.A(n_1589),
.Y(n_2467)
);

BUFx6f_ASAP7_75t_L g2468 ( 
.A(n_1556),
.Y(n_2468)
);

CKINVDCx5p33_ASAP7_75t_R g2469 ( 
.A(n_1225),
.Y(n_2469)
);

HB1xp67_ASAP7_75t_L g2470 ( 
.A(n_1228),
.Y(n_2470)
);

CKINVDCx5p33_ASAP7_75t_R g2471 ( 
.A(n_745),
.Y(n_2471)
);

INVx1_ASAP7_75t_SL g2472 ( 
.A(n_1655),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_1649),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_220),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_1045),
.Y(n_2475)
);

CKINVDCx5p33_ASAP7_75t_R g2476 ( 
.A(n_1152),
.Y(n_2476)
);

BUFx6f_ASAP7_75t_L g2477 ( 
.A(n_1299),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_984),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_1583),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_883),
.Y(n_2480)
);

CKINVDCx5p33_ASAP7_75t_R g2481 ( 
.A(n_1721),
.Y(n_2481)
);

BUFx3_ASAP7_75t_L g2482 ( 
.A(n_1551),
.Y(n_2482)
);

CKINVDCx5p33_ASAP7_75t_R g2483 ( 
.A(n_1716),
.Y(n_2483)
);

CKINVDCx5p33_ASAP7_75t_R g2484 ( 
.A(n_73),
.Y(n_2484)
);

CKINVDCx5p33_ASAP7_75t_R g2485 ( 
.A(n_830),
.Y(n_2485)
);

CKINVDCx5p33_ASAP7_75t_R g2486 ( 
.A(n_1181),
.Y(n_2486)
);

CKINVDCx5p33_ASAP7_75t_R g2487 ( 
.A(n_1097),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_821),
.Y(n_2488)
);

CKINVDCx5p33_ASAP7_75t_R g2489 ( 
.A(n_1690),
.Y(n_2489)
);

CKINVDCx5p33_ASAP7_75t_R g2490 ( 
.A(n_900),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_48),
.Y(n_2491)
);

BUFx5_ASAP7_75t_L g2492 ( 
.A(n_1700),
.Y(n_2492)
);

CKINVDCx20_ASAP7_75t_R g2493 ( 
.A(n_304),
.Y(n_2493)
);

CKINVDCx5p33_ASAP7_75t_R g2494 ( 
.A(n_1260),
.Y(n_2494)
);

INVx1_ASAP7_75t_SL g2495 ( 
.A(n_265),
.Y(n_2495)
);

CKINVDCx5p33_ASAP7_75t_R g2496 ( 
.A(n_752),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_1659),
.Y(n_2497)
);

CKINVDCx5p33_ASAP7_75t_R g2498 ( 
.A(n_1187),
.Y(n_2498)
);

CKINVDCx5p33_ASAP7_75t_R g2499 ( 
.A(n_405),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_967),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_637),
.Y(n_2501)
);

CKINVDCx5p33_ASAP7_75t_R g2502 ( 
.A(n_564),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_1651),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_162),
.Y(n_2504)
);

CKINVDCx16_ASAP7_75t_R g2505 ( 
.A(n_1591),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_1238),
.Y(n_2506)
);

CKINVDCx20_ASAP7_75t_R g2507 ( 
.A(n_1533),
.Y(n_2507)
);

CKINVDCx5p33_ASAP7_75t_R g2508 ( 
.A(n_228),
.Y(n_2508)
);

CKINVDCx5p33_ASAP7_75t_R g2509 ( 
.A(n_1631),
.Y(n_2509)
);

CKINVDCx5p33_ASAP7_75t_R g2510 ( 
.A(n_1602),
.Y(n_2510)
);

CKINVDCx5p33_ASAP7_75t_R g2511 ( 
.A(n_1628),
.Y(n_2511)
);

CKINVDCx5p33_ASAP7_75t_R g2512 ( 
.A(n_47),
.Y(n_2512)
);

BUFx10_ASAP7_75t_L g2513 ( 
.A(n_1115),
.Y(n_2513)
);

BUFx6f_ASAP7_75t_L g2514 ( 
.A(n_1578),
.Y(n_2514)
);

CKINVDCx5p33_ASAP7_75t_R g2515 ( 
.A(n_1579),
.Y(n_2515)
);

CKINVDCx20_ASAP7_75t_R g2516 ( 
.A(n_1584),
.Y(n_2516)
);

CKINVDCx20_ASAP7_75t_R g2517 ( 
.A(n_1696),
.Y(n_2517)
);

BUFx10_ASAP7_75t_L g2518 ( 
.A(n_582),
.Y(n_2518)
);

CKINVDCx5p33_ASAP7_75t_R g2519 ( 
.A(n_145),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_818),
.Y(n_2520)
);

CKINVDCx5p33_ASAP7_75t_R g2521 ( 
.A(n_219),
.Y(n_2521)
);

CKINVDCx16_ASAP7_75t_R g2522 ( 
.A(n_223),
.Y(n_2522)
);

CKINVDCx5p33_ASAP7_75t_R g2523 ( 
.A(n_1642),
.Y(n_2523)
);

CKINVDCx5p33_ASAP7_75t_R g2524 ( 
.A(n_1636),
.Y(n_2524)
);

BUFx6f_ASAP7_75t_L g2525 ( 
.A(n_1023),
.Y(n_2525)
);

CKINVDCx20_ASAP7_75t_R g2526 ( 
.A(n_1598),
.Y(n_2526)
);

CKINVDCx20_ASAP7_75t_R g2527 ( 
.A(n_1669),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_1788),
.Y(n_2528)
);

CKINVDCx5p33_ASAP7_75t_R g2529 ( 
.A(n_1685),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_1128),
.Y(n_2530)
);

BUFx2_ASAP7_75t_R g2531 ( 
.A(n_919),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_135),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_450),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_1586),
.Y(n_2534)
);

CKINVDCx5p33_ASAP7_75t_R g2535 ( 
.A(n_142),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_878),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_261),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_826),
.Y(n_2538)
);

CKINVDCx5p33_ASAP7_75t_R g2539 ( 
.A(n_153),
.Y(n_2539)
);

INVx2_ASAP7_75t_SL g2540 ( 
.A(n_949),
.Y(n_2540)
);

CKINVDCx20_ASAP7_75t_R g2541 ( 
.A(n_1601),
.Y(n_2541)
);

INVx2_ASAP7_75t_SL g2542 ( 
.A(n_458),
.Y(n_2542)
);

CKINVDCx16_ASAP7_75t_R g2543 ( 
.A(n_1025),
.Y(n_2543)
);

CKINVDCx20_ASAP7_75t_R g2544 ( 
.A(n_287),
.Y(n_2544)
);

CKINVDCx5p33_ASAP7_75t_R g2545 ( 
.A(n_1109),
.Y(n_2545)
);

CKINVDCx5p33_ASAP7_75t_R g2546 ( 
.A(n_788),
.Y(n_2546)
);

CKINVDCx20_ASAP7_75t_R g2547 ( 
.A(n_499),
.Y(n_2547)
);

BUFx6f_ASAP7_75t_L g2548 ( 
.A(n_1572),
.Y(n_2548)
);

CKINVDCx20_ASAP7_75t_R g2549 ( 
.A(n_1637),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_800),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_1218),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_203),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_1328),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_90),
.Y(n_2554)
);

CKINVDCx5p33_ASAP7_75t_R g2555 ( 
.A(n_1611),
.Y(n_2555)
);

CKINVDCx5p33_ASAP7_75t_R g2556 ( 
.A(n_580),
.Y(n_2556)
);

CKINVDCx5p33_ASAP7_75t_R g2557 ( 
.A(n_1162),
.Y(n_2557)
);

CKINVDCx5p33_ASAP7_75t_R g2558 ( 
.A(n_1570),
.Y(n_2558)
);

CKINVDCx16_ASAP7_75t_R g2559 ( 
.A(n_100),
.Y(n_2559)
);

CKINVDCx20_ASAP7_75t_R g2560 ( 
.A(n_240),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_1686),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_1576),
.Y(n_2562)
);

CKINVDCx14_ASAP7_75t_R g2563 ( 
.A(n_1148),
.Y(n_2563)
);

CKINVDCx5p33_ASAP7_75t_R g2564 ( 
.A(n_463),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_1167),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_1582),
.Y(n_2566)
);

CKINVDCx5p33_ASAP7_75t_R g2567 ( 
.A(n_23),
.Y(n_2567)
);

CKINVDCx20_ASAP7_75t_R g2568 ( 
.A(n_219),
.Y(n_2568)
);

BUFx6f_ASAP7_75t_L g2569 ( 
.A(n_1331),
.Y(n_2569)
);

CKINVDCx20_ASAP7_75t_R g2570 ( 
.A(n_800),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_1073),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_1438),
.Y(n_2572)
);

CKINVDCx5p33_ASAP7_75t_R g2573 ( 
.A(n_87),
.Y(n_2573)
);

CKINVDCx5p33_ASAP7_75t_R g2574 ( 
.A(n_736),
.Y(n_2574)
);

CKINVDCx5p33_ASAP7_75t_R g2575 ( 
.A(n_1653),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_1557),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_415),
.Y(n_2577)
);

CKINVDCx5p33_ASAP7_75t_R g2578 ( 
.A(n_1476),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_1452),
.Y(n_2579)
);

CKINVDCx14_ASAP7_75t_R g2580 ( 
.A(n_1718),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_1198),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_1159),
.Y(n_2582)
);

BUFx10_ASAP7_75t_L g2583 ( 
.A(n_345),
.Y(n_2583)
);

BUFx10_ASAP7_75t_L g2584 ( 
.A(n_663),
.Y(n_2584)
);

BUFx6f_ASAP7_75t_L g2585 ( 
.A(n_112),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_1132),
.Y(n_2586)
);

CKINVDCx5p33_ASAP7_75t_R g2587 ( 
.A(n_198),
.Y(n_2587)
);

BUFx10_ASAP7_75t_L g2588 ( 
.A(n_949),
.Y(n_2588)
);

INVx1_ASAP7_75t_SL g2589 ( 
.A(n_1680),
.Y(n_2589)
);

CKINVDCx20_ASAP7_75t_R g2590 ( 
.A(n_213),
.Y(n_2590)
);

CKINVDCx5p33_ASAP7_75t_R g2591 ( 
.A(n_301),
.Y(n_2591)
);

CKINVDCx5p33_ASAP7_75t_R g2592 ( 
.A(n_932),
.Y(n_2592)
);

INVx2_ASAP7_75t_SL g2593 ( 
.A(n_1736),
.Y(n_2593)
);

HB1xp67_ASAP7_75t_L g2594 ( 
.A(n_355),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_1516),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_464),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_1792),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_1594),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_61),
.Y(n_2599)
);

CKINVDCx20_ASAP7_75t_R g2600 ( 
.A(n_1767),
.Y(n_2600)
);

CKINVDCx5p33_ASAP7_75t_R g2601 ( 
.A(n_1080),
.Y(n_2601)
);

CKINVDCx5p33_ASAP7_75t_R g2602 ( 
.A(n_596),
.Y(n_2602)
);

CKINVDCx5p33_ASAP7_75t_R g2603 ( 
.A(n_1513),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_601),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_952),
.Y(n_2605)
);

CKINVDCx5p33_ASAP7_75t_R g2606 ( 
.A(n_438),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_120),
.Y(n_2607)
);

CKINVDCx20_ASAP7_75t_R g2608 ( 
.A(n_751),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_575),
.Y(n_2609)
);

CKINVDCx5p33_ASAP7_75t_R g2610 ( 
.A(n_397),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_1204),
.Y(n_2611)
);

BUFx6f_ASAP7_75t_L g2612 ( 
.A(n_656),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_838),
.Y(n_2613)
);

CKINVDCx5p33_ASAP7_75t_R g2614 ( 
.A(n_1691),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_640),
.Y(n_2615)
);

CKINVDCx16_ASAP7_75t_R g2616 ( 
.A(n_1673),
.Y(n_2616)
);

CKINVDCx20_ASAP7_75t_R g2617 ( 
.A(n_617),
.Y(n_2617)
);

CKINVDCx5p33_ASAP7_75t_R g2618 ( 
.A(n_583),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_468),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_1329),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_288),
.Y(n_2621)
);

CKINVDCx5p33_ASAP7_75t_R g2622 ( 
.A(n_686),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_1181),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_418),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_414),
.Y(n_2625)
);

CKINVDCx5p33_ASAP7_75t_R g2626 ( 
.A(n_612),
.Y(n_2626)
);

CKINVDCx5p33_ASAP7_75t_R g2627 ( 
.A(n_1663),
.Y(n_2627)
);

CKINVDCx5p33_ASAP7_75t_R g2628 ( 
.A(n_664),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_710),
.Y(n_2629)
);

CKINVDCx5p33_ASAP7_75t_R g2630 ( 
.A(n_1309),
.Y(n_2630)
);

CKINVDCx5p33_ASAP7_75t_R g2631 ( 
.A(n_1391),
.Y(n_2631)
);

CKINVDCx5p33_ASAP7_75t_R g2632 ( 
.A(n_183),
.Y(n_2632)
);

CKINVDCx5p33_ASAP7_75t_R g2633 ( 
.A(n_764),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_1580),
.Y(n_2634)
);

CKINVDCx5p33_ASAP7_75t_R g2635 ( 
.A(n_268),
.Y(n_2635)
);

BUFx8_ASAP7_75t_SL g2636 ( 
.A(n_386),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_49),
.Y(n_2637)
);

CKINVDCx5p33_ASAP7_75t_R g2638 ( 
.A(n_923),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_1569),
.Y(n_2639)
);

CKINVDCx5p33_ASAP7_75t_R g2640 ( 
.A(n_1008),
.Y(n_2640)
);

CKINVDCx20_ASAP7_75t_R g2641 ( 
.A(n_449),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_14),
.Y(n_2642)
);

BUFx3_ASAP7_75t_L g2643 ( 
.A(n_1662),
.Y(n_2643)
);

CKINVDCx5p33_ASAP7_75t_R g2644 ( 
.A(n_1504),
.Y(n_2644)
);

CKINVDCx5p33_ASAP7_75t_R g2645 ( 
.A(n_826),
.Y(n_2645)
);

CKINVDCx5p33_ASAP7_75t_R g2646 ( 
.A(n_1491),
.Y(n_2646)
);

CKINVDCx5p33_ASAP7_75t_R g2647 ( 
.A(n_1316),
.Y(n_2647)
);

CKINVDCx5p33_ASAP7_75t_R g2648 ( 
.A(n_663),
.Y(n_2648)
);

CKINVDCx5p33_ASAP7_75t_R g2649 ( 
.A(n_169),
.Y(n_2649)
);

CKINVDCx5p33_ASAP7_75t_R g2650 ( 
.A(n_114),
.Y(n_2650)
);

INVx1_ASAP7_75t_SL g2651 ( 
.A(n_1796),
.Y(n_2651)
);

CKINVDCx5p33_ASAP7_75t_R g2652 ( 
.A(n_947),
.Y(n_2652)
);

BUFx3_ASAP7_75t_L g2653 ( 
.A(n_202),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_1532),
.Y(n_2654)
);

INVx1_ASAP7_75t_SL g2655 ( 
.A(n_1430),
.Y(n_2655)
);

CKINVDCx5p33_ASAP7_75t_R g2656 ( 
.A(n_1505),
.Y(n_2656)
);

INVx1_ASAP7_75t_SL g2657 ( 
.A(n_178),
.Y(n_2657)
);

CKINVDCx5p33_ASAP7_75t_R g2658 ( 
.A(n_823),
.Y(n_2658)
);

CKINVDCx5p33_ASAP7_75t_R g2659 ( 
.A(n_1165),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_1252),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_1568),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_939),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_354),
.Y(n_2663)
);

INVxp67_ASAP7_75t_L g2664 ( 
.A(n_1586),
.Y(n_2664)
);

CKINVDCx16_ASAP7_75t_R g2665 ( 
.A(n_1981),
.Y(n_2665)
);

INVxp67_ASAP7_75t_SL g2666 ( 
.A(n_2379),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_1959),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_1959),
.Y(n_2668)
);

INVxp67_ASAP7_75t_SL g2669 ( 
.A(n_2379),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_1959),
.Y(n_2670)
);

CKINVDCx5p33_ASAP7_75t_R g2671 ( 
.A(n_2636),
.Y(n_2671)
);

BUFx6f_ASAP7_75t_L g2672 ( 
.A(n_2041),
.Y(n_2672)
);

INVxp33_ASAP7_75t_SL g2673 ( 
.A(n_2093),
.Y(n_2673)
);

INVxp33_ASAP7_75t_SL g2674 ( 
.A(n_2203),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_1959),
.Y(n_2675)
);

CKINVDCx5p33_ASAP7_75t_R g2676 ( 
.A(n_1917),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_1959),
.Y(n_2677)
);

INVxp67_ASAP7_75t_SL g2678 ( 
.A(n_2594),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_1961),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_1961),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_1961),
.Y(n_2681)
);

INVxp67_ASAP7_75t_SL g2682 ( 
.A(n_2041),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_1961),
.Y(n_2683)
);

CKINVDCx5p33_ASAP7_75t_R g2684 ( 
.A(n_1999),
.Y(n_2684)
);

INVxp67_ASAP7_75t_L g2685 ( 
.A(n_1812),
.Y(n_2685)
);

INVxp33_ASAP7_75t_L g2686 ( 
.A(n_1819),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_1961),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_1797),
.Y(n_2688)
);

CKINVDCx16_ASAP7_75t_R g2689 ( 
.A(n_2522),
.Y(n_2689)
);

BUFx3_ASAP7_75t_L g2690 ( 
.A(n_1851),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_1797),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_1797),
.Y(n_2692)
);

HB1xp67_ASAP7_75t_L g2693 ( 
.A(n_2446),
.Y(n_2693)
);

CKINVDCx20_ASAP7_75t_R g2694 ( 
.A(n_1976),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_1797),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_2264),
.Y(n_2696)
);

INVxp67_ASAP7_75t_L g2697 ( 
.A(n_1897),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_1797),
.Y(n_2698)
);

INVxp33_ASAP7_75t_SL g2699 ( 
.A(n_1876),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_1885),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_1885),
.Y(n_2701)
);

CKINVDCx5p33_ASAP7_75t_R g2702 ( 
.A(n_2559),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_1885),
.Y(n_2703)
);

CKINVDCx5p33_ASAP7_75t_R g2704 ( 
.A(n_2204),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_1885),
.Y(n_2705)
);

BUFx3_ASAP7_75t_L g2706 ( 
.A(n_2039),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2110),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2110),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2110),
.Y(n_2709)
);

CKINVDCx5p33_ASAP7_75t_R g2710 ( 
.A(n_2563),
.Y(n_2710)
);

CKINVDCx5p33_ASAP7_75t_R g2711 ( 
.A(n_2580),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2295),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2295),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2295),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2295),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2392),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2392),
.Y(n_2717)
);

CKINVDCx5p33_ASAP7_75t_R g2718 ( 
.A(n_1801),
.Y(n_2718)
);

BUFx3_ASAP7_75t_L g2719 ( 
.A(n_2065),
.Y(n_2719)
);

CKINVDCx5p33_ASAP7_75t_R g2720 ( 
.A(n_1914),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2392),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2392),
.Y(n_2722)
);

CKINVDCx20_ASAP7_75t_R g2723 ( 
.A(n_1963),
.Y(n_2723)
);

CKINVDCx5p33_ASAP7_75t_R g2724 ( 
.A(n_2267),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2392),
.Y(n_2725)
);

INVx1_ASAP7_75t_SL g2726 ( 
.A(n_1904),
.Y(n_2726)
);

CKINVDCx20_ASAP7_75t_R g2727 ( 
.A(n_2329),
.Y(n_2727)
);

INVxp67_ASAP7_75t_L g2728 ( 
.A(n_1906),
.Y(n_2728)
);

INVxp67_ASAP7_75t_SL g2729 ( 
.A(n_2041),
.Y(n_2729)
);

INVxp67_ASAP7_75t_SL g2730 ( 
.A(n_2585),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2492),
.Y(n_2731)
);

CKINVDCx5p33_ASAP7_75t_R g2732 ( 
.A(n_2346),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2492),
.Y(n_2733)
);

INVxp67_ASAP7_75t_SL g2734 ( 
.A(n_2585),
.Y(n_2734)
);

CKINVDCx5p33_ASAP7_75t_R g2735 ( 
.A(n_2349),
.Y(n_2735)
);

CKINVDCx20_ASAP7_75t_R g2736 ( 
.A(n_2505),
.Y(n_2736)
);

CKINVDCx20_ASAP7_75t_R g2737 ( 
.A(n_2543),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2663),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_1816),
.Y(n_2739)
);

CKINVDCx5p33_ASAP7_75t_R g2740 ( 
.A(n_2616),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_1843),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_1861),
.Y(n_2742)
);

INVxp33_ASAP7_75t_L g2743 ( 
.A(n_1892),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_1944),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_1953),
.Y(n_2745)
);

BUFx2_ASAP7_75t_L g2746 ( 
.A(n_2082),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_1958),
.Y(n_2747)
);

CKINVDCx14_ASAP7_75t_R g2748 ( 
.A(n_2157),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_1982),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2005),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2047),
.Y(n_2751)
);

INVxp33_ASAP7_75t_SL g2752 ( 
.A(n_2470),
.Y(n_2752)
);

CKINVDCx5p33_ASAP7_75t_R g2753 ( 
.A(n_1807),
.Y(n_2753)
);

INVxp33_ASAP7_75t_SL g2754 ( 
.A(n_1815),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2051),
.Y(n_2755)
);

INVxp67_ASAP7_75t_SL g2756 ( 
.A(n_2653),
.Y(n_2756)
);

NOR2xp67_ASAP7_75t_L g2757 ( 
.A(n_2664),
.B(n_0),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2056),
.Y(n_2758)
);

CKINVDCx20_ASAP7_75t_R g2759 ( 
.A(n_1798),
.Y(n_2759)
);

INVxp33_ASAP7_75t_L g2760 ( 
.A(n_2215),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2067),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2087),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2097),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2108),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2167),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2179),
.Y(n_2766)
);

BUFx2_ASAP7_75t_SL g2767 ( 
.A(n_1973),
.Y(n_2767)
);

INVxp67_ASAP7_75t_SL g2768 ( 
.A(n_2380),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2255),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2304),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2312),
.Y(n_2771)
);

CKINVDCx16_ASAP7_75t_R g2772 ( 
.A(n_1973),
.Y(n_2772)
);

INVxp67_ASAP7_75t_SL g2773 ( 
.A(n_1825),
.Y(n_2773)
);

INVxp33_ASAP7_75t_SL g2774 ( 
.A(n_1822),
.Y(n_2774)
);

INVxp67_ASAP7_75t_SL g2775 ( 
.A(n_1825),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2408),
.Y(n_2776)
);

INVxp33_ASAP7_75t_SL g2777 ( 
.A(n_1829),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2437),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2458),
.Y(n_2779)
);

CKINVDCx20_ASAP7_75t_R g2780 ( 
.A(n_1814),
.Y(n_2780)
);

INVxp33_ASAP7_75t_L g2781 ( 
.A(n_2229),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2474),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2504),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2532),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2359),
.B(n_0),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2537),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2552),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2554),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2599),
.Y(n_2789)
);

INVxp33_ASAP7_75t_SL g2790 ( 
.A(n_1860),
.Y(n_2790)
);

CKINVDCx16_ASAP7_75t_R g2791 ( 
.A(n_2160),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2621),
.Y(n_2792)
);

INVxp33_ASAP7_75t_SL g2793 ( 
.A(n_1870),
.Y(n_2793)
);

BUFx3_ASAP7_75t_L g2794 ( 
.A(n_1862),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2637),
.Y(n_2795)
);

HB1xp67_ASAP7_75t_L g2796 ( 
.A(n_1882),
.Y(n_2796)
);

INVxp67_ASAP7_75t_SL g2797 ( 
.A(n_1825),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2642),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_1899),
.Y(n_2799)
);

CKINVDCx16_ASAP7_75t_R g2800 ( 
.A(n_2160),
.Y(n_2800)
);

CKINVDCx5p33_ASAP7_75t_R g2801 ( 
.A(n_1898),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2018),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2376),
.Y(n_2803)
);

INVxp67_ASAP7_75t_L g2804 ( 
.A(n_2212),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2399),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2440),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2491),
.Y(n_2807)
);

INVxp67_ASAP7_75t_SL g2808 ( 
.A(n_1838),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2607),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_1838),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_1856),
.Y(n_2811)
);

CKINVDCx5p33_ASAP7_75t_R g2812 ( 
.A(n_1909),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_1856),
.Y(n_2813)
);

HB1xp67_ASAP7_75t_L g2814 ( 
.A(n_1943),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_1856),
.Y(n_2815)
);

INVxp33_ASAP7_75t_SL g2816 ( 
.A(n_2016),
.Y(n_2816)
);

CKINVDCx5p33_ASAP7_75t_R g2817 ( 
.A(n_2026),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_1920),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_1920),
.Y(n_2819)
);

BUFx2_ASAP7_75t_L g2820 ( 
.A(n_2032),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2036),
.Y(n_2821)
);

BUFx6f_ASAP7_75t_L g2822 ( 
.A(n_2036),
.Y(n_2822)
);

CKINVDCx5p33_ASAP7_75t_R g2823 ( 
.A(n_2040),
.Y(n_2823)
);

INVx1_ASAP7_75t_SL g2824 ( 
.A(n_2180),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2054),
.Y(n_2825)
);

CKINVDCx20_ASAP7_75t_R g2826 ( 
.A(n_1818),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2054),
.Y(n_2827)
);

HB1xp67_ASAP7_75t_L g2828 ( 
.A(n_2049),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2054),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2055),
.Y(n_2830)
);

INVxp33_ASAP7_75t_SL g2831 ( 
.A(n_2064),
.Y(n_2831)
);

CKINVDCx5p33_ASAP7_75t_R g2832 ( 
.A(n_2075),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2055),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2055),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2059),
.Y(n_2835)
);

CKINVDCx16_ASAP7_75t_R g2836 ( 
.A(n_2212),
.Y(n_2836)
);

INVxp67_ASAP7_75t_SL g2837 ( 
.A(n_2059),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2059),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2095),
.Y(n_2839)
);

BUFx6f_ASAP7_75t_L g2840 ( 
.A(n_2095),
.Y(n_2840)
);

CKINVDCx5p33_ASAP7_75t_R g2841 ( 
.A(n_2090),
.Y(n_2841)
);

INVxp67_ASAP7_75t_L g2842 ( 
.A(n_2224),
.Y(n_2842)
);

CKINVDCx5p33_ASAP7_75t_R g2843 ( 
.A(n_2103),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2095),
.Y(n_2844)
);

INVxp67_ASAP7_75t_SL g2845 ( 
.A(n_2096),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2096),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2096),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2178),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2178),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2178),
.Y(n_2850)
);

INVx1_ASAP7_75t_SL g2851 ( 
.A(n_2560),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2184),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2184),
.Y(n_2853)
);

INVx1_ASAP7_75t_SL g2854 ( 
.A(n_2367),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2190),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2190),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2192),
.Y(n_2857)
);

INVxp67_ASAP7_75t_L g2858 ( 
.A(n_2224),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2192),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2211),
.Y(n_2860)
);

INVxp67_ASAP7_75t_L g2861 ( 
.A(n_2449),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2211),
.Y(n_2862)
);

INVxp67_ASAP7_75t_SL g2863 ( 
.A(n_2211),
.Y(n_2863)
);

INVxp67_ASAP7_75t_SL g2864 ( 
.A(n_2256),
.Y(n_2864)
);

CKINVDCx20_ASAP7_75t_R g2865 ( 
.A(n_1840),
.Y(n_2865)
);

INVxp33_ASAP7_75t_SL g2866 ( 
.A(n_2109),
.Y(n_2866)
);

HB1xp67_ASAP7_75t_L g2867 ( 
.A(n_2129),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2256),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2256),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2289),
.Y(n_2870)
);

CKINVDCx20_ASAP7_75t_R g2871 ( 
.A(n_1886),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2289),
.Y(n_2872)
);

INVxp33_ASAP7_75t_SL g2873 ( 
.A(n_2130),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2813),
.Y(n_2874)
);

NOR2x1_ASAP7_75t_L g2875 ( 
.A(n_2667),
.B(n_2058),
.Y(n_2875)
);

AND2x6_ASAP7_75t_L g2876 ( 
.A(n_2690),
.B(n_2081),
.Y(n_2876)
);

NOR2xp33_ASAP7_75t_L g2877 ( 
.A(n_2754),
.B(n_2194),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2819),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2666),
.B(n_2289),
.Y(n_2879)
);

AND2x2_ASAP7_75t_L g2880 ( 
.A(n_2693),
.B(n_2669),
.Y(n_2880)
);

NAND2xp33_ASAP7_75t_L g2881 ( 
.A(n_2704),
.B(n_2710),
.Y(n_2881)
);

OA21x2_ASAP7_75t_L g2882 ( 
.A1(n_2668),
.A2(n_1799),
.B(n_1833),
.Y(n_2882)
);

HB1xp67_ASAP7_75t_L g2883 ( 
.A(n_2718),
.Y(n_2883)
);

AND2x4_ASAP7_75t_L g2884 ( 
.A(n_2678),
.B(n_2168),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2773),
.Y(n_2885)
);

AND2x4_ASAP7_75t_L g2886 ( 
.A(n_2756),
.B(n_2245),
.Y(n_2886)
);

INVx2_ASAP7_75t_SL g2887 ( 
.A(n_2753),
.Y(n_2887)
);

AND2x2_ASAP7_75t_L g2888 ( 
.A(n_2768),
.B(n_2260),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_SL g2889 ( 
.A(n_2711),
.B(n_2320),
.Y(n_2889)
);

OAI22x1_ASAP7_75t_SL g2890 ( 
.A1(n_2759),
.A2(n_1998),
.B1(n_2122),
.B2(n_1863),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2775),
.Y(n_2891)
);

INVx3_ASAP7_75t_L g2892 ( 
.A(n_2672),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2825),
.Y(n_2893)
);

INVx2_ASAP7_75t_L g2894 ( 
.A(n_2860),
.Y(n_2894)
);

BUFx6f_ASAP7_75t_L g2895 ( 
.A(n_2672),
.Y(n_2895)
);

OA21x2_ASAP7_75t_L g2896 ( 
.A1(n_2670),
.A2(n_2000),
.B(n_1865),
.Y(n_2896)
);

BUFx6f_ASAP7_75t_L g2897 ( 
.A(n_2822),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2862),
.Y(n_2898)
);

INVxp67_ASAP7_75t_L g2899 ( 
.A(n_2767),
.Y(n_2899)
);

CKINVDCx20_ASAP7_75t_R g2900 ( 
.A(n_2780),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2797),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2808),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2837),
.Y(n_2903)
);

BUFx6f_ASAP7_75t_L g2904 ( 
.A(n_2822),
.Y(n_2904)
);

NOR2xp33_ASAP7_75t_L g2905 ( 
.A(n_2774),
.B(n_1905),
.Y(n_2905)
);

BUFx3_ASAP7_75t_L g2906 ( 
.A(n_2706),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2822),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2845),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2682),
.B(n_2320),
.Y(n_2909)
);

OAI22xp5_ASAP7_75t_L g2910 ( 
.A1(n_2699),
.A2(n_2146),
.B1(n_2150),
.B2(n_2147),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2863),
.Y(n_2911)
);

OA21x2_ASAP7_75t_L g2912 ( 
.A1(n_2675),
.A2(n_2044),
.B(n_2025),
.Y(n_2912)
);

BUFx3_ASAP7_75t_L g2913 ( 
.A(n_2719),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2729),
.B(n_2730),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2864),
.Y(n_2915)
);

BUFx6f_ASAP7_75t_L g2916 ( 
.A(n_2840),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2734),
.Y(n_2917)
);

BUFx6f_ASAP7_75t_L g2918 ( 
.A(n_2840),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2677),
.Y(n_2919)
);

BUFx6f_ASAP7_75t_L g2920 ( 
.A(n_2747),
.Y(n_2920)
);

OAI21x1_ASAP7_75t_L g2921 ( 
.A1(n_2679),
.A2(n_2050),
.B(n_2048),
.Y(n_2921)
);

BUFx3_ASAP7_75t_L g2922 ( 
.A(n_2794),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2680),
.Y(n_2923)
);

NOR2x1_ASAP7_75t_L g2924 ( 
.A(n_2681),
.B(n_2276),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2683),
.Y(n_2925)
);

BUFx2_ASAP7_75t_L g2926 ( 
.A(n_2723),
.Y(n_2926)
);

AOI22xp5_ASAP7_75t_L g2927 ( 
.A1(n_2752),
.A2(n_2173),
.B1(n_2195),
.B2(n_2171),
.Y(n_2927)
);

CKINVDCx6p67_ASAP7_75t_R g2928 ( 
.A(n_2694),
.Y(n_2928)
);

OAI21x1_ASAP7_75t_L g2929 ( 
.A1(n_2687),
.A2(n_2070),
.B(n_2060),
.Y(n_2929)
);

CKINVDCx5p33_ASAP7_75t_R g2930 ( 
.A(n_2676),
.Y(n_2930)
);

AND2x2_ASAP7_75t_L g2931 ( 
.A(n_2820),
.B(n_2301),
.Y(n_2931)
);

OA21x2_ASAP7_75t_L g2932 ( 
.A1(n_2688),
.A2(n_2092),
.B(n_2072),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2810),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2811),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2815),
.Y(n_2935)
);

AND2x2_ASAP7_75t_L g2936 ( 
.A(n_2796),
.B(n_2382),
.Y(n_2936)
);

CKINVDCx20_ASAP7_75t_R g2937 ( 
.A(n_2826),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2818),
.Y(n_2938)
);

BUFx2_ASAP7_75t_L g2939 ( 
.A(n_2727),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2821),
.Y(n_2940)
);

NOR2xp33_ASAP7_75t_L g2941 ( 
.A(n_2777),
.B(n_1960),
.Y(n_2941)
);

AOI22xp5_ASAP7_75t_L g2942 ( 
.A1(n_2673),
.A2(n_2216),
.B1(n_2217),
.B2(n_2197),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2827),
.Y(n_2943)
);

OAI22xp5_ASAP7_75t_L g2944 ( 
.A1(n_2674),
.A2(n_2247),
.B1(n_2252),
.B2(n_2230),
.Y(n_2944)
);

BUFx3_ASAP7_75t_L g2945 ( 
.A(n_2829),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2830),
.Y(n_2946)
);

BUFx6f_ASAP7_75t_L g2947 ( 
.A(n_2763),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2833),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2834),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2835),
.Y(n_2950)
);

INVxp67_ASAP7_75t_L g2951 ( 
.A(n_2814),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2838),
.Y(n_2952)
);

AND2x4_ASAP7_75t_L g2953 ( 
.A(n_2685),
.B(n_2386),
.Y(n_2953)
);

AOI22xp5_ASAP7_75t_L g2954 ( 
.A1(n_2720),
.A2(n_2270),
.B1(n_2281),
.B2(n_2263),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2839),
.Y(n_2955)
);

OA21x2_ASAP7_75t_L g2956 ( 
.A1(n_2691),
.A2(n_2121),
.B(n_2120),
.Y(n_2956)
);

AND2x4_ASAP7_75t_L g2957 ( 
.A(n_2697),
.B(n_2728),
.Y(n_2957)
);

INVx5_ASAP7_75t_L g2958 ( 
.A(n_2772),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2844),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2846),
.Y(n_2960)
);

OA21x2_ASAP7_75t_L g2961 ( 
.A1(n_2692),
.A2(n_2164),
.B(n_2132),
.Y(n_2961)
);

INVx3_ASAP7_75t_L g2962 ( 
.A(n_2806),
.Y(n_2962)
);

INVx6_ASAP7_75t_L g2963 ( 
.A(n_2791),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2847),
.Y(n_2964)
);

BUFx8_ASAP7_75t_L g2965 ( 
.A(n_2746),
.Y(n_2965)
);

BUFx6f_ASAP7_75t_L g2966 ( 
.A(n_2765),
.Y(n_2966)
);

BUFx2_ASAP7_75t_L g2967 ( 
.A(n_2736),
.Y(n_2967)
);

BUFx6f_ASAP7_75t_L g2968 ( 
.A(n_2782),
.Y(n_2968)
);

BUFx6f_ASAP7_75t_L g2969 ( 
.A(n_2789),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2848),
.Y(n_2970)
);

AOI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2724),
.A2(n_2291),
.B1(n_2292),
.B2(n_2283),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2849),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2850),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2852),
.Y(n_2974)
);

BUFx6f_ASAP7_75t_L g2975 ( 
.A(n_2795),
.Y(n_2975)
);

AND2x4_ASAP7_75t_L g2976 ( 
.A(n_2828),
.B(n_2423),
.Y(n_2976)
);

INVx2_ASAP7_75t_SL g2977 ( 
.A(n_2801),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2853),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2867),
.B(n_2429),
.Y(n_2979)
);

AND2x2_ASAP7_75t_L g2980 ( 
.A(n_2748),
.B(n_2435),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2855),
.Y(n_2981)
);

INVx5_ASAP7_75t_L g2982 ( 
.A(n_2800),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2812),
.B(n_2330),
.Y(n_2983)
);

AND2x4_ASAP7_75t_L g2984 ( 
.A(n_2804),
.B(n_2454),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2817),
.B(n_2339),
.Y(n_2985)
);

AND2x6_ASAP7_75t_L g2986 ( 
.A(n_2726),
.B(n_2136),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2856),
.Y(n_2987)
);

CKINVDCx5p33_ASAP7_75t_R g2988 ( 
.A(n_2684),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2857),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2859),
.Y(n_2990)
);

INVx3_ASAP7_75t_L g2991 ( 
.A(n_2868),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2869),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2870),
.Y(n_2993)
);

OA21x2_ASAP7_75t_L g2994 ( 
.A1(n_2695),
.A2(n_2272),
.B(n_2251),
.Y(n_2994)
);

AOI22x1_ASAP7_75t_SL g2995 ( 
.A1(n_2737),
.A2(n_2343),
.B1(n_2424),
.B2(n_2202),
.Y(n_2995)
);

HB1xp67_ASAP7_75t_L g2996 ( 
.A(n_2732),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2872),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2698),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2700),
.Y(n_2999)
);

BUFx6f_ASAP7_75t_L g3000 ( 
.A(n_2738),
.Y(n_3000)
);

INVx3_ASAP7_75t_L g3001 ( 
.A(n_2739),
.Y(n_3001)
);

CKINVDCx16_ASAP7_75t_R g3002 ( 
.A(n_2665),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2701),
.Y(n_3003)
);

XNOR2xp5_ASAP7_75t_L g3004 ( 
.A(n_2865),
.B(n_2493),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2703),
.Y(n_3005)
);

OA21x2_ASAP7_75t_L g3006 ( 
.A1(n_2705),
.A2(n_2708),
.B(n_2707),
.Y(n_3006)
);

AND2x4_ASAP7_75t_L g3007 ( 
.A(n_2842),
.B(n_2482),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2709),
.Y(n_3008)
);

INVx3_ASAP7_75t_L g3009 ( 
.A(n_2741),
.Y(n_3009)
);

AND2x4_ASAP7_75t_L g3010 ( 
.A(n_2858),
.B(n_2643),
.Y(n_3010)
);

BUFx3_ASAP7_75t_L g3011 ( 
.A(n_2712),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2713),
.Y(n_3012)
);

NOR2xp33_ASAP7_75t_L g3013 ( 
.A(n_2790),
.B(n_2277),
.Y(n_3013)
);

AOI22xp5_ASAP7_75t_SL g3014 ( 
.A1(n_2760),
.A2(n_2568),
.B1(n_2590),
.B2(n_2544),
.Y(n_3014)
);

INVx3_ASAP7_75t_L g3015 ( 
.A(n_2742),
.Y(n_3015)
);

BUFx6f_ASAP7_75t_L g3016 ( 
.A(n_2744),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2714),
.Y(n_3017)
);

AND2x2_ASAP7_75t_L g3018 ( 
.A(n_2823),
.B(n_2449),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2715),
.Y(n_3019)
);

CKINVDCx20_ASAP7_75t_R g3020 ( 
.A(n_2871),
.Y(n_3020)
);

BUFx6f_ASAP7_75t_L g3021 ( 
.A(n_2745),
.Y(n_3021)
);

INVx5_ASAP7_75t_L g3022 ( 
.A(n_2836),
.Y(n_3022)
);

CKINVDCx6p67_ASAP7_75t_R g3023 ( 
.A(n_2689),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2716),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2717),
.Y(n_3025)
);

INVx6_ASAP7_75t_L g3026 ( 
.A(n_2793),
.Y(n_3026)
);

OA21x2_ASAP7_75t_L g3027 ( 
.A1(n_2721),
.A2(n_2294),
.B(n_2278),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2722),
.Y(n_3028)
);

INVx4_ASAP7_75t_L g3029 ( 
.A(n_2832),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2725),
.Y(n_3030)
);

AND2x4_ASAP7_75t_L g3031 ( 
.A(n_2861),
.B(n_1820),
.Y(n_3031)
);

BUFx6f_ASAP7_75t_L g3032 ( 
.A(n_2749),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_2731),
.Y(n_3033)
);

NAND2xp33_ASAP7_75t_L g3034 ( 
.A(n_2841),
.B(n_2300),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2733),
.Y(n_3035)
);

AND2x4_ASAP7_75t_L g3036 ( 
.A(n_2843),
.B(n_1877),
.Y(n_3036)
);

NAND2xp33_ASAP7_75t_L g3037 ( 
.A(n_2702),
.B(n_2323),
.Y(n_3037)
);

BUFx6f_ASAP7_75t_L g3038 ( 
.A(n_2750),
.Y(n_3038)
);

BUFx6f_ASAP7_75t_L g3039 ( 
.A(n_2751),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2755),
.Y(n_3040)
);

BUFx2_ASAP7_75t_L g3041 ( 
.A(n_2735),
.Y(n_3041)
);

AND2x6_ASAP7_75t_L g3042 ( 
.A(n_2785),
.B(n_2495),
.Y(n_3042)
);

BUFx6f_ASAP7_75t_L g3043 ( 
.A(n_2758),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_2781),
.B(n_2583),
.Y(n_3044)
);

CKINVDCx5p33_ASAP7_75t_R g3045 ( 
.A(n_2696),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2761),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2816),
.B(n_2339),
.Y(n_3047)
);

CKINVDCx5p33_ASAP7_75t_R g3048 ( 
.A(n_2930),
.Y(n_3048)
);

CKINVDCx5p33_ASAP7_75t_R g3049 ( 
.A(n_2988),
.Y(n_3049)
);

BUFx2_ASAP7_75t_L g3050 ( 
.A(n_2986),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_3040),
.Y(n_3051)
);

CKINVDCx5p33_ASAP7_75t_R g3052 ( 
.A(n_3045),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_2907),
.Y(n_3053)
);

CKINVDCx5p33_ASAP7_75t_R g3054 ( 
.A(n_2900),
.Y(n_3054)
);

CKINVDCx5p33_ASAP7_75t_R g3055 ( 
.A(n_2937),
.Y(n_3055)
);

INVxp67_ASAP7_75t_L g3056 ( 
.A(n_2877),
.Y(n_3056)
);

CKINVDCx5p33_ASAP7_75t_R g3057 ( 
.A(n_3020),
.Y(n_3057)
);

CKINVDCx5p33_ASAP7_75t_R g3058 ( 
.A(n_2928),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_3046),
.Y(n_3059)
);

BUFx6f_ASAP7_75t_SL g3060 ( 
.A(n_2986),
.Y(n_3060)
);

CKINVDCx5p33_ASAP7_75t_R g3061 ( 
.A(n_3023),
.Y(n_3061)
);

CKINVDCx5p33_ASAP7_75t_R g3062 ( 
.A(n_3002),
.Y(n_3062)
);

CKINVDCx5p33_ASAP7_75t_R g3063 ( 
.A(n_3029),
.Y(n_3063)
);

CKINVDCx5p33_ASAP7_75t_R g3064 ( 
.A(n_2887),
.Y(n_3064)
);

CKINVDCx20_ASAP7_75t_R g3065 ( 
.A(n_2926),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2874),
.Y(n_3066)
);

CKINVDCx5p33_ASAP7_75t_R g3067 ( 
.A(n_2977),
.Y(n_3067)
);

CKINVDCx5p33_ASAP7_75t_R g3068 ( 
.A(n_2939),
.Y(n_3068)
);

CKINVDCx5p33_ASAP7_75t_R g3069 ( 
.A(n_2967),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_3000),
.Y(n_3070)
);

CKINVDCx5p33_ASAP7_75t_R g3071 ( 
.A(n_3004),
.Y(n_3071)
);

AND2x2_ASAP7_75t_L g3072 ( 
.A(n_3044),
.B(n_2740),
.Y(n_3072)
);

CKINVDCx5p33_ASAP7_75t_R g3073 ( 
.A(n_3026),
.Y(n_3073)
);

HB1xp67_ASAP7_75t_L g3074 ( 
.A(n_2980),
.Y(n_3074)
);

CKINVDCx5p33_ASAP7_75t_R g3075 ( 
.A(n_2958),
.Y(n_3075)
);

CKINVDCx5p33_ASAP7_75t_R g3076 ( 
.A(n_2982),
.Y(n_3076)
);

CKINVDCx5p33_ASAP7_75t_R g3077 ( 
.A(n_3022),
.Y(n_3077)
);

CKINVDCx16_ASAP7_75t_R g3078 ( 
.A(n_2883),
.Y(n_3078)
);

CKINVDCx5p33_ASAP7_75t_R g3079 ( 
.A(n_2963),
.Y(n_3079)
);

CKINVDCx5p33_ASAP7_75t_R g3080 ( 
.A(n_2996),
.Y(n_3080)
);

CKINVDCx5p33_ASAP7_75t_R g3081 ( 
.A(n_2922),
.Y(n_3081)
);

CKINVDCx5p33_ASAP7_75t_R g3082 ( 
.A(n_2906),
.Y(n_3082)
);

BUFx6f_ASAP7_75t_L g3083 ( 
.A(n_2897),
.Y(n_3083)
);

CKINVDCx5p33_ASAP7_75t_R g3084 ( 
.A(n_2913),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2878),
.Y(n_3085)
);

OAI22xp5_ASAP7_75t_SL g3086 ( 
.A1(n_2942),
.A2(n_1921),
.B1(n_1927),
.B2(n_1893),
.Y(n_3086)
);

CKINVDCx5p33_ASAP7_75t_R g3087 ( 
.A(n_2899),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_2893),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_3016),
.Y(n_3089)
);

INVx2_ASAP7_75t_L g3090 ( 
.A(n_2894),
.Y(n_3090)
);

CKINVDCx5p33_ASAP7_75t_R g3091 ( 
.A(n_2983),
.Y(n_3091)
);

NOR2xp33_ASAP7_75t_R g3092 ( 
.A(n_2881),
.B(n_2671),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2985),
.B(n_2831),
.Y(n_3093)
);

NOR2xp33_ASAP7_75t_R g3094 ( 
.A(n_3034),
.B(n_2824),
.Y(n_3094)
);

NOR2xp33_ASAP7_75t_R g3095 ( 
.A(n_3037),
.B(n_2851),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2898),
.Y(n_3096)
);

CKINVDCx5p33_ASAP7_75t_R g3097 ( 
.A(n_2965),
.Y(n_3097)
);

AND2x2_ASAP7_75t_L g3098 ( 
.A(n_2880),
.B(n_2686),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_2931),
.B(n_2888),
.Y(n_3099)
);

CKINVDCx20_ASAP7_75t_R g3100 ( 
.A(n_2951),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_3021),
.Y(n_3101)
);

INVx2_ASAP7_75t_L g3102 ( 
.A(n_2920),
.Y(n_3102)
);

CKINVDCx5p33_ASAP7_75t_R g3103 ( 
.A(n_3018),
.Y(n_3103)
);

NOR2xp33_ASAP7_75t_R g3104 ( 
.A(n_2917),
.B(n_2854),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_3032),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_3038),
.Y(n_3106)
);

CKINVDCx5p33_ASAP7_75t_R g3107 ( 
.A(n_3047),
.Y(n_3107)
);

NOR2xp33_ASAP7_75t_L g3108 ( 
.A(n_2914),
.B(n_2866),
.Y(n_3108)
);

INVxp67_ASAP7_75t_SL g3109 ( 
.A(n_2909),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_3039),
.Y(n_3110)
);

INVx11_ASAP7_75t_L g3111 ( 
.A(n_2876),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_SL g3112 ( 
.A(n_3036),
.B(n_2873),
.Y(n_3112)
);

CKINVDCx5p33_ASAP7_75t_R g3113 ( 
.A(n_2890),
.Y(n_3113)
);

NOR2xp33_ASAP7_75t_R g3114 ( 
.A(n_2885),
.B(n_1965),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_3011),
.B(n_2762),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_3043),
.Y(n_3116)
);

BUFx6f_ASAP7_75t_L g3117 ( 
.A(n_2904),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2923),
.Y(n_3118)
);

CKINVDCx5p33_ASAP7_75t_R g3119 ( 
.A(n_2995),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2947),
.Y(n_3120)
);

BUFx10_ASAP7_75t_L g3121 ( 
.A(n_2957),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2998),
.Y(n_3122)
);

NOR2xp33_ASAP7_75t_SL g3123 ( 
.A(n_2876),
.B(n_2531),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2999),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_3005),
.Y(n_3125)
);

CKINVDCx5p33_ASAP7_75t_R g3126 ( 
.A(n_2954),
.Y(n_3126)
);

CKINVDCx5p33_ASAP7_75t_R g3127 ( 
.A(n_2971),
.Y(n_3127)
);

CKINVDCx5p33_ASAP7_75t_R g3128 ( 
.A(n_3042),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_2966),
.Y(n_3129)
);

CKINVDCx5p33_ASAP7_75t_R g3130 ( 
.A(n_2910),
.Y(n_3130)
);

INVxp67_ASAP7_75t_L g3131 ( 
.A(n_2905),
.Y(n_3131)
);

CKINVDCx5p33_ASAP7_75t_R g3132 ( 
.A(n_2941),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_3017),
.Y(n_3133)
);

CKINVDCx20_ASAP7_75t_R g3134 ( 
.A(n_3014),
.Y(n_3134)
);

CKINVDCx5p33_ASAP7_75t_R g3135 ( 
.A(n_3013),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_3019),
.Y(n_3136)
);

NOR2xp33_ASAP7_75t_R g3137 ( 
.A(n_2891),
.B(n_1967),
.Y(n_3137)
);

NOR2xp33_ASAP7_75t_L g3138 ( 
.A(n_2889),
.B(n_2743),
.Y(n_3138)
);

CKINVDCx5p33_ASAP7_75t_R g3139 ( 
.A(n_2944),
.Y(n_3139)
);

CKINVDCx6p67_ASAP7_75t_R g3140 ( 
.A(n_2984),
.Y(n_3140)
);

CKINVDCx5p33_ASAP7_75t_R g3141 ( 
.A(n_2886),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_3024),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_3028),
.Y(n_3143)
);

INVxp67_ASAP7_75t_L g3144 ( 
.A(n_2936),
.Y(n_3144)
);

CKINVDCx5p33_ASAP7_75t_R g3145 ( 
.A(n_2927),
.Y(n_3145)
);

CKINVDCx20_ASAP7_75t_R g3146 ( 
.A(n_2979),
.Y(n_3146)
);

BUFx2_ASAP7_75t_L g3147 ( 
.A(n_3007),
.Y(n_3147)
);

CKINVDCx5p33_ASAP7_75t_R g3148 ( 
.A(n_2901),
.Y(n_3148)
);

CKINVDCx20_ASAP7_75t_R g3149 ( 
.A(n_2879),
.Y(n_3149)
);

CKINVDCx5p33_ASAP7_75t_R g3150 ( 
.A(n_2902),
.Y(n_3150)
);

CKINVDCx16_ASAP7_75t_R g3151 ( 
.A(n_2976),
.Y(n_3151)
);

BUFx3_ASAP7_75t_L g3152 ( 
.A(n_2882),
.Y(n_3152)
);

CKINVDCx5p33_ASAP7_75t_R g3153 ( 
.A(n_2903),
.Y(n_3153)
);

INVx2_ASAP7_75t_L g3154 ( 
.A(n_2968),
.Y(n_3154)
);

NOR2xp33_ASAP7_75t_R g3155 ( 
.A(n_2908),
.B(n_1970),
.Y(n_3155)
);

CKINVDCx5p33_ASAP7_75t_R g3156 ( 
.A(n_2911),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_3030),
.Y(n_3157)
);

CKINVDCx5p33_ASAP7_75t_R g3158 ( 
.A(n_2915),
.Y(n_3158)
);

BUFx6f_ASAP7_75t_L g3159 ( 
.A(n_2916),
.Y(n_3159)
);

CKINVDCx5p33_ASAP7_75t_R g3160 ( 
.A(n_2884),
.Y(n_3160)
);

CKINVDCx20_ASAP7_75t_R g3161 ( 
.A(n_2945),
.Y(n_3161)
);

CKINVDCx5p33_ASAP7_75t_R g3162 ( 
.A(n_2953),
.Y(n_3162)
);

INVx2_ASAP7_75t_L g3163 ( 
.A(n_2969),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2919),
.Y(n_3164)
);

CKINVDCx5p33_ASAP7_75t_R g3165 ( 
.A(n_3010),
.Y(n_3165)
);

CKINVDCx5p33_ASAP7_75t_R g3166 ( 
.A(n_3031),
.Y(n_3166)
);

NOR2xp67_ASAP7_75t_L g3167 ( 
.A(n_3001),
.B(n_2764),
.Y(n_3167)
);

CKINVDCx5p33_ASAP7_75t_R g3168 ( 
.A(n_2975),
.Y(n_3168)
);

BUFx10_ASAP7_75t_L g3169 ( 
.A(n_2935),
.Y(n_3169)
);

NOR2xp33_ASAP7_75t_R g3170 ( 
.A(n_3009),
.B(n_2008),
.Y(n_3170)
);

NOR2xp33_ASAP7_75t_R g3171 ( 
.A(n_3015),
.B(n_2030),
.Y(n_3171)
);

INVx3_ASAP7_75t_L g3172 ( 
.A(n_2925),
.Y(n_3172)
);

CKINVDCx5p33_ASAP7_75t_R g3173 ( 
.A(n_3003),
.Y(n_3173)
);

INVx4_ASAP7_75t_L g3174 ( 
.A(n_3006),
.Y(n_3174)
);

HB1xp67_ASAP7_75t_L g3175 ( 
.A(n_2892),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_3008),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_3012),
.Y(n_3177)
);

CKINVDCx5p33_ASAP7_75t_R g3178 ( 
.A(n_3025),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2933),
.Y(n_3179)
);

CKINVDCx5p33_ASAP7_75t_R g3180 ( 
.A(n_3033),
.Y(n_3180)
);

CKINVDCx5p33_ASAP7_75t_R g3181 ( 
.A(n_3035),
.Y(n_3181)
);

CKINVDCx5p33_ASAP7_75t_R g3182 ( 
.A(n_2918),
.Y(n_3182)
);

INVx2_ASAP7_75t_L g3183 ( 
.A(n_2934),
.Y(n_3183)
);

CKINVDCx5p33_ASAP7_75t_R g3184 ( 
.A(n_2895),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_SL g3185 ( 
.A(n_2875),
.B(n_2757),
.Y(n_3185)
);

INVx2_ASAP7_75t_SL g3186 ( 
.A(n_2924),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2896),
.Y(n_3187)
);

CKINVDCx5p33_ASAP7_75t_R g3188 ( 
.A(n_2962),
.Y(n_3188)
);

CKINVDCx5p33_ASAP7_75t_R g3189 ( 
.A(n_2943),
.Y(n_3189)
);

BUFx2_ASAP7_75t_L g3190 ( 
.A(n_2912),
.Y(n_3190)
);

CKINVDCx5p33_ASAP7_75t_R g3191 ( 
.A(n_2949),
.Y(n_3191)
);

CKINVDCx5p33_ASAP7_75t_R g3192 ( 
.A(n_2950),
.Y(n_3192)
);

CKINVDCx5p33_ASAP7_75t_R g3193 ( 
.A(n_2955),
.Y(n_3193)
);

HB1xp67_ASAP7_75t_L g3194 ( 
.A(n_2932),
.Y(n_3194)
);

CKINVDCx20_ASAP7_75t_R g3195 ( 
.A(n_2956),
.Y(n_3195)
);

CKINVDCx5p33_ASAP7_75t_R g3196 ( 
.A(n_2964),
.Y(n_3196)
);

CKINVDCx5p33_ASAP7_75t_R g3197 ( 
.A(n_2978),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2961),
.Y(n_3198)
);

CKINVDCx5p33_ASAP7_75t_R g3199 ( 
.A(n_2987),
.Y(n_3199)
);

CKINVDCx5p33_ASAP7_75t_R g3200 ( 
.A(n_2990),
.Y(n_3200)
);

CKINVDCx5p33_ASAP7_75t_R g3201 ( 
.A(n_2993),
.Y(n_3201)
);

CKINVDCx5p33_ASAP7_75t_R g3202 ( 
.A(n_2997),
.Y(n_3202)
);

CKINVDCx5p33_ASAP7_75t_R g3203 ( 
.A(n_2938),
.Y(n_3203)
);

CKINVDCx20_ASAP7_75t_R g3204 ( 
.A(n_2994),
.Y(n_3204)
);

HB1xp67_ASAP7_75t_L g3205 ( 
.A(n_3027),
.Y(n_3205)
);

CKINVDCx16_ASAP7_75t_R g3206 ( 
.A(n_2940),
.Y(n_3206)
);

INVx3_ASAP7_75t_L g3207 ( 
.A(n_2921),
.Y(n_3207)
);

INVx3_ASAP7_75t_L g3208 ( 
.A(n_2929),
.Y(n_3208)
);

CKINVDCx5p33_ASAP7_75t_R g3209 ( 
.A(n_2946),
.Y(n_3209)
);

NOR2xp33_ASAP7_75t_R g3210 ( 
.A(n_2991),
.B(n_2043),
.Y(n_3210)
);

CKINVDCx5p33_ASAP7_75t_R g3211 ( 
.A(n_2948),
.Y(n_3211)
);

CKINVDCx5p33_ASAP7_75t_R g3212 ( 
.A(n_2952),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_2959),
.Y(n_3213)
);

INVx3_ASAP7_75t_L g3214 ( 
.A(n_2992),
.Y(n_3214)
);

NAND2xp33_ASAP7_75t_L g3215 ( 
.A(n_2960),
.B(n_2356),
.Y(n_3215)
);

CKINVDCx20_ASAP7_75t_R g3216 ( 
.A(n_2970),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_2972),
.Y(n_3217)
);

CKINVDCx20_ASAP7_75t_R g3218 ( 
.A(n_2973),
.Y(n_3218)
);

NOR2xp33_ASAP7_75t_R g3219 ( 
.A(n_2974),
.B(n_2084),
.Y(n_3219)
);

HB1xp67_ASAP7_75t_L g3220 ( 
.A(n_2981),
.Y(n_3220)
);

BUFx6f_ASAP7_75t_L g3221 ( 
.A(n_2989),
.Y(n_3221)
);

NOR2xp33_ASAP7_75t_SL g3222 ( 
.A(n_3002),
.B(n_2089),
.Y(n_3222)
);

CKINVDCx5p33_ASAP7_75t_R g3223 ( 
.A(n_2930),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_2907),
.Y(n_3224)
);

CKINVDCx5p33_ASAP7_75t_R g3225 ( 
.A(n_2930),
.Y(n_3225)
);

BUFx6f_ASAP7_75t_SL g3226 ( 
.A(n_2986),
.Y(n_3226)
);

CKINVDCx5p33_ASAP7_75t_R g3227 ( 
.A(n_2930),
.Y(n_3227)
);

NAND2xp33_ASAP7_75t_R g3228 ( 
.A(n_3041),
.B(n_2370),
.Y(n_3228)
);

CKINVDCx20_ASAP7_75t_R g3229 ( 
.A(n_2900),
.Y(n_3229)
);

NOR2x1p5_ASAP7_75t_L g3230 ( 
.A(n_3023),
.B(n_2393),
.Y(n_3230)
);

NOR2xp33_ASAP7_75t_R g3231 ( 
.A(n_2930),
.B(n_2126),
.Y(n_3231)
);

BUFx8_ASAP7_75t_SL g3232 ( 
.A(n_3229),
.Y(n_3232)
);

NOR2xp33_ASAP7_75t_L g3233 ( 
.A(n_3056),
.B(n_1806),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3051),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_SL g3235 ( 
.A(n_3099),
.B(n_2356),
.Y(n_3235)
);

OR2x6_ASAP7_75t_L g3236 ( 
.A(n_3050),
.B(n_1937),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_3109),
.B(n_2356),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_3059),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3066),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_3085),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_3131),
.B(n_1828),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_3088),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_3090),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_3091),
.B(n_2363),
.Y(n_3244)
);

INVx4_ASAP7_75t_L g3245 ( 
.A(n_3168),
.Y(n_3245)
);

INVx3_ASAP7_75t_L g3246 ( 
.A(n_3083),
.Y(n_3246)
);

INVxp33_ASAP7_75t_L g3247 ( 
.A(n_3231),
.Y(n_3247)
);

INVx2_ASAP7_75t_L g3248 ( 
.A(n_3096),
.Y(n_3248)
);

AND2x6_ASAP7_75t_L g3249 ( 
.A(n_3187),
.B(n_2406),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3118),
.Y(n_3250)
);

INVx4_ASAP7_75t_L g3251 ( 
.A(n_3182),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_3122),
.Y(n_3252)
);

BUFx6f_ASAP7_75t_L g3253 ( 
.A(n_3083),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_3108),
.B(n_2406),
.Y(n_3254)
);

INVx3_ASAP7_75t_L g3255 ( 
.A(n_3083),
.Y(n_3255)
);

BUFx3_ASAP7_75t_L g3256 ( 
.A(n_3161),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3124),
.Y(n_3257)
);

INVx2_ASAP7_75t_L g3258 ( 
.A(n_3172),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3125),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_3194),
.B(n_2409),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_3205),
.B(n_2409),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_3107),
.B(n_2409),
.Y(n_3262)
);

NOR2xp33_ASAP7_75t_L g3263 ( 
.A(n_3132),
.B(n_1864),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_3172),
.Y(n_3264)
);

BUFx4f_ASAP7_75t_L g3265 ( 
.A(n_3140),
.Y(n_3265)
);

BUFx10_ASAP7_75t_L g3266 ( 
.A(n_3060),
.Y(n_3266)
);

INVx5_ASAP7_75t_L g3267 ( 
.A(n_3121),
.Y(n_3267)
);

INVx2_ASAP7_75t_L g3268 ( 
.A(n_3179),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3133),
.Y(n_3269)
);

INVx4_ASAP7_75t_L g3270 ( 
.A(n_3184),
.Y(n_3270)
);

INVx5_ASAP7_75t_L g3271 ( 
.A(n_3121),
.Y(n_3271)
);

CKINVDCx5p33_ASAP7_75t_R g3272 ( 
.A(n_3048),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3136),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3142),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_SL g3275 ( 
.A(n_3148),
.B(n_2419),
.Y(n_3275)
);

OR2x2_ASAP7_75t_SL g3276 ( 
.A(n_3151),
.B(n_2302),
.Y(n_3276)
);

AND2x2_ASAP7_75t_SL g3277 ( 
.A(n_3123),
.B(n_2419),
.Y(n_3277)
);

CKINVDCx5p33_ASAP7_75t_R g3278 ( 
.A(n_3049),
.Y(n_3278)
);

CKINVDCx5p33_ASAP7_75t_R g3279 ( 
.A(n_3052),
.Y(n_3279)
);

BUFx6f_ASAP7_75t_L g3280 ( 
.A(n_3117),
.Y(n_3280)
);

INVx2_ASAP7_75t_SL g3281 ( 
.A(n_3188),
.Y(n_3281)
);

INVx2_ASAP7_75t_SL g3282 ( 
.A(n_3098),
.Y(n_3282)
);

AOI22xp5_ASAP7_75t_L g3283 ( 
.A1(n_3195),
.A2(n_2172),
.B1(n_2199),
.B2(n_2185),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_3183),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3143),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_3157),
.B(n_2468),
.Y(n_3286)
);

CKINVDCx5p33_ASAP7_75t_R g3287 ( 
.A(n_3223),
.Y(n_3287)
);

AOI22xp5_ASAP7_75t_L g3288 ( 
.A1(n_3204),
.A2(n_2200),
.B1(n_2220),
.B2(n_2219),
.Y(n_3288)
);

OR2x6_ASAP7_75t_SL g3289 ( 
.A(n_3135),
.B(n_2394),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_3220),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_3152),
.B(n_2468),
.Y(n_3291)
);

CKINVDCx5p33_ASAP7_75t_R g3292 ( 
.A(n_3225),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_3144),
.B(n_2766),
.Y(n_3293)
);

INVx1_ASAP7_75t_SL g3294 ( 
.A(n_3146),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3213),
.Y(n_3295)
);

NOR2x1p5_ASAP7_75t_L g3296 ( 
.A(n_3079),
.B(n_2402),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_3164),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3217),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_SL g3299 ( 
.A(n_3150),
.B(n_2477),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_3072),
.B(n_2769),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3214),
.Y(n_3301)
);

INVx5_ASAP7_75t_L g3302 ( 
.A(n_3117),
.Y(n_3302)
);

BUFx6f_ASAP7_75t_L g3303 ( 
.A(n_3117),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_SL g3304 ( 
.A(n_3153),
.B(n_2477),
.Y(n_3304)
);

OAI21xp33_ASAP7_75t_L g3305 ( 
.A1(n_3138),
.A2(n_3158),
.B(n_3156),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3214),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3175),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_3053),
.Y(n_3308)
);

AND2x4_ASAP7_75t_L g3309 ( 
.A(n_3120),
.B(n_2770),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3190),
.B(n_2477),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_SL g3311 ( 
.A(n_3093),
.B(n_2514),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3174),
.B(n_2514),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_SL g3313 ( 
.A(n_3064),
.B(n_2514),
.Y(n_3313)
);

BUFx3_ASAP7_75t_L g3314 ( 
.A(n_3159),
.Y(n_3314)
);

INVx2_ASAP7_75t_SL g3315 ( 
.A(n_3169),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3224),
.Y(n_3316)
);

OR2x6_ASAP7_75t_L g3317 ( 
.A(n_3147),
.B(n_2227),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3176),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3177),
.Y(n_3319)
);

AND2x2_ASAP7_75t_L g3320 ( 
.A(n_3103),
.B(n_2771),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_3067),
.B(n_3104),
.Y(n_3321)
);

NOR2xp33_ASAP7_75t_L g3322 ( 
.A(n_3149),
.B(n_1866),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3198),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_SL g3324 ( 
.A(n_3094),
.B(n_2525),
.Y(n_3324)
);

CKINVDCx20_ASAP7_75t_R g3325 ( 
.A(n_3054),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_3173),
.B(n_2525),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_3115),
.Y(n_3327)
);

INVx4_ASAP7_75t_L g3328 ( 
.A(n_3073),
.Y(n_3328)
);

AOI22xp33_ASAP7_75t_L g3329 ( 
.A1(n_3207),
.A2(n_2569),
.B1(n_2612),
.B2(n_2548),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_SL g3330 ( 
.A(n_3095),
.B(n_2548),
.Y(n_3330)
);

OR2x2_ASAP7_75t_L g3331 ( 
.A(n_3206),
.B(n_2657),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3167),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_3189),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_3221),
.Y(n_3334)
);

NOR2xp33_ASAP7_75t_L g3335 ( 
.A(n_3178),
.B(n_1887),
.Y(n_3335)
);

CKINVDCx16_ASAP7_75t_R g3336 ( 
.A(n_3222),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_3180),
.B(n_2569),
.Y(n_3337)
);

OR2x2_ASAP7_75t_L g3338 ( 
.A(n_3078),
.B(n_1983),
.Y(n_3338)
);

HB1xp67_ASAP7_75t_SL g3339 ( 
.A(n_3062),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3191),
.Y(n_3340)
);

AOI22xp33_ASAP7_75t_L g3341 ( 
.A1(n_3207),
.A2(n_2612),
.B1(n_2569),
.B2(n_1989),
.Y(n_3341)
);

BUFx6f_ASAP7_75t_L g3342 ( 
.A(n_3159),
.Y(n_3342)
);

BUFx6f_ASAP7_75t_L g3343 ( 
.A(n_3159),
.Y(n_3343)
);

INVx3_ASAP7_75t_L g3344 ( 
.A(n_3129),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_SL g3345 ( 
.A(n_3181),
.B(n_2612),
.Y(n_3345)
);

INVx4_ASAP7_75t_L g3346 ( 
.A(n_3081),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3192),
.Y(n_3347)
);

INVxp33_ASAP7_75t_L g3348 ( 
.A(n_3170),
.Y(n_3348)
);

AOI22xp5_ASAP7_75t_L g3349 ( 
.A1(n_3126),
.A2(n_2315),
.B1(n_2331),
.B2(n_2327),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3193),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_3221),
.Y(n_3351)
);

BUFx8_ASAP7_75t_SL g3352 ( 
.A(n_3061),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3196),
.Y(n_3353)
);

NOR2xp33_ASAP7_75t_L g3354 ( 
.A(n_3087),
.B(n_1985),
.Y(n_3354)
);

HB1xp67_ASAP7_75t_L g3355 ( 
.A(n_3210),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3197),
.Y(n_3356)
);

OAI22xp5_ASAP7_75t_L g3357 ( 
.A1(n_3130),
.A2(n_3139),
.B1(n_3127),
.B2(n_3145),
.Y(n_3357)
);

NOR2xp33_ASAP7_75t_L g3358 ( 
.A(n_3203),
.B(n_1994),
.Y(n_3358)
);

BUFx3_ASAP7_75t_L g3359 ( 
.A(n_3082),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3199),
.Y(n_3360)
);

NOR2xp33_ASAP7_75t_L g3361 ( 
.A(n_3209),
.B(n_2015),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3200),
.Y(n_3362)
);

INVx3_ASAP7_75t_L g3363 ( 
.A(n_3154),
.Y(n_3363)
);

BUFx6f_ASAP7_75t_L g3364 ( 
.A(n_3221),
.Y(n_3364)
);

OR2x2_ASAP7_75t_L g3365 ( 
.A(n_3112),
.B(n_3166),
.Y(n_3365)
);

OR2x2_ASAP7_75t_L g3366 ( 
.A(n_3071),
.B(n_2061),
.Y(n_3366)
);

AND2x2_ASAP7_75t_L g3367 ( 
.A(n_3171),
.B(n_2776),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3201),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_3211),
.B(n_2105),
.Y(n_3369)
);

OR2x6_ASAP7_75t_L g3370 ( 
.A(n_3230),
.B(n_1956),
.Y(n_3370)
);

CKINVDCx5p33_ASAP7_75t_R g3371 ( 
.A(n_3227),
.Y(n_3371)
);

BUFx6f_ASAP7_75t_L g3372 ( 
.A(n_3163),
.Y(n_3372)
);

INVx6_ASAP7_75t_L g3373 ( 
.A(n_3169),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3202),
.Y(n_3374)
);

AND2x2_ASAP7_75t_L g3375 ( 
.A(n_3114),
.B(n_2778),
.Y(n_3375)
);

NOR2xp33_ASAP7_75t_L g3376 ( 
.A(n_3212),
.B(n_2113),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_3186),
.B(n_3063),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3208),
.B(n_2234),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_SL g3379 ( 
.A(n_3141),
.B(n_1802),
.Y(n_3379)
);

INVx1_ASAP7_75t_SL g3380 ( 
.A(n_3137),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3185),
.B(n_2290),
.Y(n_3381)
);

INVx2_ASAP7_75t_SL g3382 ( 
.A(n_3219),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_3070),
.Y(n_3383)
);

AND2x2_ASAP7_75t_L g3384 ( 
.A(n_3155),
.B(n_2779),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_SL g3385 ( 
.A(n_3160),
.B(n_1805),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3089),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_3101),
.Y(n_3387)
);

OR2x2_ASAP7_75t_L g3388 ( 
.A(n_3086),
.B(n_2235),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_SL g3389 ( 
.A(n_3092),
.B(n_1808),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_SL g3390 ( 
.A(n_3128),
.B(n_1811),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3105),
.Y(n_3391)
);

INVx3_ASAP7_75t_L g3392 ( 
.A(n_3106),
.Y(n_3392)
);

INVxp67_ASAP7_75t_L g3393 ( 
.A(n_3228),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3110),
.Y(n_3394)
);

INVx4_ASAP7_75t_L g3395 ( 
.A(n_3084),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3116),
.Y(n_3396)
);

BUFx3_ASAP7_75t_L g3397 ( 
.A(n_3065),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3216),
.Y(n_3398)
);

NAND3xp33_ASAP7_75t_L g3399 ( 
.A(n_3080),
.B(n_2433),
.C(n_2407),
.Y(n_3399)
);

INVx5_ASAP7_75t_L g3400 ( 
.A(n_3111),
.Y(n_3400)
);

NOR2xp33_ASAP7_75t_L g3401 ( 
.A(n_3162),
.B(n_2274),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_3218),
.Y(n_3402)
);

CKINVDCx16_ASAP7_75t_R g3403 ( 
.A(n_3060),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3215),
.Y(n_3404)
);

AND2x4_ASAP7_75t_L g3405 ( 
.A(n_3165),
.B(n_2783),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_3226),
.Y(n_3406)
);

NOR2x1p5_ASAP7_75t_L g3407 ( 
.A(n_3075),
.B(n_2439),
.Y(n_3407)
);

BUFx3_ASAP7_75t_L g3408 ( 
.A(n_3055),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_3226),
.Y(n_3409)
);

OR2x6_ASAP7_75t_L g3410 ( 
.A(n_3057),
.B(n_2540),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3100),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_3076),
.B(n_2542),
.Y(n_3412)
);

AND2x2_ASAP7_75t_L g3413 ( 
.A(n_3068),
.B(n_2784),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_3077),
.Y(n_3414)
);

NOR2xp33_ASAP7_75t_SL g3415 ( 
.A(n_3058),
.B(n_3069),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3134),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3119),
.B(n_2593),
.Y(n_3417)
);

AND2x6_ASAP7_75t_L g3418 ( 
.A(n_3113),
.B(n_1800),
.Y(n_3418)
);

AND2x2_ASAP7_75t_L g3419 ( 
.A(n_3097),
.B(n_2786),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_3066),
.Y(n_3420)
);

INVx4_ASAP7_75t_L g3421 ( 
.A(n_3168),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3051),
.Y(n_3422)
);

AND2x2_ASAP7_75t_L g3423 ( 
.A(n_3098),
.B(n_2787),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3051),
.Y(n_3424)
);

BUFx3_ASAP7_75t_L g3425 ( 
.A(n_3168),
.Y(n_3425)
);

BUFx8_ASAP7_75t_SL g3426 ( 
.A(n_3229),
.Y(n_3426)
);

NOR2xp33_ASAP7_75t_L g3427 ( 
.A(n_3056),
.B(n_2472),
.Y(n_3427)
);

BUFx6f_ASAP7_75t_L g3428 ( 
.A(n_3083),
.Y(n_3428)
);

INVx2_ASAP7_75t_L g3429 ( 
.A(n_3066),
.Y(n_3429)
);

NAND2x1p5_ASAP7_75t_L g3430 ( 
.A(n_3099),
.B(n_2788),
.Y(n_3430)
);

NAND3xp33_ASAP7_75t_L g3431 ( 
.A(n_3056),
.B(n_2484),
.C(n_2448),
.Y(n_3431)
);

AND2x2_ASAP7_75t_L g3432 ( 
.A(n_3098),
.B(n_2792),
.Y(n_3432)
);

BUFx6f_ASAP7_75t_L g3433 ( 
.A(n_3083),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_SL g3434 ( 
.A(n_3099),
.B(n_1813),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3109),
.B(n_2798),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_SL g3436 ( 
.A(n_3099),
.B(n_1817),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3109),
.B(n_1821),
.Y(n_3437)
);

AND2x6_ASAP7_75t_L g3438 ( 
.A(n_3187),
.B(n_1803),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3051),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3051),
.Y(n_3440)
);

AND2x4_ASAP7_75t_L g3441 ( 
.A(n_3102),
.B(n_2799),
.Y(n_3441)
);

INVx2_ASAP7_75t_L g3442 ( 
.A(n_3066),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3051),
.Y(n_3443)
);

INVx2_ASAP7_75t_SL g3444 ( 
.A(n_3074),
.Y(n_3444)
);

INVx3_ASAP7_75t_L g3445 ( 
.A(n_3083),
.Y(n_3445)
);

OR2x6_ASAP7_75t_L g3446 ( 
.A(n_3050),
.B(n_1804),
.Y(n_3446)
);

CKINVDCx5p33_ASAP7_75t_R g3447 ( 
.A(n_3048),
.Y(n_3447)
);

CKINVDCx5p33_ASAP7_75t_R g3448 ( 
.A(n_3048),
.Y(n_3448)
);

AND2x4_ASAP7_75t_L g3449 ( 
.A(n_3102),
.B(n_2802),
.Y(n_3449)
);

CKINVDCx20_ASAP7_75t_R g3450 ( 
.A(n_3229),
.Y(n_3450)
);

BUFx8_ASAP7_75t_SL g3451 ( 
.A(n_3229),
.Y(n_3451)
);

INVx2_ASAP7_75t_L g3452 ( 
.A(n_3066),
.Y(n_3452)
);

INVx2_ASAP7_75t_SL g3453 ( 
.A(n_3074),
.Y(n_3453)
);

INVxp67_ASAP7_75t_L g3454 ( 
.A(n_3138),
.Y(n_3454)
);

INVx4_ASAP7_75t_L g3455 ( 
.A(n_3168),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_SL g3456 ( 
.A(n_3099),
.B(n_1823),
.Y(n_3456)
);

NOR2xp33_ASAP7_75t_L g3457 ( 
.A(n_3056),
.B(n_2589),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_3109),
.B(n_1824),
.Y(n_3458)
);

INVx4_ASAP7_75t_L g3459 ( 
.A(n_3168),
.Y(n_3459)
);

AND2x2_ASAP7_75t_L g3460 ( 
.A(n_3098),
.B(n_1924),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3109),
.B(n_1826),
.Y(n_3461)
);

OR2x6_ASAP7_75t_L g3462 ( 
.A(n_3050),
.B(n_1809),
.Y(n_3462)
);

CKINVDCx20_ASAP7_75t_R g3463 ( 
.A(n_3229),
.Y(n_3463)
);

INVx3_ASAP7_75t_L g3464 ( 
.A(n_3083),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3066),
.Y(n_3465)
);

INVx2_ASAP7_75t_L g3466 ( 
.A(n_3066),
.Y(n_3466)
);

AND2x4_ASAP7_75t_L g3467 ( 
.A(n_3102),
.B(n_2803),
.Y(n_3467)
);

AND2x2_ASAP7_75t_L g3468 ( 
.A(n_3098),
.B(n_1924),
.Y(n_3468)
);

BUFx6f_ASAP7_75t_L g3469 ( 
.A(n_3083),
.Y(n_3469)
);

NOR2xp33_ASAP7_75t_L g3470 ( 
.A(n_3056),
.B(n_2651),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_L g3471 ( 
.A(n_3056),
.B(n_2655),
.Y(n_3471)
);

CKINVDCx20_ASAP7_75t_R g3472 ( 
.A(n_3229),
.Y(n_3472)
);

OAI22xp5_ASAP7_75t_L g3473 ( 
.A1(n_3195),
.A2(n_1839),
.B1(n_1844),
.B2(n_1831),
.Y(n_3473)
);

OR2x6_ASAP7_75t_L g3474 ( 
.A(n_3050),
.B(n_1810),
.Y(n_3474)
);

NOR2xp33_ASAP7_75t_L g3475 ( 
.A(n_3056),
.B(n_2499),
.Y(n_3475)
);

NOR2xp33_ASAP7_75t_L g3476 ( 
.A(n_3056),
.B(n_2508),
.Y(n_3476)
);

INVx4_ASAP7_75t_SL g3477 ( 
.A(n_3060),
.Y(n_3477)
);

BUFx3_ASAP7_75t_L g3478 ( 
.A(n_3168),
.Y(n_3478)
);

OR2x2_ASAP7_75t_L g3479 ( 
.A(n_3098),
.B(n_2512),
.Y(n_3479)
);

BUFx6f_ASAP7_75t_L g3480 ( 
.A(n_3083),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_SL g3481 ( 
.A(n_3305),
.B(n_2365),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3234),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3454),
.B(n_1845),
.Y(n_3483)
);

AOI22xp33_ASAP7_75t_L g3484 ( 
.A1(n_3438),
.A2(n_3277),
.B1(n_3378),
.B2(n_3323),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3435),
.B(n_1849),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3254),
.B(n_1853),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3233),
.B(n_1854),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3238),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3427),
.B(n_1857),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3250),
.Y(n_3490)
);

AND2x6_ASAP7_75t_SL g3491 ( 
.A(n_3410),
.B(n_1827),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3252),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3240),
.Y(n_3493)
);

AOI22xp5_ASAP7_75t_L g3494 ( 
.A1(n_3393),
.A2(n_2428),
.B1(n_2441),
.B2(n_2397),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3257),
.Y(n_3495)
);

O2A1O1Ixp33_ASAP7_75t_L g3496 ( 
.A1(n_3235),
.A2(n_1832),
.B(n_1834),
.C(n_1830),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3259),
.Y(n_3497)
);

INVx8_ASAP7_75t_L g3498 ( 
.A(n_3302),
.Y(n_3498)
);

AOI22xp33_ASAP7_75t_L g3499 ( 
.A1(n_3438),
.A2(n_2465),
.B1(n_2466),
.B2(n_2453),
.Y(n_3499)
);

AOI22xp33_ASAP7_75t_L g3500 ( 
.A1(n_3438),
.A2(n_2516),
.B1(n_2517),
.B2(n_2507),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3457),
.B(n_1859),
.Y(n_3501)
);

AND2x6_ASAP7_75t_L g3502 ( 
.A(n_3300),
.B(n_1835),
.Y(n_3502)
);

NOR2xp33_ASAP7_75t_L g3503 ( 
.A(n_3263),
.B(n_2526),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3470),
.B(n_1868),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_SL g3505 ( 
.A(n_3321),
.B(n_2527),
.Y(n_3505)
);

BUFx3_ASAP7_75t_L g3506 ( 
.A(n_3425),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3471),
.B(n_1869),
.Y(n_3507)
);

NOR2xp33_ASAP7_75t_L g3508 ( 
.A(n_3358),
.B(n_2541),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3241),
.B(n_1872),
.Y(n_3509)
);

AOI221xp5_ASAP7_75t_L g3510 ( 
.A1(n_3361),
.A2(n_2535),
.B1(n_2539),
.B2(n_2521),
.C(n_2519),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3437),
.B(n_1874),
.Y(n_3511)
);

INVx2_ASAP7_75t_SL g3512 ( 
.A(n_3405),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3248),
.Y(n_3513)
);

AND2x2_ASAP7_75t_L g3514 ( 
.A(n_3320),
.B(n_2038),
.Y(n_3514)
);

INVx2_ASAP7_75t_SL g3515 ( 
.A(n_3423),
.Y(n_3515)
);

NOR2xp33_ASAP7_75t_L g3516 ( 
.A(n_3369),
.B(n_2547),
.Y(n_3516)
);

BUFx3_ASAP7_75t_L g3517 ( 
.A(n_3478),
.Y(n_3517)
);

NOR2xp33_ASAP7_75t_L g3518 ( 
.A(n_3376),
.B(n_2549),
.Y(n_3518)
);

INVx2_ASAP7_75t_SL g3519 ( 
.A(n_3432),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_3420),
.Y(n_3520)
);

NOR2xp33_ASAP7_75t_L g3521 ( 
.A(n_3354),
.B(n_2570),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3458),
.B(n_1879),
.Y(n_3522)
);

AOI21x1_ASAP7_75t_L g3523 ( 
.A1(n_3312),
.A2(n_2807),
.B(n_2805),
.Y(n_3523)
);

AOI22xp33_ASAP7_75t_L g3524 ( 
.A1(n_3269),
.A2(n_2608),
.B1(n_2617),
.B2(n_2600),
.Y(n_3524)
);

NOR2xp33_ASAP7_75t_L g3525 ( 
.A(n_3380),
.B(n_2641),
.Y(n_3525)
);

AOI22xp5_ASAP7_75t_L g3526 ( 
.A1(n_3282),
.A2(n_1888),
.B1(n_1889),
.B2(n_1883),
.Y(n_3526)
);

OAI221xp5_ASAP7_75t_L g3527 ( 
.A1(n_3475),
.A2(n_1841),
.B1(n_1842),
.B2(n_1837),
.C(n_1836),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3461),
.B(n_1891),
.Y(n_3528)
);

AOI22xp33_ASAP7_75t_L g3529 ( 
.A1(n_3273),
.A2(n_2345),
.B1(n_2352),
.B2(n_2344),
.Y(n_3529)
);

NOR3xp33_ASAP7_75t_L g3530 ( 
.A(n_3322),
.B(n_1895),
.C(n_1894),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3274),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_3429),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_3244),
.B(n_1896),
.Y(n_3533)
);

NOR2xp33_ASAP7_75t_L g3534 ( 
.A(n_3335),
.B(n_1902),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_SL g3535 ( 
.A(n_3333),
.B(n_1903),
.Y(n_3535)
);

AOI221xp5_ASAP7_75t_L g3536 ( 
.A1(n_3476),
.A2(n_2587),
.B1(n_2591),
.B2(n_2573),
.C(n_2567),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3285),
.Y(n_3537)
);

NAND2xp5_ASAP7_75t_SL g3538 ( 
.A(n_3340),
.B(n_3347),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3301),
.B(n_1908),
.Y(n_3539)
);

INVx4_ASAP7_75t_L g3540 ( 
.A(n_3267),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_SL g3541 ( 
.A(n_3350),
.B(n_1913),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3306),
.B(n_1916),
.Y(n_3542)
);

AND2x6_ASAP7_75t_SL g3543 ( 
.A(n_3410),
.B(n_1846),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3262),
.B(n_1918),
.Y(n_3544)
);

INVx2_ASAP7_75t_L g3545 ( 
.A(n_3442),
.Y(n_3545)
);

OAI22x1_ASAP7_75t_L g3546 ( 
.A1(n_3349),
.A2(n_2632),
.B1(n_2635),
.B2(n_2610),
.Y(n_3546)
);

NOR2xp33_ASAP7_75t_L g3547 ( 
.A(n_3348),
.B(n_1919),
.Y(n_3547)
);

AOI22xp33_ASAP7_75t_L g3548 ( 
.A1(n_3422),
.A2(n_2374),
.B1(n_2405),
.B2(n_2362),
.Y(n_3548)
);

NOR2xp33_ASAP7_75t_L g3549 ( 
.A(n_3366),
.B(n_1923),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3424),
.Y(n_3550)
);

INVx3_ASAP7_75t_L g3551 ( 
.A(n_3253),
.Y(n_3551)
);

INVx2_ASAP7_75t_L g3552 ( 
.A(n_3452),
.Y(n_3552)
);

A2O1A1Ixp33_ASAP7_75t_L g3553 ( 
.A1(n_3439),
.A2(n_1848),
.B(n_1850),
.C(n_1847),
.Y(n_3553)
);

INVx2_ASAP7_75t_L g3554 ( 
.A(n_3465),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_SL g3555 ( 
.A(n_3353),
.B(n_1925),
.Y(n_3555)
);

AND2x6_ASAP7_75t_L g3556 ( 
.A(n_3367),
.B(n_1852),
.Y(n_3556)
);

AND2x4_ASAP7_75t_L g3557 ( 
.A(n_3267),
.B(n_2809),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3375),
.B(n_3384),
.Y(n_3558)
);

OR2x2_ASAP7_75t_L g3559 ( 
.A(n_3331),
.B(n_2649),
.Y(n_3559)
);

OR2x2_ASAP7_75t_L g3560 ( 
.A(n_3479),
.B(n_2650),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3466),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3440),
.B(n_1926),
.Y(n_3562)
);

NAND2xp33_ASAP7_75t_L g3563 ( 
.A(n_3355),
.B(n_1928),
.Y(n_3563)
);

AOI22xp5_ASAP7_75t_L g3564 ( 
.A1(n_3443),
.A2(n_1931),
.B1(n_1933),
.B2(n_1929),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3293),
.B(n_1936),
.Y(n_3565)
);

INVx2_ASAP7_75t_L g3566 ( 
.A(n_3268),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3239),
.Y(n_3567)
);

AOI22xp5_ASAP7_75t_L g3568 ( 
.A1(n_3295),
.A2(n_1941),
.B1(n_1942),
.B2(n_1939),
.Y(n_3568)
);

INVx4_ASAP7_75t_L g3569 ( 
.A(n_3271),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3334),
.B(n_1945),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3242),
.Y(n_3571)
);

AOI22xp5_ASAP7_75t_L g3572 ( 
.A1(n_3298),
.A2(n_1948),
.B1(n_1949),
.B2(n_1946),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_SL g3573 ( 
.A(n_3356),
.B(n_1950),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3351),
.B(n_1952),
.Y(n_3574)
);

NOR3xp33_ASAP7_75t_L g3575 ( 
.A(n_3357),
.B(n_1955),
.C(n_1954),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3310),
.B(n_1957),
.Y(n_3576)
);

BUFx3_ASAP7_75t_L g3577 ( 
.A(n_3256),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3237),
.B(n_1962),
.Y(n_3578)
);

O2A1O1Ixp33_ASAP7_75t_L g3579 ( 
.A1(n_3260),
.A2(n_1858),
.B(n_1867),
.C(n_1855),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3460),
.B(n_3468),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3261),
.B(n_3284),
.Y(n_3581)
);

NOR2xp33_ASAP7_75t_L g3582 ( 
.A(n_3401),
.B(n_3247),
.Y(n_3582)
);

BUFx6f_ASAP7_75t_L g3583 ( 
.A(n_3253),
.Y(n_3583)
);

O2A1O1Ixp5_ASAP7_75t_L g3584 ( 
.A1(n_3291),
.A2(n_2447),
.B(n_2479),
.C(n_2438),
.Y(n_3584)
);

NOR2xp33_ASAP7_75t_L g3585 ( 
.A(n_3382),
.B(n_1964),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3243),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3332),
.B(n_1966),
.Y(n_3587)
);

A2O1A1Ixp33_ASAP7_75t_L g3588 ( 
.A1(n_3431),
.A2(n_1873),
.B(n_1875),
.C(n_1871),
.Y(n_3588)
);

A2O1A1Ixp33_ASAP7_75t_L g3589 ( 
.A1(n_3318),
.A2(n_1880),
.B(n_1881),
.C(n_1878),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3326),
.B(n_1968),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3319),
.Y(n_3591)
);

INVx2_ASAP7_75t_SL g3592 ( 
.A(n_3413),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3337),
.B(n_3297),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3430),
.B(n_1971),
.Y(n_3594)
);

NOR2xp33_ASAP7_75t_L g3595 ( 
.A(n_3283),
.B(n_1972),
.Y(n_3595)
);

BUFx6f_ASAP7_75t_SL g3596 ( 
.A(n_3266),
.Y(n_3596)
);

INVx2_ASAP7_75t_L g3597 ( 
.A(n_3308),
.Y(n_3597)
);

INVx3_ASAP7_75t_L g3598 ( 
.A(n_3280),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3316),
.B(n_1974),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3258),
.B(n_3264),
.Y(n_3600)
);

NOR2xp33_ASAP7_75t_L g3601 ( 
.A(n_3288),
.B(n_1975),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3377),
.B(n_1977),
.Y(n_3602)
);

INVx3_ASAP7_75t_L g3603 ( 
.A(n_3280),
.Y(n_3603)
);

AOI22xp33_ASAP7_75t_L g3604 ( 
.A1(n_3388),
.A2(n_2571),
.B1(n_2576),
.B2(n_2497),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3441),
.Y(n_3605)
);

AOI22xp33_ASAP7_75t_L g3606 ( 
.A1(n_3341),
.A2(n_2586),
.B1(n_2613),
.B2(n_2579),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3329),
.B(n_3360),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_SL g3608 ( 
.A(n_3362),
.B(n_1979),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3449),
.Y(n_3609)
);

AND2x2_ASAP7_75t_L g3610 ( 
.A(n_3368),
.B(n_2078),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3467),
.Y(n_3611)
);

OR2x6_ASAP7_75t_L g3612 ( 
.A(n_3245),
.B(n_1884),
.Y(n_3612)
);

INVx2_ASAP7_75t_SL g3613 ( 
.A(n_3303),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3374),
.B(n_1984),
.Y(n_3614)
);

OAI22xp5_ASAP7_75t_L g3615 ( 
.A1(n_3290),
.A2(n_3444),
.B1(n_3453),
.B2(n_3315),
.Y(n_3615)
);

NAND3xp33_ASAP7_75t_L g3616 ( 
.A(n_3473),
.B(n_1988),
.C(n_1986),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_L g3617 ( 
.A(n_3249),
.B(n_3286),
.Y(n_3617)
);

AOI22xp33_ASAP7_75t_L g3618 ( 
.A1(n_3434),
.A2(n_2660),
.B1(n_2639),
.B2(n_1890),
.Y(n_3618)
);

NOR2x1p5_ASAP7_75t_L g3619 ( 
.A(n_3421),
.B(n_1990),
.Y(n_3619)
);

AOI22xp5_ASAP7_75t_L g3620 ( 
.A1(n_3436),
.A2(n_2001),
.B1(n_2002),
.B2(n_1996),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_SL g3621 ( 
.A(n_3281),
.B(n_2003),
.Y(n_3621)
);

INVx2_ASAP7_75t_L g3622 ( 
.A(n_3309),
.Y(n_3622)
);

INVx8_ASAP7_75t_L g3623 ( 
.A(n_3302),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3383),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3381),
.B(n_2004),
.Y(n_3625)
);

INVx1_ASAP7_75t_SL g3626 ( 
.A(n_3294),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3386),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3391),
.Y(n_3628)
);

NOR2xp33_ASAP7_75t_L g3629 ( 
.A(n_3338),
.B(n_2006),
.Y(n_3629)
);

INVx4_ASAP7_75t_L g3630 ( 
.A(n_3271),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_SL g3631 ( 
.A(n_3336),
.B(n_3346),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3456),
.B(n_2007),
.Y(n_3632)
);

CKINVDCx20_ASAP7_75t_R g3633 ( 
.A(n_3232),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3311),
.B(n_2009),
.Y(n_3634)
);

BUFx3_ASAP7_75t_L g3635 ( 
.A(n_3450),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_SL g3636 ( 
.A(n_3395),
.B(n_2010),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_SL g3637 ( 
.A(n_3359),
.B(n_2011),
.Y(n_3637)
);

INVxp33_ASAP7_75t_L g3638 ( 
.A(n_3419),
.Y(n_3638)
);

INVx2_ASAP7_75t_L g3639 ( 
.A(n_3387),
.Y(n_3639)
);

AND2x6_ASAP7_75t_L g3640 ( 
.A(n_3409),
.B(n_1900),
.Y(n_3640)
);

NOR2xp33_ASAP7_75t_L g3641 ( 
.A(n_3390),
.B(n_2012),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_SL g3642 ( 
.A(n_3455),
.B(n_2013),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3394),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3392),
.Y(n_3644)
);

AOI22xp33_ASAP7_75t_SL g3645 ( 
.A1(n_3415),
.A2(n_2091),
.B1(n_2198),
.B2(n_2078),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3396),
.Y(n_3646)
);

INVx2_ASAP7_75t_L g3647 ( 
.A(n_3344),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_3404),
.B(n_2014),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_3373),
.B(n_2091),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_SL g3650 ( 
.A(n_3459),
.B(n_2017),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3307),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3324),
.B(n_2019),
.Y(n_3652)
);

AND2x2_ASAP7_75t_L g3653 ( 
.A(n_3251),
.B(n_2198),
.Y(n_3653)
);

BUFx3_ASAP7_75t_L g3654 ( 
.A(n_3463),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3363),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3372),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_SL g3657 ( 
.A(n_3272),
.B(n_3278),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3330),
.B(n_2020),
.Y(n_3658)
);

AND2x2_ASAP7_75t_L g3659 ( 
.A(n_3270),
.B(n_2213),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_SL g3660 ( 
.A(n_3279),
.B(n_3287),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_3246),
.Y(n_3661)
);

INVx4_ASAP7_75t_L g3662 ( 
.A(n_3292),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3389),
.B(n_2021),
.Y(n_3663)
);

AND2x2_ASAP7_75t_L g3664 ( 
.A(n_3371),
.B(n_2213),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3255),
.Y(n_3665)
);

NOR2xp33_ASAP7_75t_L g3666 ( 
.A(n_3365),
.B(n_2022),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3445),
.Y(n_3667)
);

INVx2_ASAP7_75t_L g3668 ( 
.A(n_3464),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3345),
.B(n_3275),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3299),
.B(n_2023),
.Y(n_3670)
);

BUFx3_ASAP7_75t_L g3671 ( 
.A(n_3472),
.Y(n_3671)
);

AOI22xp5_ASAP7_75t_L g3672 ( 
.A1(n_3399),
.A2(n_2029),
.B1(n_2031),
.B2(n_2027),
.Y(n_3672)
);

A2O1A1Ixp33_ASAP7_75t_L g3673 ( 
.A1(n_3304),
.A2(n_1907),
.B(n_1910),
.C(n_1901),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3314),
.Y(n_3674)
);

AOI22xp5_ASAP7_75t_L g3675 ( 
.A1(n_3379),
.A2(n_2034),
.B1(n_2035),
.B2(n_2033),
.Y(n_3675)
);

AOI22xp5_ASAP7_75t_L g3676 ( 
.A1(n_3385),
.A2(n_3236),
.B1(n_3317),
.B2(n_3446),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_SL g3677 ( 
.A(n_3447),
.B(n_2037),
.Y(n_3677)
);

O2A1O1Ixp5_ASAP7_75t_L g3678 ( 
.A1(n_3313),
.A2(n_1912),
.B(n_1915),
.C(n_1911),
.Y(n_3678)
);

AND2x2_ASAP7_75t_L g3679 ( 
.A(n_3448),
.B(n_2232),
.Y(n_3679)
);

AND2x2_ASAP7_75t_L g3680 ( 
.A(n_3402),
.B(n_2232),
.Y(n_3680)
);

NAND2xp33_ASAP7_75t_L g3681 ( 
.A(n_3400),
.B(n_2042),
.Y(n_3681)
);

INVx2_ASAP7_75t_SL g3682 ( 
.A(n_3342),
.Y(n_3682)
);

INVx2_ASAP7_75t_L g3683 ( 
.A(n_3480),
.Y(n_3683)
);

INVx2_ASAP7_75t_SL g3684 ( 
.A(n_3342),
.Y(n_3684)
);

NOR2xp33_ASAP7_75t_L g3685 ( 
.A(n_3411),
.B(n_3328),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3412),
.B(n_2045),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3343),
.Y(n_3687)
);

AOI22xp5_ASAP7_75t_L g3688 ( 
.A1(n_3317),
.A2(n_2052),
.B1(n_2053),
.B2(n_2046),
.Y(n_3688)
);

INVx2_ASAP7_75t_L g3689 ( 
.A(n_3428),
.Y(n_3689)
);

NOR2xp33_ASAP7_75t_L g3690 ( 
.A(n_3398),
.B(n_3417),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3433),
.Y(n_3691)
);

INVx5_ASAP7_75t_L g3692 ( 
.A(n_3469),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_SL g3693 ( 
.A(n_3400),
.B(n_2062),
.Y(n_3693)
);

AND2x2_ASAP7_75t_L g3694 ( 
.A(n_3408),
.B(n_2237),
.Y(n_3694)
);

INVx2_ASAP7_75t_L g3695 ( 
.A(n_3469),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_L g3696 ( 
.A(n_3397),
.B(n_2063),
.Y(n_3696)
);

INVx4_ASAP7_75t_L g3697 ( 
.A(n_3265),
.Y(n_3697)
);

NOR2xp67_ASAP7_75t_L g3698 ( 
.A(n_3414),
.B(n_2066),
.Y(n_3698)
);

INVx2_ASAP7_75t_L g3699 ( 
.A(n_3276),
.Y(n_3699)
);

AOI22xp5_ASAP7_75t_L g3700 ( 
.A1(n_3446),
.A2(n_2069),
.B1(n_2073),
.B2(n_2068),
.Y(n_3700)
);

INVx2_ASAP7_75t_L g3701 ( 
.A(n_3462),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_3296),
.B(n_2076),
.Y(n_3702)
);

INVx2_ASAP7_75t_L g3703 ( 
.A(n_3462),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3474),
.B(n_2079),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3406),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3407),
.B(n_2085),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_L g3707 ( 
.A(n_3370),
.B(n_2094),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3370),
.B(n_2099),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3418),
.B(n_2100),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3418),
.B(n_2101),
.Y(n_3710)
);

AND2x6_ASAP7_75t_SL g3711 ( 
.A(n_3416),
.B(n_1922),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3477),
.B(n_2104),
.Y(n_3712)
);

NOR3xp33_ASAP7_75t_L g3713 ( 
.A(n_3403),
.B(n_2107),
.C(n_2106),
.Y(n_3713)
);

AOI22xp33_ASAP7_75t_L g3714 ( 
.A1(n_3325),
.A2(n_1932),
.B1(n_1934),
.B2(n_1930),
.Y(n_3714)
);

NOR2xp33_ASAP7_75t_L g3715 ( 
.A(n_3339),
.B(n_2112),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_3289),
.B(n_2115),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_SL g3717 ( 
.A(n_3426),
.B(n_2116),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3451),
.Y(n_3718)
);

INVxp67_ASAP7_75t_SL g3719 ( 
.A(n_3352),
.Y(n_3719)
);

OAI22xp33_ASAP7_75t_L g3720 ( 
.A1(n_3454),
.A2(n_2119),
.B1(n_2124),
.B2(n_2117),
.Y(n_3720)
);

NOR2xp33_ASAP7_75t_L g3721 ( 
.A(n_3454),
.B(n_2125),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_3327),
.B(n_2133),
.Y(n_3722)
);

BUFx6f_ASAP7_75t_SL g3723 ( 
.A(n_3266),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_SL g3724 ( 
.A(n_3305),
.B(n_2134),
.Y(n_3724)
);

AOI21xp5_ASAP7_75t_L g3725 ( 
.A1(n_3312),
.A2(n_1938),
.B(n_1935),
.Y(n_3725)
);

OAI22xp5_ASAP7_75t_L g3726 ( 
.A1(n_3454),
.A2(n_2138),
.B1(n_2143),
.B2(n_2137),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3327),
.B(n_2144),
.Y(n_3727)
);

NOR2xp33_ASAP7_75t_L g3728 ( 
.A(n_3454),
.B(n_2148),
.Y(n_3728)
);

NOR2xp33_ASAP7_75t_L g3729 ( 
.A(n_3454),
.B(n_2149),
.Y(n_3729)
);

BUFx6f_ASAP7_75t_L g3730 ( 
.A(n_3253),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3327),
.B(n_2152),
.Y(n_3731)
);

OAI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_3454),
.A2(n_2154),
.B1(n_2156),
.B2(n_2153),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3327),
.B(n_2159),
.Y(n_3733)
);

NOR2xp33_ASAP7_75t_L g3734 ( 
.A(n_3454),
.B(n_2162),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_SL g3735 ( 
.A(n_3305),
.B(n_2163),
.Y(n_3735)
);

INVx4_ASAP7_75t_L g3736 ( 
.A(n_3425),
.Y(n_3736)
);

NOR2xp33_ASAP7_75t_L g3737 ( 
.A(n_3454),
.B(n_2165),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3234),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_SL g3739 ( 
.A(n_3305),
.B(n_2169),
.Y(n_3739)
);

NOR2xp33_ASAP7_75t_L g3740 ( 
.A(n_3454),
.B(n_2170),
.Y(n_3740)
);

OR2x6_ASAP7_75t_L g3741 ( 
.A(n_3425),
.B(n_1940),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3327),
.B(n_2174),
.Y(n_3742)
);

AOI22xp5_ASAP7_75t_L g3743 ( 
.A1(n_3327),
.A2(n_2176),
.B1(n_2181),
.B2(n_2175),
.Y(n_3743)
);

AOI22xp5_ASAP7_75t_L g3744 ( 
.A1(n_3327),
.A2(n_2183),
.B1(n_2186),
.B2(n_2182),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3240),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3234),
.Y(n_3746)
);

OAI22xp5_ASAP7_75t_L g3747 ( 
.A1(n_3454),
.A2(n_2188),
.B1(n_2189),
.B2(n_2187),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_SL g3748 ( 
.A(n_3305),
.B(n_2191),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3240),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3327),
.B(n_2196),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3327),
.B(n_2201),
.Y(n_3751)
);

BUFx5_ASAP7_75t_L g3752 ( 
.A(n_3323),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_SL g3753 ( 
.A(n_3305),
.B(n_2205),
.Y(n_3753)
);

NOR2xp33_ASAP7_75t_L g3754 ( 
.A(n_3454),
.B(n_2206),
.Y(n_3754)
);

OAI22xp5_ASAP7_75t_L g3755 ( 
.A1(n_3454),
.A2(n_2209),
.B1(n_2210),
.B2(n_2208),
.Y(n_3755)
);

NOR2xp33_ASAP7_75t_L g3756 ( 
.A(n_3454),
.B(n_2214),
.Y(n_3756)
);

AOI22xp5_ASAP7_75t_L g3757 ( 
.A1(n_3327),
.A2(n_2221),
.B1(n_2222),
.B2(n_2218),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3234),
.Y(n_3758)
);

INVxp67_ASAP7_75t_SL g3759 ( 
.A(n_3364),
.Y(n_3759)
);

INVx2_ASAP7_75t_SL g3760 ( 
.A(n_3405),
.Y(n_3760)
);

INVx4_ASAP7_75t_L g3761 ( 
.A(n_3425),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3233),
.B(n_2250),
.Y(n_3762)
);

NOR2xp33_ASAP7_75t_L g3763 ( 
.A(n_3454),
.B(n_2223),
.Y(n_3763)
);

INVx2_ASAP7_75t_L g3764 ( 
.A(n_3240),
.Y(n_3764)
);

NAND2xp33_ASAP7_75t_L g3765 ( 
.A(n_3438),
.B(n_2225),
.Y(n_3765)
);

INVx2_ASAP7_75t_SL g3766 ( 
.A(n_3405),
.Y(n_3766)
);

AOI221xp5_ASAP7_75t_L g3767 ( 
.A1(n_3241),
.A2(n_1969),
.B1(n_1978),
.B2(n_1951),
.C(n_1947),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3240),
.Y(n_3768)
);

OR2x6_ASAP7_75t_L g3769 ( 
.A(n_3736),
.B(n_1980),
.Y(n_3769)
);

AOI21xp5_ASAP7_75t_L g3770 ( 
.A1(n_3581),
.A2(n_1991),
.B(n_1987),
.Y(n_3770)
);

NAND2xp5_ASAP7_75t_L g3771 ( 
.A(n_3558),
.B(n_3534),
.Y(n_3771)
);

AOI21xp5_ASAP7_75t_L g3772 ( 
.A1(n_3593),
.A2(n_1993),
.B(n_1992),
.Y(n_3772)
);

AOI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_3607),
.A2(n_1997),
.B(n_1995),
.Y(n_3773)
);

CKINVDCx5p33_ASAP7_75t_R g3774 ( 
.A(n_3633),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3515),
.B(n_2226),
.Y(n_3775)
);

AOI21xp5_ASAP7_75t_L g3776 ( 
.A1(n_3617),
.A2(n_3580),
.B(n_3600),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3519),
.B(n_2228),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3511),
.A2(n_2028),
.B(n_2024),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_SL g3779 ( 
.A(n_3592),
.B(n_2231),
.Y(n_3779)
);

NAND2xp33_ASAP7_75t_L g3780 ( 
.A(n_3752),
.B(n_2236),
.Y(n_3780)
);

AOI21xp5_ASAP7_75t_L g3781 ( 
.A1(n_3522),
.A2(n_2071),
.B(n_2057),
.Y(n_3781)
);

O2A1O1Ixp33_ASAP7_75t_L g3782 ( 
.A1(n_3503),
.A2(n_2077),
.B(n_2080),
.C(n_2074),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_L g3783 ( 
.A(n_3508),
.B(n_2238),
.Y(n_3783)
);

BUFx12f_ASAP7_75t_L g3784 ( 
.A(n_3697),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3516),
.B(n_2241),
.Y(n_3785)
);

OAI21xp5_ASAP7_75t_L g3786 ( 
.A1(n_3484),
.A2(n_2086),
.B(n_2083),
.Y(n_3786)
);

OAI22xp5_ASAP7_75t_L g3787 ( 
.A1(n_3518),
.A2(n_2246),
.B1(n_2248),
.B2(n_2244),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_SL g3788 ( 
.A(n_3582),
.B(n_2249),
.Y(n_3788)
);

AOI21xp5_ASAP7_75t_L g3789 ( 
.A1(n_3528),
.A2(n_2098),
.B(n_2088),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_3487),
.B(n_2253),
.Y(n_3790)
);

NAND2xp33_ASAP7_75t_L g3791 ( 
.A(n_3752),
.B(n_2257),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3489),
.B(n_2259),
.Y(n_3792)
);

BUFx12f_ASAP7_75t_L g3793 ( 
.A(n_3540),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_3501),
.B(n_2261),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_SL g3795 ( 
.A(n_3690),
.B(n_3638),
.Y(n_3795)
);

CKINVDCx10_ASAP7_75t_R g3796 ( 
.A(n_3596),
.Y(n_3796)
);

NOR2x1p5_ASAP7_75t_SL g3797 ( 
.A(n_3752),
.B(n_2102),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3482),
.Y(n_3798)
);

INVx2_ASAP7_75t_L g3799 ( 
.A(n_3493),
.Y(n_3799)
);

O2A1O1Ixp33_ASAP7_75t_L g3800 ( 
.A1(n_3521),
.A2(n_2114),
.B(n_2118),
.C(n_2111),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3762),
.B(n_2286),
.Y(n_3801)
);

NOR2xp67_ASAP7_75t_L g3802 ( 
.A(n_3761),
.B(n_2262),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3504),
.B(n_2266),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3488),
.Y(n_3804)
);

BUFx12f_ASAP7_75t_L g3805 ( 
.A(n_3569),
.Y(n_3805)
);

OAI22xp5_ASAP7_75t_L g3806 ( 
.A1(n_3490),
.A2(n_2273),
.B1(n_2275),
.B2(n_2271),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_L g3807 ( 
.A(n_3507),
.B(n_2279),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_3509),
.B(n_2284),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_SL g3809 ( 
.A(n_3602),
.B(n_2285),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3492),
.Y(n_3810)
);

NOR2xp33_ASAP7_75t_L g3811 ( 
.A(n_3525),
.B(n_2287),
.Y(n_3811)
);

INVx2_ASAP7_75t_L g3812 ( 
.A(n_3513),
.Y(n_3812)
);

O2A1O1Ixp33_ASAP7_75t_SL g3813 ( 
.A1(n_3588),
.A2(n_2127),
.B(n_2128),
.C(n_2123),
.Y(n_3813)
);

BUFx3_ASAP7_75t_L g3814 ( 
.A(n_3506),
.Y(n_3814)
);

AOI21xp5_ASAP7_75t_L g3815 ( 
.A1(n_3578),
.A2(n_2135),
.B(n_2131),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_3485),
.B(n_2288),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_3520),
.Y(n_3817)
);

AOI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_3576),
.A2(n_2140),
.B(n_2139),
.Y(n_3818)
);

NOR2xp33_ASAP7_75t_L g3819 ( 
.A(n_3549),
.B(n_2293),
.Y(n_3819)
);

AOI21xp5_ASAP7_75t_L g3820 ( 
.A1(n_3538),
.A2(n_2142),
.B(n_2141),
.Y(n_3820)
);

AO21x1_ASAP7_75t_L g3821 ( 
.A1(n_3725),
.A2(n_2151),
.B(n_2145),
.Y(n_3821)
);

OAI22xp5_ASAP7_75t_L g3822 ( 
.A1(n_3495),
.A2(n_2297),
.B1(n_2299),
.B2(n_2296),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3497),
.Y(n_3823)
);

AO21x1_ASAP7_75t_L g3824 ( 
.A1(n_3486),
.A2(n_2158),
.B(n_2155),
.Y(n_3824)
);

A2O1A1Ixp33_ASAP7_75t_L g3825 ( 
.A1(n_3595),
.A2(n_2166),
.B(n_2177),
.C(n_2161),
.Y(n_3825)
);

OAI22xp5_ASAP7_75t_L g3826 ( 
.A1(n_3531),
.A2(n_2305),
.B1(n_2306),
.B2(n_2303),
.Y(n_3826)
);

OAI21xp5_ASAP7_75t_L g3827 ( 
.A1(n_3584),
.A2(n_2207),
.B(n_2193),
.Y(n_3827)
);

NOR2xp33_ASAP7_75t_L g3828 ( 
.A(n_3721),
.B(n_2307),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3537),
.B(n_2310),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3550),
.B(n_2313),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3738),
.B(n_2314),
.Y(n_3831)
);

AND2x2_ASAP7_75t_L g3832 ( 
.A(n_3514),
.B(n_2286),
.Y(n_3832)
);

OAI21xp33_ASAP7_75t_L g3833 ( 
.A1(n_3601),
.A2(n_3500),
.B(n_3499),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_L g3834 ( 
.A(n_3746),
.B(n_2316),
.Y(n_3834)
);

AO21x1_ASAP7_75t_L g3835 ( 
.A1(n_3724),
.A2(n_2239),
.B(n_2233),
.Y(n_3835)
);

AO21x1_ASAP7_75t_L g3836 ( 
.A1(n_3735),
.A2(n_2242),
.B(n_2240),
.Y(n_3836)
);

OAI22xp5_ASAP7_75t_L g3837 ( 
.A1(n_3758),
.A2(n_2319),
.B1(n_2321),
.B2(n_2317),
.Y(n_3837)
);

BUFx2_ASAP7_75t_L g3838 ( 
.A(n_3635),
.Y(n_3838)
);

OAI21xp33_ASAP7_75t_L g3839 ( 
.A1(n_3510),
.A2(n_2324),
.B(n_2322),
.Y(n_3839)
);

AOI21xp5_ASAP7_75t_L g3840 ( 
.A1(n_3533),
.A2(n_2254),
.B(n_2243),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3728),
.B(n_2328),
.Y(n_3841)
);

A2O1A1Ixp33_ASAP7_75t_L g3842 ( 
.A1(n_3666),
.A2(n_2265),
.B(n_2268),
.C(n_2258),
.Y(n_3842)
);

NOR2xp33_ASAP7_75t_L g3843 ( 
.A(n_3729),
.B(n_2333),
.Y(n_3843)
);

AOI22xp33_ASAP7_75t_L g3844 ( 
.A1(n_3575),
.A2(n_2280),
.B1(n_2282),
.B2(n_2269),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3532),
.Y(n_3845)
);

NAND2x1_ASAP7_75t_L g3846 ( 
.A(n_3545),
.B(n_2298),
.Y(n_3846)
);

AOI22xp5_ASAP7_75t_L g3847 ( 
.A1(n_3502),
.A2(n_2337),
.B1(n_2341),
.B2(n_2336),
.Y(n_3847)
);

AO21x1_ASAP7_75t_L g3848 ( 
.A1(n_3739),
.A2(n_3753),
.B(n_3748),
.Y(n_3848)
);

INVx3_ASAP7_75t_L g3849 ( 
.A(n_3517),
.Y(n_3849)
);

A2O1A1Ixp33_ASAP7_75t_L g3850 ( 
.A1(n_3641),
.A2(n_2309),
.B(n_2311),
.C(n_2308),
.Y(n_3850)
);

OAI21xp5_ASAP7_75t_L g3851 ( 
.A1(n_3722),
.A2(n_2325),
.B(n_2318),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_3734),
.B(n_2342),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3591),
.Y(n_3853)
);

INVx3_ASAP7_75t_L g3854 ( 
.A(n_3498),
.Y(n_3854)
);

NAND2x1_ASAP7_75t_L g3855 ( 
.A(n_3552),
.B(n_2326),
.Y(n_3855)
);

NOR2xp33_ASAP7_75t_L g3856 ( 
.A(n_3737),
.B(n_2347),
.Y(n_3856)
);

O2A1O1Ixp33_ASAP7_75t_L g3857 ( 
.A1(n_3527),
.A2(n_2334),
.B(n_2335),
.C(n_2332),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_SL g3858 ( 
.A(n_3727),
.B(n_2350),
.Y(n_3858)
);

AOI21xp5_ASAP7_75t_L g3859 ( 
.A1(n_3544),
.A2(n_2340),
.B(n_2338),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3740),
.B(n_2351),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3754),
.B(n_2353),
.Y(n_3861)
);

AOI22xp5_ASAP7_75t_L g3862 ( 
.A1(n_3502),
.A2(n_2355),
.B1(n_2357),
.B2(n_2354),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3756),
.B(n_2360),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3763),
.B(n_2361),
.Y(n_3864)
);

AOI21xp5_ASAP7_75t_L g3865 ( 
.A1(n_3590),
.A2(n_2372),
.B(n_2368),
.Y(n_3865)
);

AOI21x1_ASAP7_75t_L g3866 ( 
.A1(n_3523),
.A2(n_3571),
.B(n_3567),
.Y(n_3866)
);

AOI22xp5_ASAP7_75t_L g3867 ( 
.A1(n_3502),
.A2(n_2366),
.B1(n_2369),
.B2(n_2364),
.Y(n_3867)
);

OAI22xp5_ASAP7_75t_L g3868 ( 
.A1(n_3731),
.A2(n_2373),
.B1(n_2375),
.B2(n_2371),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3565),
.B(n_2377),
.Y(n_3869)
);

NOR2xp67_ASAP7_75t_L g3870 ( 
.A(n_3662),
.B(n_2381),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_SL g3871 ( 
.A(n_3733),
.B(n_2383),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_3742),
.B(n_2385),
.Y(n_3872)
);

AOI21xp5_ASAP7_75t_L g3873 ( 
.A1(n_3570),
.A2(n_2388),
.B(n_2384),
.Y(n_3873)
);

OAI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_3750),
.A2(n_2398),
.B(n_2390),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_SL g3875 ( 
.A(n_3751),
.B(n_2387),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_3483),
.B(n_2389),
.Y(n_3876)
);

AOI21xp5_ASAP7_75t_L g3877 ( 
.A1(n_3574),
.A2(n_2411),
.B(n_2410),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_SL g3878 ( 
.A(n_3644),
.B(n_2391),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3624),
.Y(n_3879)
);

OAI21xp5_ASAP7_75t_L g3880 ( 
.A1(n_3648),
.A2(n_2415),
.B(n_2413),
.Y(n_3880)
);

AOI21xp5_ASAP7_75t_L g3881 ( 
.A1(n_3539),
.A2(n_2442),
.B(n_2417),
.Y(n_3881)
);

INVx2_ASAP7_75t_SL g3882 ( 
.A(n_3623),
.Y(n_3882)
);

BUFx6f_ASAP7_75t_L g3883 ( 
.A(n_3583),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3627),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3628),
.Y(n_3885)
);

NAND3xp33_ASAP7_75t_L g3886 ( 
.A(n_3536),
.B(n_2396),
.C(n_2395),
.Y(n_3886)
);

BUFx6f_ASAP7_75t_L g3887 ( 
.A(n_3583),
.Y(n_3887)
);

NAND2xp33_ASAP7_75t_L g3888 ( 
.A(n_3752),
.B(n_2400),
.Y(n_3888)
);

AOI21xp5_ASAP7_75t_L g3889 ( 
.A1(n_3542),
.A2(n_2450),
.B(n_2445),
.Y(n_3889)
);

AOI21xp33_ASAP7_75t_L g3890 ( 
.A1(n_3629),
.A2(n_2403),
.B(n_2401),
.Y(n_3890)
);

AOI21xp5_ASAP7_75t_L g3891 ( 
.A1(n_3759),
.A2(n_2456),
.B(n_2451),
.Y(n_3891)
);

HB1xp67_ASAP7_75t_L g3892 ( 
.A(n_3626),
.Y(n_3892)
);

AOI21xp5_ASAP7_75t_L g3893 ( 
.A1(n_3554),
.A2(n_2473),
.B(n_2459),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_SL g3894 ( 
.A(n_3512),
.B(n_2404),
.Y(n_3894)
);

HB1xp67_ASAP7_75t_L g3895 ( 
.A(n_3699),
.Y(n_3895)
);

AOI21xp5_ASAP7_75t_L g3896 ( 
.A1(n_3561),
.A2(n_2478),
.B(n_2475),
.Y(n_3896)
);

OAI21xp5_ASAP7_75t_L g3897 ( 
.A1(n_3586),
.A2(n_3562),
.B(n_3663),
.Y(n_3897)
);

AOI21xp5_ASAP7_75t_L g3898 ( 
.A1(n_3566),
.A2(n_2501),
.B(n_2500),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3643),
.Y(n_3899)
);

INVx1_ASAP7_75t_SL g3900 ( 
.A(n_3654),
.Y(n_3900)
);

AOI21xp33_ASAP7_75t_L g3901 ( 
.A1(n_3560),
.A2(n_2418),
.B(n_2416),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3556),
.B(n_2420),
.Y(n_3902)
);

INVx2_ASAP7_75t_L g3903 ( 
.A(n_3745),
.Y(n_3903)
);

NOR2xp33_ASAP7_75t_L g3904 ( 
.A(n_3505),
.B(n_2421),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_L g3905 ( 
.A(n_3597),
.B(n_2422),
.Y(n_3905)
);

NOR2xp33_ASAP7_75t_L g3906 ( 
.A(n_3494),
.B(n_3481),
.Y(n_3906)
);

OAI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_3749),
.A2(n_2530),
.B(n_2528),
.Y(n_3907)
);

AOI21xp5_ASAP7_75t_L g3908 ( 
.A1(n_3764),
.A2(n_2534),
.B(n_2533),
.Y(n_3908)
);

OAI21xp5_ASAP7_75t_L g3909 ( 
.A1(n_3768),
.A2(n_2538),
.B(n_2536),
.Y(n_3909)
);

NOR3xp33_ASAP7_75t_L g3910 ( 
.A(n_3715),
.B(n_2426),
.C(n_2425),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3646),
.Y(n_3911)
);

INVx4_ASAP7_75t_L g3912 ( 
.A(n_3623),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_L g3913 ( 
.A(n_3547),
.B(n_2427),
.Y(n_3913)
);

HB1xp67_ASAP7_75t_L g3914 ( 
.A(n_3730),
.Y(n_3914)
);

OAI321xp33_ASAP7_75t_L g3915 ( 
.A1(n_3767),
.A2(n_2562),
.A3(n_2551),
.B1(n_2566),
.B2(n_2553),
.C(n_2550),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_3585),
.B(n_2430),
.Y(n_3916)
);

AOI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3587),
.A2(n_2577),
.B(n_2572),
.Y(n_3917)
);

AOI21xp5_ASAP7_75t_L g3918 ( 
.A1(n_3632),
.A2(n_3625),
.B(n_3669),
.Y(n_3918)
);

NOR2xp33_ASAP7_75t_L g3919 ( 
.A(n_3696),
.B(n_3685),
.Y(n_3919)
);

INVx3_ASAP7_75t_L g3920 ( 
.A(n_3692),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3651),
.Y(n_3921)
);

AOI21xp5_ASAP7_75t_L g3922 ( 
.A1(n_3599),
.A2(n_2582),
.B(n_2581),
.Y(n_3922)
);

INVx2_ASAP7_75t_SL g3923 ( 
.A(n_3760),
.Y(n_3923)
);

OAI22xp5_ASAP7_75t_L g3924 ( 
.A1(n_3639),
.A2(n_2432),
.B1(n_2434),
.B2(n_2431),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_L g3925 ( 
.A(n_3686),
.B(n_2436),
.Y(n_3925)
);

AOI21xp5_ASAP7_75t_L g3926 ( 
.A1(n_3594),
.A2(n_2598),
.B(n_2596),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3655),
.Y(n_3927)
);

AOI21xp5_ASAP7_75t_L g3928 ( 
.A1(n_3535),
.A2(n_2605),
.B(n_2604),
.Y(n_3928)
);

AOI21xp5_ASAP7_75t_L g3929 ( 
.A1(n_3541),
.A2(n_2619),
.B(n_2615),
.Y(n_3929)
);

NOR2xp33_ASAP7_75t_L g3930 ( 
.A(n_3559),
.B(n_2443),
.Y(n_3930)
);

CKINVDCx5p33_ASAP7_75t_R g3931 ( 
.A(n_3671),
.Y(n_3931)
);

BUFx6f_ASAP7_75t_L g3932 ( 
.A(n_3730),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_L g3933 ( 
.A(n_3614),
.B(n_3530),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3656),
.B(n_2444),
.Y(n_3934)
);

AOI21xp5_ASAP7_75t_L g3935 ( 
.A1(n_3555),
.A2(n_2623),
.B(n_2620),
.Y(n_3935)
);

BUFx2_ASAP7_75t_L g3936 ( 
.A(n_3577),
.Y(n_3936)
);

NOR2xp33_ASAP7_75t_L g3937 ( 
.A(n_3677),
.B(n_2452),
.Y(n_3937)
);

NOR2xp33_ASAP7_75t_L g3938 ( 
.A(n_3720),
.B(n_2455),
.Y(n_3938)
);

O2A1O1Ixp5_ASAP7_75t_L g3939 ( 
.A1(n_3573),
.A2(n_2629),
.B(n_2634),
.C(n_2625),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3743),
.B(n_2460),
.Y(n_3940)
);

NOR2xp33_ASAP7_75t_L g3941 ( 
.A(n_3657),
.B(n_2461),
.Y(n_3941)
);

BUFx6f_ASAP7_75t_L g3942 ( 
.A(n_3692),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3647),
.Y(n_3943)
);

AO21x1_ASAP7_75t_L g3944 ( 
.A1(n_3579),
.A2(n_2662),
.B(n_407),
.Y(n_3944)
);

OAI22xp5_ASAP7_75t_L g3945 ( 
.A1(n_3524),
.A2(n_2463),
.B1(n_2464),
.B2(n_2462),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3665),
.Y(n_3946)
);

INVx3_ASAP7_75t_L g3947 ( 
.A(n_3692),
.Y(n_3947)
);

CKINVDCx10_ASAP7_75t_R g3948 ( 
.A(n_3723),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3744),
.B(n_2467),
.Y(n_3949)
);

AOI21xp5_ASAP7_75t_L g3950 ( 
.A1(n_3608),
.A2(n_2471),
.B(n_2469),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3661),
.Y(n_3951)
);

NOR3xp33_ASAP7_75t_L g3952 ( 
.A(n_3717),
.B(n_2480),
.C(n_2476),
.Y(n_3952)
);

NOR2xp33_ASAP7_75t_L g3953 ( 
.A(n_3660),
.B(n_2481),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_L g3954 ( 
.A(n_3757),
.B(n_3610),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_SL g3955 ( 
.A(n_3766),
.B(n_3615),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3618),
.B(n_2483),
.Y(n_3956)
);

AND2x2_ASAP7_75t_L g3957 ( 
.A(n_3664),
.B(n_2348),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_3680),
.B(n_2485),
.Y(n_3958)
);

INVx2_ASAP7_75t_L g3959 ( 
.A(n_3667),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3674),
.B(n_2486),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3653),
.B(n_2487),
.Y(n_3961)
);

AOI21xp5_ASAP7_75t_L g3962 ( 
.A1(n_3765),
.A2(n_2489),
.B(n_2488),
.Y(n_3962)
);

INVx2_ASAP7_75t_L g3963 ( 
.A(n_3668),
.Y(n_3963)
);

NAND3xp33_ASAP7_75t_L g3964 ( 
.A(n_3616),
.B(n_3645),
.C(n_3563),
.Y(n_3964)
);

NOR2xp33_ASAP7_75t_L g3965 ( 
.A(n_3631),
.B(n_2490),
.Y(n_3965)
);

AND2x2_ASAP7_75t_L g3966 ( 
.A(n_3679),
.B(n_2348),
.Y(n_3966)
);

OAI22xp5_ASAP7_75t_L g3967 ( 
.A1(n_3676),
.A2(n_2496),
.B1(n_2498),
.B2(n_2494),
.Y(n_3967)
);

AOI21xp5_ASAP7_75t_L g3968 ( 
.A1(n_3622),
.A2(n_2503),
.B(n_2502),
.Y(n_3968)
);

OAI21xp5_ASAP7_75t_L g3969 ( 
.A1(n_3702),
.A2(n_2509),
.B(n_2506),
.Y(n_3969)
);

BUFx4f_ASAP7_75t_L g3970 ( 
.A(n_3718),
.Y(n_3970)
);

AND2x4_ASAP7_75t_L g3971 ( 
.A(n_3705),
.B(n_2510),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_L g3972 ( 
.A(n_3659),
.B(n_2511),
.Y(n_3972)
);

BUFx6f_ASAP7_75t_L g3973 ( 
.A(n_3613),
.Y(n_3973)
);

INVx2_ASAP7_75t_L g3974 ( 
.A(n_3683),
.Y(n_3974)
);

NOR2xp33_ASAP7_75t_L g3975 ( 
.A(n_3755),
.B(n_2515),
.Y(n_3975)
);

AND2x2_ASAP7_75t_L g3976 ( 
.A(n_3694),
.B(n_2358),
.Y(n_3976)
);

AOI21xp5_ASAP7_75t_L g3977 ( 
.A1(n_3605),
.A2(n_2523),
.B(n_2520),
.Y(n_3977)
);

OAI21xp5_ASAP7_75t_L g3978 ( 
.A1(n_3526),
.A2(n_2529),
.B(n_2524),
.Y(n_3978)
);

INVxp67_ASAP7_75t_L g3979 ( 
.A(n_3649),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3714),
.B(n_2358),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_L g3981 ( 
.A(n_3689),
.B(n_2545),
.Y(n_3981)
);

OR2x2_ASAP7_75t_L g3982 ( 
.A(n_3726),
.B(n_2546),
.Y(n_3982)
);

NOR2xp33_ASAP7_75t_L g3983 ( 
.A(n_3747),
.B(n_2555),
.Y(n_3983)
);

O2A1O1Ixp33_ASAP7_75t_L g3984 ( 
.A1(n_3673),
.A2(n_2412),
.B(n_2414),
.C(n_2378),
.Y(n_3984)
);

AOI21xp33_ASAP7_75t_L g3985 ( 
.A1(n_3546),
.A2(n_2557),
.B(n_2556),
.Y(n_3985)
);

OAI21xp5_ASAP7_75t_L g3986 ( 
.A1(n_3706),
.A2(n_2561),
.B(n_2558),
.Y(n_3986)
);

BUFx3_ASAP7_75t_L g3987 ( 
.A(n_3551),
.Y(n_3987)
);

OAI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_3670),
.A2(n_2565),
.B(n_2564),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_SL g3989 ( 
.A(n_3630),
.B(n_2574),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_L g3990 ( 
.A(n_3695),
.B(n_2575),
.Y(n_3990)
);

AO21x1_ASAP7_75t_L g3991 ( 
.A1(n_3496),
.A2(n_409),
.B(n_408),
.Y(n_3991)
);

AOI21xp5_ASAP7_75t_L g3992 ( 
.A1(n_3609),
.A2(n_3611),
.B(n_3621),
.Y(n_3992)
);

INVx3_ASAP7_75t_L g3993 ( 
.A(n_3598),
.Y(n_3993)
);

AND2x4_ASAP7_75t_L g3994 ( 
.A(n_3701),
.B(n_2578),
.Y(n_3994)
);

O2A1O1Ixp5_ASAP7_75t_L g3995 ( 
.A1(n_3634),
.A2(n_2412),
.B(n_2414),
.C(n_2378),
.Y(n_3995)
);

O2A1O1Ixp5_ASAP7_75t_L g3996 ( 
.A1(n_3636),
.A2(n_2513),
.B(n_2518),
.C(n_2457),
.Y(n_3996)
);

NOR2xp33_ASAP7_75t_R g3997 ( 
.A(n_3681),
.B(n_2592),
.Y(n_3997)
);

BUFx6f_ASAP7_75t_L g3998 ( 
.A(n_3682),
.Y(n_3998)
);

INVx8_ASAP7_75t_L g3999 ( 
.A(n_3640),
.Y(n_3999)
);

OAI21xp5_ASAP7_75t_L g4000 ( 
.A1(n_3652),
.A2(n_2597),
.B(n_2595),
.Y(n_4000)
);

NOR2x1_ASAP7_75t_L g4001 ( 
.A(n_3619),
.B(n_2584),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3732),
.B(n_2601),
.Y(n_4002)
);

AOI21xp5_ASAP7_75t_L g4003 ( 
.A1(n_3918),
.A2(n_3650),
.B(n_3642),
.Y(n_4003)
);

O2A1O1Ixp33_ASAP7_75t_L g4004 ( 
.A1(n_3833),
.A2(n_3716),
.B(n_3553),
.C(n_3589),
.Y(n_4004)
);

OR2x2_ASAP7_75t_L g4005 ( 
.A(n_3771),
.B(n_3704),
.Y(n_4005)
);

AOI21xp33_ASAP7_75t_L g4006 ( 
.A1(n_3819),
.A2(n_3919),
.B(n_3843),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3921),
.Y(n_4007)
);

AOI21xp5_ASAP7_75t_L g4008 ( 
.A1(n_3776),
.A2(n_3637),
.B(n_3693),
.Y(n_4008)
);

BUFx6f_ASAP7_75t_L g4009 ( 
.A(n_3942),
.Y(n_4009)
);

A2O1A1Ixp33_ASAP7_75t_L g4010 ( 
.A1(n_3906),
.A2(n_3698),
.B(n_3678),
.C(n_3658),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_3828),
.B(n_3604),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_3856),
.B(n_3564),
.Y(n_4012)
);

INVxp67_ASAP7_75t_L g4013 ( 
.A(n_3892),
.Y(n_4013)
);

NOR2xp33_ASAP7_75t_SL g4014 ( 
.A(n_3784),
.B(n_3719),
.Y(n_4014)
);

INVx2_ASAP7_75t_L g4015 ( 
.A(n_3798),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3804),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_SL g4017 ( 
.A(n_3795),
.B(n_3703),
.Y(n_4017)
);

AOI22xp33_ASAP7_75t_L g4018 ( 
.A1(n_3938),
.A2(n_3713),
.B1(n_3709),
.B2(n_3710),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_3810),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_SL g4020 ( 
.A(n_3954),
.B(n_3933),
.Y(n_4020)
);

AOI21xp5_ASAP7_75t_L g4021 ( 
.A1(n_3897),
.A2(n_3791),
.B(n_3780),
.Y(n_4021)
);

INVx2_ASAP7_75t_L g4022 ( 
.A(n_3823),
.Y(n_4022)
);

INVx3_ASAP7_75t_L g4023 ( 
.A(n_3814),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3783),
.B(n_3675),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3853),
.Y(n_4025)
);

INVx2_ASAP7_75t_L g4026 ( 
.A(n_3879),
.Y(n_4026)
);

BUFx6f_ASAP7_75t_L g4027 ( 
.A(n_3942),
.Y(n_4027)
);

HB1xp67_ASAP7_75t_L g4028 ( 
.A(n_3936),
.Y(n_4028)
);

NOR2xp33_ASAP7_75t_L g4029 ( 
.A(n_3811),
.B(n_3688),
.Y(n_4029)
);

OAI22xp33_ASAP7_75t_L g4030 ( 
.A1(n_3785),
.A2(n_3741),
.B1(n_3612),
.B2(n_3700),
.Y(n_4030)
);

INVx2_ASAP7_75t_L g4031 ( 
.A(n_3884),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3885),
.Y(n_4032)
);

BUFx6f_ASAP7_75t_L g4033 ( 
.A(n_3883),
.Y(n_4033)
);

AND3x1_ASAP7_75t_SL g4034 ( 
.A(n_3899),
.B(n_3691),
.C(n_3687),
.Y(n_4034)
);

INVx3_ASAP7_75t_L g4035 ( 
.A(n_3849),
.Y(n_4035)
);

OAI22xp5_ASAP7_75t_L g4036 ( 
.A1(n_3911),
.A2(n_3684),
.B1(n_3603),
.B2(n_3620),
.Y(n_4036)
);

OR2x6_ASAP7_75t_L g4037 ( 
.A(n_3999),
.B(n_3912),
.Y(n_4037)
);

AOI21xp5_ASAP7_75t_L g4038 ( 
.A1(n_3888),
.A2(n_3708),
.B(n_3707),
.Y(n_4038)
);

O2A1O1Ixp33_ASAP7_75t_SL g4039 ( 
.A1(n_3842),
.A2(n_3712),
.B(n_3672),
.C(n_3572),
.Y(n_4039)
);

A2O1A1Ixp33_ASAP7_75t_L g4040 ( 
.A1(n_3851),
.A2(n_3568),
.B(n_3606),
.C(n_3557),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_SL g4041 ( 
.A(n_3931),
.B(n_3529),
.Y(n_4041)
);

AND2x4_ASAP7_75t_L g4042 ( 
.A(n_3854),
.B(n_3612),
.Y(n_4042)
);

A2O1A1Ixp33_ASAP7_75t_L g4043 ( 
.A1(n_3874),
.A2(n_3548),
.B(n_2603),
.C(n_2606),
.Y(n_4043)
);

BUFx3_ASAP7_75t_L g4044 ( 
.A(n_3883),
.Y(n_4044)
);

BUFx3_ASAP7_75t_L g4045 ( 
.A(n_3932),
.Y(n_4045)
);

BUFx2_ASAP7_75t_L g4046 ( 
.A(n_3932),
.Y(n_4046)
);

NOR2xp33_ASAP7_75t_R g4047 ( 
.A(n_3774),
.B(n_3491),
.Y(n_4047)
);

O2A1O1Ixp33_ASAP7_75t_L g4048 ( 
.A1(n_3890),
.A2(n_3800),
.B(n_3782),
.C(n_3880),
.Y(n_4048)
);

O2A1O1Ixp33_ASAP7_75t_L g4049 ( 
.A1(n_3975),
.A2(n_3711),
.B(n_3543),
.C(n_2588),
.Y(n_4049)
);

NOR2xp33_ASAP7_75t_L g4050 ( 
.A(n_3913),
.B(n_3841),
.Y(n_4050)
);

AOI21xp5_ASAP7_75t_L g4051 ( 
.A1(n_3848),
.A2(n_2609),
.B(n_2602),
.Y(n_4051)
);

INVx2_ASAP7_75t_L g4052 ( 
.A(n_3799),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_3852),
.B(n_2611),
.Y(n_4053)
);

O2A1O1Ixp33_ASAP7_75t_L g4054 ( 
.A1(n_3983),
.A2(n_2588),
.B(n_2584),
.C(n_2614),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_3860),
.B(n_2618),
.Y(n_4055)
);

INVx2_ASAP7_75t_L g4056 ( 
.A(n_3812),
.Y(n_4056)
);

OAI21xp33_ASAP7_75t_L g4057 ( 
.A1(n_3980),
.A2(n_2624),
.B(n_2622),
.Y(n_4057)
);

BUFx12f_ASAP7_75t_L g4058 ( 
.A(n_3793),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3817),
.Y(n_4059)
);

A2O1A1Ixp33_ASAP7_75t_L g4060 ( 
.A1(n_3964),
.A2(n_2627),
.B(n_2628),
.C(n_2626),
.Y(n_4060)
);

AND3x1_ASAP7_75t_SL g4061 ( 
.A(n_3927),
.B(n_2631),
.C(n_2630),
.Y(n_4061)
);

NOR2x1p5_ASAP7_75t_L g4062 ( 
.A(n_3805),
.B(n_2633),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_SL g4063 ( 
.A(n_3941),
.B(n_2638),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3861),
.B(n_2640),
.Y(n_4064)
);

HB1xp67_ASAP7_75t_L g4065 ( 
.A(n_3895),
.Y(n_4065)
);

INVx3_ASAP7_75t_L g4066 ( 
.A(n_3987),
.Y(n_4066)
);

A2O1A1Ixp33_ASAP7_75t_L g4067 ( 
.A1(n_3904),
.A2(n_2645),
.B(n_2646),
.C(n_2644),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_L g4068 ( 
.A(n_3863),
.B(n_2647),
.Y(n_4068)
);

NOR2xp33_ASAP7_75t_L g4069 ( 
.A(n_3864),
.B(n_2648),
.Y(n_4069)
);

NOR2xp33_ASAP7_75t_L g4070 ( 
.A(n_3916),
.B(n_2652),
.Y(n_4070)
);

NAND2x1_ASAP7_75t_L g4071 ( 
.A(n_3920),
.B(n_412),
.Y(n_4071)
);

AND2x4_ASAP7_75t_L g4072 ( 
.A(n_3882),
.B(n_2654),
.Y(n_4072)
);

AO21x1_ASAP7_75t_L g4073 ( 
.A1(n_3786),
.A2(n_413),
.B(n_412),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3845),
.Y(n_4074)
);

OAI22xp5_ASAP7_75t_L g4075 ( 
.A1(n_3790),
.A2(n_2658),
.B1(n_2659),
.B2(n_2656),
.Y(n_4075)
);

INVx2_ASAP7_75t_L g4076 ( 
.A(n_3903),
.Y(n_4076)
);

AO21x2_ASAP7_75t_L g4077 ( 
.A1(n_3773),
.A2(n_1),
.B(n_2),
.Y(n_4077)
);

INVx4_ASAP7_75t_L g4078 ( 
.A(n_3887),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_3801),
.B(n_3832),
.Y(n_4079)
);

AOI21xp5_ASAP7_75t_L g4080 ( 
.A1(n_3792),
.A2(n_2661),
.B(n_414),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_SL g4081 ( 
.A(n_3953),
.B(n_413),
.Y(n_4081)
);

A2O1A1Ixp33_ASAP7_75t_L g4082 ( 
.A1(n_3937),
.A2(n_3),
.B(n_1),
.C(n_2),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_L g4083 ( 
.A(n_3794),
.B(n_3803),
.Y(n_4083)
);

OAI22xp5_ASAP7_75t_L g4084 ( 
.A1(n_3807),
.A2(n_417),
.B1(n_418),
.B2(n_416),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_3808),
.B(n_1),
.Y(n_4085)
);

A2O1A1Ixp33_ASAP7_75t_L g4086 ( 
.A1(n_3930),
.A2(n_4),
.B(n_2),
.C(n_3),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_L g4087 ( 
.A(n_3816),
.B(n_3),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_3946),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3943),
.Y(n_4089)
);

OR2x2_ASAP7_75t_L g4090 ( 
.A(n_3958),
.B(n_4),
.Y(n_4090)
);

OR2x4_ASAP7_75t_L g4091 ( 
.A(n_3965),
.B(n_4),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_3869),
.B(n_5),
.Y(n_4092)
);

OAI22xp5_ASAP7_75t_L g4093 ( 
.A1(n_3872),
.A2(n_420),
.B1(n_421),
.B2(n_419),
.Y(n_4093)
);

BUFx6f_ASAP7_75t_L g4094 ( 
.A(n_3887),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_3974),
.Y(n_4095)
);

INVx5_ASAP7_75t_L g4096 ( 
.A(n_3947),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3876),
.B(n_5),
.Y(n_4097)
);

NOR2xp33_ASAP7_75t_L g4098 ( 
.A(n_3788),
.B(n_420),
.Y(n_4098)
);

BUFx2_ASAP7_75t_L g4099 ( 
.A(n_3838),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_SL g4100 ( 
.A(n_3979),
.B(n_422),
.Y(n_4100)
);

BUFx2_ASAP7_75t_L g4101 ( 
.A(n_3914),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_3925),
.B(n_5),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3951),
.Y(n_4103)
);

BUFx3_ASAP7_75t_L g4104 ( 
.A(n_3973),
.Y(n_4104)
);

O2A1O1Ixp33_ASAP7_75t_L g4105 ( 
.A1(n_3901),
.A2(n_424),
.B(n_425),
.C(n_423),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_3959),
.Y(n_4106)
);

HB1xp67_ASAP7_75t_L g4107 ( 
.A(n_3973),
.Y(n_4107)
);

INVx2_ASAP7_75t_L g4108 ( 
.A(n_3963),
.Y(n_4108)
);

BUFx6f_ASAP7_75t_L g4109 ( 
.A(n_3998),
.Y(n_4109)
);

AOI21xp5_ASAP7_75t_L g4110 ( 
.A1(n_3809),
.A2(n_424),
.B(n_423),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_3846),
.Y(n_4111)
);

A2O1A1Ixp33_ASAP7_75t_L g4112 ( 
.A1(n_3797),
.A2(n_8),
.B(n_6),
.C(n_7),
.Y(n_4112)
);

INVx3_ASAP7_75t_SL g4113 ( 
.A(n_3769),
.Y(n_4113)
);

HB1xp67_ASAP7_75t_L g4114 ( 
.A(n_3998),
.Y(n_4114)
);

NOR3xp33_ASAP7_75t_SL g4115 ( 
.A(n_3839),
.B(n_6),
.C(n_7),
.Y(n_4115)
);

NOR2xp33_ASAP7_75t_L g4116 ( 
.A(n_3900),
.B(n_426),
.Y(n_4116)
);

NAND2x1p5_ASAP7_75t_L g4117 ( 
.A(n_3993),
.B(n_428),
.Y(n_4117)
);

NOR2xp33_ASAP7_75t_L g4118 ( 
.A(n_3961),
.B(n_429),
.Y(n_4118)
);

O2A1O1Ixp33_ASAP7_75t_L g4119 ( 
.A1(n_3825),
.A2(n_431),
.B(n_432),
.C(n_430),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_SL g4120 ( 
.A(n_3957),
.B(n_430),
.Y(n_4120)
);

AOI22xp5_ASAP7_75t_L g4121 ( 
.A1(n_3910),
.A2(n_433),
.B1(n_434),
.B2(n_431),
.Y(n_4121)
);

INVx2_ASAP7_75t_L g4122 ( 
.A(n_3855),
.Y(n_4122)
);

HB1xp67_ASAP7_75t_L g4123 ( 
.A(n_3923),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_L g4124 ( 
.A(n_3829),
.B(n_7),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_3905),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_L g4126 ( 
.A(n_3830),
.B(n_8),
.Y(n_4126)
);

BUFx2_ASAP7_75t_L g4127 ( 
.A(n_3994),
.Y(n_4127)
);

AOI21xp5_ASAP7_75t_L g4128 ( 
.A1(n_3858),
.A2(n_3875),
.B(n_3871),
.Y(n_4128)
);

INVx3_ASAP7_75t_L g4129 ( 
.A(n_3970),
.Y(n_4129)
);

OAI21xp33_ASAP7_75t_L g4130 ( 
.A1(n_3787),
.A2(n_9),
.B(n_10),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_3831),
.B(n_9),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_SL g4132 ( 
.A(n_3966),
.B(n_433),
.Y(n_4132)
);

BUFx6f_ASAP7_75t_L g4133 ( 
.A(n_3999),
.Y(n_4133)
);

A2O1A1Ixp33_ASAP7_75t_L g4134 ( 
.A1(n_4002),
.A2(n_12),
.B(n_9),
.C(n_11),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_3976),
.B(n_434),
.Y(n_4135)
);

NAND2xp33_ASAP7_75t_SL g4136 ( 
.A(n_3997),
.B(n_3955),
.Y(n_4136)
);

O2A1O1Ixp33_ASAP7_75t_L g4137 ( 
.A1(n_3850),
.A2(n_436),
.B(n_437),
.C(n_435),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_3834),
.B(n_11),
.Y(n_4138)
);

BUFx2_ASAP7_75t_SL g4139 ( 
.A(n_3802),
.Y(n_4139)
);

AOI22xp33_ASAP7_75t_L g4140 ( 
.A1(n_3886),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_4140)
);

AOI22xp33_ASAP7_75t_L g4141 ( 
.A1(n_3978),
.A2(n_3982),
.B1(n_3940),
.B2(n_3949),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_3772),
.B(n_3770),
.Y(n_4142)
);

BUFx6f_ASAP7_75t_L g4143 ( 
.A(n_3971),
.Y(n_4143)
);

BUFx6f_ASAP7_75t_L g4144 ( 
.A(n_3894),
.Y(n_4144)
);

OAI22x1_ASAP7_75t_L g4145 ( 
.A1(n_4001),
.A2(n_3779),
.B1(n_3862),
.B2(n_3847),
.Y(n_4145)
);

NAND2x1_ASAP7_75t_L g4146 ( 
.A(n_3992),
.B(n_439),
.Y(n_4146)
);

OAI22x1_ASAP7_75t_L g4147 ( 
.A1(n_3867),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_4147)
);

NOR2xp33_ASAP7_75t_L g4148 ( 
.A(n_3972),
.B(n_439),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_L g4149 ( 
.A(n_3844),
.B(n_13),
.Y(n_4149)
);

CKINVDCx5p33_ASAP7_75t_R g4150 ( 
.A(n_3796),
.Y(n_4150)
);

INVx2_ASAP7_75t_L g4151 ( 
.A(n_3934),
.Y(n_4151)
);

AOI21xp5_ASAP7_75t_L g4152 ( 
.A1(n_3878),
.A2(n_441),
.B(n_440),
.Y(n_4152)
);

NAND3xp33_ASAP7_75t_SL g4153 ( 
.A(n_3857),
.B(n_15),
.C(n_16),
.Y(n_4153)
);

AOI21xp5_ASAP7_75t_L g4154 ( 
.A1(n_3968),
.A2(n_443),
.B(n_442),
.Y(n_4154)
);

AOI21xp5_ASAP7_75t_L g4155 ( 
.A1(n_3977),
.A2(n_444),
.B(n_442),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3981),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3990),
.Y(n_4157)
);

BUFx8_ASAP7_75t_SL g4158 ( 
.A(n_3948),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3827),
.Y(n_4159)
);

O2A1O1Ixp33_ASAP7_75t_L g4160 ( 
.A1(n_3985),
.A2(n_445),
.B(n_446),
.C(n_444),
.Y(n_4160)
);

AO22x1_ASAP7_75t_L g4161 ( 
.A1(n_3952),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_4161)
);

INVx2_ASAP7_75t_L g4162 ( 
.A(n_3960),
.Y(n_4162)
);

OAI22xp5_ASAP7_75t_L g4163 ( 
.A1(n_3775),
.A2(n_447),
.B1(n_448),
.B2(n_445),
.Y(n_4163)
);

AND2x2_ASAP7_75t_L g4164 ( 
.A(n_3988),
.B(n_447),
.Y(n_4164)
);

INVx3_ASAP7_75t_SL g4165 ( 
.A(n_3989),
.Y(n_4165)
);

NOR3xp33_ASAP7_75t_L g4166 ( 
.A(n_3996),
.B(n_3995),
.C(n_3902),
.Y(n_4166)
);

A2O1A1Ixp33_ASAP7_75t_L g4167 ( 
.A1(n_3969),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_4167)
);

AOI21xp5_ASAP7_75t_L g4168 ( 
.A1(n_3907),
.A2(n_452),
.B(n_451),
.Y(n_4168)
);

INVx4_ASAP7_75t_L g4169 ( 
.A(n_3870),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_L g4170 ( 
.A(n_3778),
.B(n_18),
.Y(n_4170)
);

AOI21xp5_ASAP7_75t_L g4171 ( 
.A1(n_3909),
.A2(n_453),
.B(n_451),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_L g4172 ( 
.A(n_3781),
.B(n_19),
.Y(n_4172)
);

BUFx2_ASAP7_75t_L g4173 ( 
.A(n_3777),
.Y(n_4173)
);

BUFx4f_ASAP7_75t_L g4174 ( 
.A(n_3835),
.Y(n_4174)
);

NAND2x1p5_ASAP7_75t_L g4175 ( 
.A(n_3893),
.B(n_455),
.Y(n_4175)
);

INVx2_ASAP7_75t_SL g4176 ( 
.A(n_3924),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_3873),
.Y(n_4177)
);

AOI21xp5_ASAP7_75t_L g4178 ( 
.A1(n_3926),
.A2(n_457),
.B(n_456),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_SL g4179 ( 
.A(n_3915),
.B(n_458),
.Y(n_4179)
);

NOR2xp33_ASAP7_75t_L g4180 ( 
.A(n_3868),
.B(n_460),
.Y(n_4180)
);

AOI22xp5_ASAP7_75t_L g4181 ( 
.A1(n_3836),
.A2(n_461),
.B1(n_462),
.B2(n_460),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_3789),
.B(n_21),
.Y(n_4182)
);

AOI21x1_ASAP7_75t_L g4183 ( 
.A1(n_3824),
.A2(n_463),
.B(n_462),
.Y(n_4183)
);

CKINVDCx8_ASAP7_75t_R g4184 ( 
.A(n_3939),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_3986),
.B(n_23),
.Y(n_4185)
);

NOR2xp33_ASAP7_75t_SL g4186 ( 
.A(n_3984),
.B(n_23),
.Y(n_4186)
);

AOI21xp5_ASAP7_75t_L g4187 ( 
.A1(n_3896),
.A2(n_466),
.B(n_464),
.Y(n_4187)
);

NOR2xp33_ASAP7_75t_L g4188 ( 
.A(n_3945),
.B(n_467),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_4000),
.B(n_24),
.Y(n_4189)
);

OAI22x1_ASAP7_75t_L g4190 ( 
.A1(n_3991),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_4190)
);

AOI21xp5_ASAP7_75t_L g4191 ( 
.A1(n_3898),
.A2(n_471),
.B(n_470),
.Y(n_4191)
);

CKINVDCx5p33_ASAP7_75t_R g4192 ( 
.A(n_3967),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_3877),
.Y(n_4193)
);

BUFx2_ASAP7_75t_L g4194 ( 
.A(n_3956),
.Y(n_4194)
);

OAI22x1_ASAP7_75t_L g4195 ( 
.A1(n_3944),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_4195)
);

HB1xp67_ASAP7_75t_L g4196 ( 
.A(n_3891),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_3840),
.B(n_28),
.Y(n_4197)
);

BUFx6f_ASAP7_75t_L g4198 ( 
.A(n_3820),
.Y(n_4198)
);

OAI22xp5_ASAP7_75t_L g4199 ( 
.A1(n_3962),
.A2(n_472),
.B1(n_473),
.B2(n_471),
.Y(n_4199)
);

BUFx6f_ASAP7_75t_L g4200 ( 
.A(n_3821),
.Y(n_4200)
);

NAND2xp33_ASAP7_75t_SL g4201 ( 
.A(n_3806),
.B(n_3822),
.Y(n_4201)
);

NOR2xp33_ASAP7_75t_L g4202 ( 
.A(n_3826),
.B(n_474),
.Y(n_4202)
);

BUFx6f_ASAP7_75t_L g4203 ( 
.A(n_3813),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_3859),
.B(n_30),
.Y(n_4204)
);

NOR2xp33_ASAP7_75t_L g4205 ( 
.A(n_3837),
.B(n_475),
.Y(n_4205)
);

BUFx6f_ASAP7_75t_L g4206 ( 
.A(n_3928),
.Y(n_4206)
);

BUFx12f_ASAP7_75t_L g4207 ( 
.A(n_3929),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_3865),
.B(n_31),
.Y(n_4208)
);

O2A1O1Ixp33_ASAP7_75t_L g4209 ( 
.A1(n_3917),
.A2(n_477),
.B(n_478),
.C(n_476),
.Y(n_4209)
);

O2A1O1Ixp33_ASAP7_75t_L g4210 ( 
.A1(n_3881),
.A2(n_479),
.B(n_480),
.C(n_478),
.Y(n_4210)
);

BUFx2_ASAP7_75t_L g4211 ( 
.A(n_3889),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_3922),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_3818),
.Y(n_4213)
);

AOI221xp5_ASAP7_75t_L g4214 ( 
.A1(n_3935),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.C(n_35),
.Y(n_4214)
);

BUFx2_ASAP7_75t_L g4215 ( 
.A(n_3815),
.Y(n_4215)
);

OAI22xp5_ASAP7_75t_L g4216 ( 
.A1(n_3950),
.A2(n_483),
.B1(n_484),
.B2(n_482),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_3908),
.Y(n_4217)
);

INVx8_ASAP7_75t_L g4218 ( 
.A(n_3784),
.Y(n_4218)
);

AO21x2_ASAP7_75t_L g4219 ( 
.A1(n_3848),
.A2(n_33),
.B(n_34),
.Y(n_4219)
);

O2A1O1Ixp5_ASAP7_75t_L g4220 ( 
.A1(n_3819),
.A2(n_485),
.B(n_486),
.C(n_484),
.Y(n_4220)
);

NOR2xp33_ASAP7_75t_SL g4221 ( 
.A(n_3919),
.B(n_34),
.Y(n_4221)
);

A2O1A1Ixp33_ASAP7_75t_L g4222 ( 
.A1(n_3833),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_4222)
);

NOR2xp33_ASAP7_75t_L g4223 ( 
.A(n_3919),
.B(n_485),
.Y(n_4223)
);

NOR2xp33_ASAP7_75t_L g4224 ( 
.A(n_3919),
.B(n_486),
.Y(n_4224)
);

AO32x2_ASAP7_75t_L g4225 ( 
.A1(n_3945),
.A2(n_38),
.A3(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_SL g4226 ( 
.A(n_3919),
.B(n_487),
.Y(n_4226)
);

OAI22xp5_ASAP7_75t_L g4227 ( 
.A1(n_3919),
.A2(n_489),
.B1(n_490),
.B2(n_488),
.Y(n_4227)
);

CKINVDCx5p33_ASAP7_75t_R g4228 ( 
.A(n_3796),
.Y(n_4228)
);

AOI21x1_ASAP7_75t_L g4229 ( 
.A1(n_3866),
.A2(n_491),
.B(n_490),
.Y(n_4229)
);

INVx2_ASAP7_75t_L g4230 ( 
.A(n_3798),
.Y(n_4230)
);

BUFx2_ASAP7_75t_L g4231 ( 
.A(n_3892),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_3771),
.B(n_36),
.Y(n_4232)
);

AOI21xp5_ASAP7_75t_L g4233 ( 
.A1(n_3918),
.A2(n_492),
.B(n_491),
.Y(n_4233)
);

O2A1O1Ixp5_ASAP7_75t_SL g4234 ( 
.A1(n_3827),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_4234)
);

AOI21xp5_ASAP7_75t_L g4235 ( 
.A1(n_3918),
.A2(n_494),
.B(n_493),
.Y(n_4235)
);

AOI21x1_ASAP7_75t_L g4236 ( 
.A1(n_3866),
.A2(n_496),
.B(n_495),
.Y(n_4236)
);

AND2x4_ASAP7_75t_L g4237 ( 
.A(n_3814),
.B(n_495),
.Y(n_4237)
);

HB1xp67_ASAP7_75t_L g4238 ( 
.A(n_3892),
.Y(n_4238)
);

O2A1O1Ixp33_ASAP7_75t_L g4239 ( 
.A1(n_3833),
.A2(n_499),
.B(n_500),
.C(n_498),
.Y(n_4239)
);

AOI21xp5_ASAP7_75t_L g4240 ( 
.A1(n_3918),
.A2(n_501),
.B(n_500),
.Y(n_4240)
);

AOI21x1_ASAP7_75t_L g4241 ( 
.A1(n_4021),
.A2(n_38),
.B(n_39),
.Y(n_4241)
);

NOR4xp25_ASAP7_75t_L g4242 ( 
.A(n_4006),
.B(n_42),
.C(n_40),
.D(n_41),
.Y(n_4242)
);

AOI21xp5_ASAP7_75t_L g4243 ( 
.A1(n_4003),
.A2(n_503),
.B(n_502),
.Y(n_4243)
);

AO31x2_ASAP7_75t_L g4244 ( 
.A1(n_4159),
.A2(n_44),
.A3(n_41),
.B(n_43),
.Y(n_4244)
);

AND2x4_ASAP7_75t_L g4245 ( 
.A(n_4023),
.B(n_4104),
.Y(n_4245)
);

OAI21xp5_ASAP7_75t_L g4246 ( 
.A1(n_4048),
.A2(n_43),
.B(n_44),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_4050),
.B(n_44),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_L g4248 ( 
.A(n_4020),
.B(n_45),
.Y(n_4248)
);

AO31x2_ASAP7_75t_L g4249 ( 
.A1(n_4073),
.A2(n_47),
.A3(n_45),
.B(n_46),
.Y(n_4249)
);

INVxp67_ASAP7_75t_L g4250 ( 
.A(n_4238),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_4015),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_L g4252 ( 
.A(n_4005),
.B(n_45),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_SL g4253 ( 
.A(n_4029),
.B(n_4012),
.Y(n_4253)
);

OAI21xp5_ASAP7_75t_L g4254 ( 
.A1(n_4070),
.A2(n_4069),
.B(n_4141),
.Y(n_4254)
);

INVxp67_ASAP7_75t_L g4255 ( 
.A(n_4231),
.Y(n_4255)
);

OAI21xp5_ASAP7_75t_L g4256 ( 
.A1(n_4011),
.A2(n_46),
.B(n_47),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_4083),
.B(n_46),
.Y(n_4257)
);

OR2x6_ASAP7_75t_L g4258 ( 
.A(n_4218),
.B(n_502),
.Y(n_4258)
);

CKINVDCx20_ASAP7_75t_R g4259 ( 
.A(n_4158),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_4019),
.Y(n_4260)
);

NAND3xp33_ASAP7_75t_SL g4261 ( 
.A(n_4221),
.B(n_48),
.C(n_49),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4022),
.Y(n_4262)
);

OAI21x1_ASAP7_75t_L g4263 ( 
.A1(n_4008),
.A2(n_50),
.B(n_51),
.Y(n_4263)
);

AOI21xp5_ASAP7_75t_L g4264 ( 
.A1(n_4142),
.A2(n_504),
.B(n_503),
.Y(n_4264)
);

BUFx3_ASAP7_75t_L g4265 ( 
.A(n_4109),
.Y(n_4265)
);

INVx2_ASAP7_75t_SL g4266 ( 
.A(n_4109),
.Y(n_4266)
);

BUFx2_ASAP7_75t_L g4267 ( 
.A(n_4099),
.Y(n_4267)
);

INVx2_ASAP7_75t_L g4268 ( 
.A(n_4026),
.Y(n_4268)
);

OAI22xp5_ASAP7_75t_L g4269 ( 
.A1(n_4223),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_4269)
);

NAND3xp33_ASAP7_75t_L g4270 ( 
.A(n_4224),
.B(n_51),
.C(n_52),
.Y(n_4270)
);

OAI21xp5_ASAP7_75t_L g4271 ( 
.A1(n_4189),
.A2(n_52),
.B(n_53),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4031),
.Y(n_4272)
);

OAI21x1_ASAP7_75t_L g4273 ( 
.A1(n_4146),
.A2(n_53),
.B(n_54),
.Y(n_4273)
);

NOR2x1_ASAP7_75t_SL g4274 ( 
.A(n_4139),
.B(n_4200),
.Y(n_4274)
);

AND2x4_ASAP7_75t_L g4275 ( 
.A(n_4066),
.B(n_506),
.Y(n_4275)
);

AOI21xp5_ASAP7_75t_L g4276 ( 
.A1(n_4038),
.A2(n_509),
.B(n_507),
.Y(n_4276)
);

OAI21xp5_ASAP7_75t_SL g4277 ( 
.A1(n_4049),
.A2(n_55),
.B(n_56),
.Y(n_4277)
);

INVx4_ASAP7_75t_L g4278 ( 
.A(n_4009),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_4230),
.Y(n_4279)
);

AOI21xp5_ASAP7_75t_L g4280 ( 
.A1(n_4136),
.A2(n_511),
.B(n_510),
.Y(n_4280)
);

AOI21x1_ASAP7_75t_SL g4281 ( 
.A1(n_4185),
.A2(n_57),
.B(n_58),
.Y(n_4281)
);

AOI21x1_ASAP7_75t_L g4282 ( 
.A1(n_4229),
.A2(n_58),
.B(n_59),
.Y(n_4282)
);

AOI21x1_ASAP7_75t_L g4283 ( 
.A1(n_4236),
.A2(n_4215),
.B(n_4211),
.Y(n_4283)
);

O2A1O1Ixp33_ASAP7_75t_SL g4284 ( 
.A1(n_4167),
.A2(n_511),
.B(n_512),
.C(n_510),
.Y(n_4284)
);

AOI21xp5_ASAP7_75t_L g4285 ( 
.A1(n_4024),
.A2(n_513),
.B(n_512),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4007),
.Y(n_4286)
);

NOR2xp67_ASAP7_75t_L g4287 ( 
.A(n_4169),
.B(n_60),
.Y(n_4287)
);

NOR2xp67_ASAP7_75t_L g4288 ( 
.A(n_4035),
.B(n_60),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_L g4289 ( 
.A(n_4125),
.B(n_61),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4016),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_L g4291 ( 
.A(n_4162),
.B(n_62),
.Y(n_4291)
);

AO21x2_ASAP7_75t_L g4292 ( 
.A1(n_4166),
.A2(n_62),
.B(n_63),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4025),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_4088),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_SL g4295 ( 
.A(n_4030),
.B(n_514),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4032),
.Y(n_4296)
);

NAND3xp33_ASAP7_75t_L g4297 ( 
.A(n_4180),
.B(n_63),
.C(n_64),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_L g4298 ( 
.A(n_4156),
.B(n_65),
.Y(n_4298)
);

OR2x2_ASAP7_75t_L g4299 ( 
.A(n_4232),
.B(n_514),
.Y(n_4299)
);

NAND2xp33_ASAP7_75t_L g4300 ( 
.A(n_4192),
.B(n_4133),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_4157),
.B(n_65),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_L g4302 ( 
.A(n_4151),
.B(n_4173),
.Y(n_4302)
);

A2O1A1Ixp33_ASAP7_75t_L g4303 ( 
.A1(n_4201),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_4303)
);

A2O1A1Ixp33_ASAP7_75t_L g4304 ( 
.A1(n_4004),
.A2(n_4054),
.B(n_4188),
.C(n_4148),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_L g4305 ( 
.A(n_4079),
.B(n_66),
.Y(n_4305)
);

NAND3x1_ASAP7_75t_L g4306 ( 
.A(n_4121),
.B(n_67),
.C(n_68),
.Y(n_4306)
);

O2A1O1Ixp33_ASAP7_75t_SL g4307 ( 
.A1(n_4222),
.A2(n_516),
.B(n_517),
.C(n_515),
.Y(n_4307)
);

NOR2xp33_ASAP7_75t_L g4308 ( 
.A(n_4013),
.B(n_515),
.Y(n_4308)
);

INVx5_ASAP7_75t_L g4309 ( 
.A(n_4033),
.Y(n_4309)
);

NOR2xp33_ASAP7_75t_SL g4310 ( 
.A(n_4150),
.B(n_68),
.Y(n_4310)
);

INVx2_ASAP7_75t_SL g4311 ( 
.A(n_4044),
.Y(n_4311)
);

AND2x4_ASAP7_75t_L g4312 ( 
.A(n_4037),
.B(n_4045),
.Y(n_4312)
);

NAND2xp5_ASAP7_75t_SL g4313 ( 
.A(n_4018),
.B(n_516),
.Y(n_4313)
);

AO21x2_ASAP7_75t_L g4314 ( 
.A1(n_4233),
.A2(n_4240),
.B(n_4235),
.Y(n_4314)
);

AOI211x1_ASAP7_75t_L g4315 ( 
.A1(n_4161),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_4315)
);

AOI22xp5_ASAP7_75t_L g4316 ( 
.A1(n_4098),
.A2(n_73),
.B1(n_70),
.B2(n_72),
.Y(n_4316)
);

INVx3_ASAP7_75t_L g4317 ( 
.A(n_4129),
.Y(n_4317)
);

AOI21xp5_ASAP7_75t_L g4318 ( 
.A1(n_4010),
.A2(n_519),
.B(n_518),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_L g4319 ( 
.A(n_4092),
.B(n_72),
.Y(n_4319)
);

NAND2xp5_ASAP7_75t_L g4320 ( 
.A(n_4085),
.B(n_74),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_4087),
.B(n_75),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_4102),
.B(n_75),
.Y(n_4322)
);

NAND2xp5_ASAP7_75t_L g4323 ( 
.A(n_4118),
.B(n_76),
.Y(n_4323)
);

A2O1A1Ixp33_ASAP7_75t_L g4324 ( 
.A1(n_4164),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_4089),
.Y(n_4325)
);

OAI21x1_ASAP7_75t_SL g4326 ( 
.A1(n_4168),
.A2(n_76),
.B(n_77),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_4097),
.B(n_78),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4059),
.Y(n_4328)
);

AND2x4_ASAP7_75t_L g4329 ( 
.A(n_4037),
.B(n_518),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_L g4330 ( 
.A(n_4194),
.B(n_79),
.Y(n_4330)
);

BUFx6f_ASAP7_75t_L g4331 ( 
.A(n_4009),
.Y(n_4331)
);

AOI211x1_ASAP7_75t_L g4332 ( 
.A1(n_4081),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_L g4333 ( 
.A(n_4053),
.B(n_81),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_L g4334 ( 
.A(n_4055),
.B(n_82),
.Y(n_4334)
);

AND2x6_ASAP7_75t_L g4335 ( 
.A(n_4203),
.B(n_520),
.Y(n_4335)
);

BUFx3_ASAP7_75t_L g4336 ( 
.A(n_4046),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4074),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_L g4338 ( 
.A(n_4064),
.B(n_83),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4103),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_4068),
.B(n_83),
.Y(n_4340)
);

AOI21xp5_ASAP7_75t_L g4341 ( 
.A1(n_4128),
.A2(n_523),
.B(n_522),
.Y(n_4341)
);

INVx2_ASAP7_75t_L g4342 ( 
.A(n_4052),
.Y(n_4342)
);

OAI22x1_ASAP7_75t_L g4343 ( 
.A1(n_4202),
.A2(n_4205),
.B1(n_4181),
.B2(n_4226),
.Y(n_4343)
);

AOI21xp5_ASAP7_75t_L g4344 ( 
.A1(n_4213),
.A2(n_525),
.B(n_524),
.Y(n_4344)
);

AO22x2_ASAP7_75t_L g4345 ( 
.A1(n_4153),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_4345)
);

OA22x2_ASAP7_75t_L g4346 ( 
.A1(n_4147),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_4346)
);

OAI21x1_ASAP7_75t_SL g4347 ( 
.A1(n_4171),
.A2(n_84),
.B(n_85),
.Y(n_4347)
);

INVx1_ASAP7_75t_L g4348 ( 
.A(n_4106),
.Y(n_4348)
);

OAI21x1_ASAP7_75t_L g4349 ( 
.A1(n_4217),
.A2(n_87),
.B(n_88),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4095),
.Y(n_4350)
);

OAI21x1_ASAP7_75t_L g4351 ( 
.A1(n_4177),
.A2(n_87),
.B(n_88),
.Y(n_4351)
);

AO31x2_ASAP7_75t_L g4352 ( 
.A1(n_4190),
.A2(n_92),
.A3(n_89),
.B(n_91),
.Y(n_4352)
);

AOI211x1_ASAP7_75t_L g4353 ( 
.A1(n_4130),
.A2(n_92),
.B(n_89),
.C(n_91),
.Y(n_4353)
);

OAI21x1_ASAP7_75t_L g4354 ( 
.A1(n_4193),
.A2(n_89),
.B(n_91),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_SL g4355 ( 
.A(n_4144),
.B(n_524),
.Y(n_4355)
);

AOI21xp5_ASAP7_75t_L g4356 ( 
.A1(n_4212),
.A2(n_526),
.B(n_525),
.Y(n_4356)
);

NOR2xp67_ASAP7_75t_SL g4357 ( 
.A(n_4058),
.B(n_93),
.Y(n_4357)
);

BUFx2_ASAP7_75t_L g4358 ( 
.A(n_4028),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_4056),
.Y(n_4359)
);

BUFx12f_ASAP7_75t_L g4360 ( 
.A(n_4228),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4076),
.Y(n_4361)
);

NAND3xp33_ASAP7_75t_L g4362 ( 
.A(n_4186),
.B(n_93),
.C(n_94),
.Y(n_4362)
);

NAND3xp33_ASAP7_75t_L g4363 ( 
.A(n_4086),
.B(n_94),
.C(n_95),
.Y(n_4363)
);

INVx2_ASAP7_75t_L g4364 ( 
.A(n_4108),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_SL g4365 ( 
.A(n_4144),
.B(n_527),
.Y(n_4365)
);

CKINVDCx5p33_ASAP7_75t_R g4366 ( 
.A(n_4047),
.Y(n_4366)
);

AOI21xp5_ASAP7_75t_L g4367 ( 
.A1(n_4196),
.A2(n_528),
.B(n_527),
.Y(n_4367)
);

OAI21x1_ASAP7_75t_L g4368 ( 
.A1(n_4111),
.A2(n_4122),
.B(n_4183),
.Y(n_4368)
);

AOI21xp5_ASAP7_75t_L g4369 ( 
.A1(n_4039),
.A2(n_530),
.B(n_529),
.Y(n_4369)
);

O2A1O1Ixp33_ASAP7_75t_L g4370 ( 
.A1(n_4082),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_4370)
);

OAI21x1_ASAP7_75t_L g4371 ( 
.A1(n_4234),
.A2(n_99),
.B(n_100),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4219),
.Y(n_4372)
);

AND2x4_ASAP7_75t_L g4373 ( 
.A(n_4101),
.B(n_4107),
.Y(n_4373)
);

OAI21x1_ASAP7_75t_L g4374 ( 
.A1(n_4154),
.A2(n_4155),
.B(n_4051),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_L g4375 ( 
.A(n_4124),
.B(n_100),
.Y(n_4375)
);

AOI21xp5_ASAP7_75t_SL g4376 ( 
.A1(n_4040),
.A2(n_531),
.B(n_529),
.Y(n_4376)
);

A2O1A1Ixp33_ASAP7_75t_L g4377 ( 
.A1(n_4080),
.A2(n_103),
.B(n_101),
.C(n_102),
.Y(n_4377)
);

NAND2x1p5_ASAP7_75t_L g4378 ( 
.A(n_4096),
.B(n_531),
.Y(n_4378)
);

AOI21xp5_ASAP7_75t_SL g4379 ( 
.A1(n_4239),
.A2(n_533),
.B(n_532),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_L g4380 ( 
.A(n_4126),
.B(n_101),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_4065),
.Y(n_4381)
);

OAI21xp5_ASAP7_75t_SL g4382 ( 
.A1(n_4140),
.A2(n_104),
.B(n_105),
.Y(n_4382)
);

OAI21xp5_ASAP7_75t_L g4383 ( 
.A1(n_4063),
.A2(n_105),
.B(n_106),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_4206),
.Y(n_4384)
);

NAND2xp5_ASAP7_75t_L g4385 ( 
.A(n_4131),
.B(n_106),
.Y(n_4385)
);

BUFx3_ASAP7_75t_L g4386 ( 
.A(n_4027),
.Y(n_4386)
);

AOI21xp5_ASAP7_75t_L g4387 ( 
.A1(n_4198),
.A2(n_533),
.B(n_532),
.Y(n_4387)
);

AOI21xp5_ASAP7_75t_L g4388 ( 
.A1(n_4198),
.A2(n_535),
.B(n_534),
.Y(n_4388)
);

OA21x2_ASAP7_75t_L g4389 ( 
.A1(n_4112),
.A2(n_107),
.B(n_108),
.Y(n_4389)
);

A2O1A1Ixp33_ASAP7_75t_L g4390 ( 
.A1(n_4176),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_4390)
);

AND2x6_ASAP7_75t_SL g4391 ( 
.A(n_4116),
.B(n_107),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4138),
.Y(n_4392)
);

OAI21xp33_ASAP7_75t_L g4393 ( 
.A1(n_4057),
.A2(n_109),
.B(n_110),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_L g4394 ( 
.A(n_4149),
.B(n_109),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_SL g4395 ( 
.A(n_4174),
.B(n_535),
.Y(n_4395)
);

INVx2_ASAP7_75t_L g4396 ( 
.A(n_4206),
.Y(n_4396)
);

OAI21xp5_ASAP7_75t_L g4397 ( 
.A1(n_4067),
.A2(n_110),
.B(n_111),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_4090),
.B(n_4017),
.Y(n_4398)
);

INVx2_ASAP7_75t_L g4399 ( 
.A(n_4077),
.Y(n_4399)
);

INVx2_ASAP7_75t_SL g4400 ( 
.A(n_4027),
.Y(n_4400)
);

OAI21x1_ASAP7_75t_L g4401 ( 
.A1(n_4220),
.A2(n_111),
.B(n_112),
.Y(n_4401)
);

OAI21x1_ASAP7_75t_L g4402 ( 
.A1(n_4187),
.A2(n_112),
.B(n_113),
.Y(n_4402)
);

OR2x6_ASAP7_75t_L g4403 ( 
.A(n_4218),
.B(n_536),
.Y(n_4403)
);

AOI21xp5_ASAP7_75t_L g4404 ( 
.A1(n_4145),
.A2(n_537),
.B(n_536),
.Y(n_4404)
);

INVx1_ASAP7_75t_SL g4405 ( 
.A(n_4123),
.Y(n_4405)
);

AOI21x1_ASAP7_75t_L g4406 ( 
.A1(n_4195),
.A2(n_113),
.B(n_114),
.Y(n_4406)
);

AOI21xp5_ASAP7_75t_L g4407 ( 
.A1(n_4179),
.A2(n_538),
.B(n_537),
.Y(n_4407)
);

NOR2xp33_ASAP7_75t_L g4408 ( 
.A(n_4041),
.B(n_538),
.Y(n_4408)
);

INVx3_ASAP7_75t_L g4409 ( 
.A(n_4078),
.Y(n_4409)
);

OAI22xp5_ASAP7_75t_L g4410 ( 
.A1(n_4036),
.A2(n_4184),
.B1(n_4091),
.B2(n_4115),
.Y(n_4410)
);

A2O1A1Ixp33_ASAP7_75t_L g4411 ( 
.A1(n_4110),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_4411)
);

OAI21x1_ASAP7_75t_L g4412 ( 
.A1(n_4191),
.A2(n_115),
.B(n_116),
.Y(n_4412)
);

INVx2_ASAP7_75t_L g4413 ( 
.A(n_4200),
.Y(n_4413)
);

NOR2xp33_ASAP7_75t_L g4414 ( 
.A(n_4165),
.B(n_539),
.Y(n_4414)
);

AO21x2_ASAP7_75t_L g4415 ( 
.A1(n_4178),
.A2(n_116),
.B(n_117),
.Y(n_4415)
);

NAND2xp5_ASAP7_75t_L g4416 ( 
.A(n_4143),
.B(n_117),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4170),
.Y(n_4417)
);

AOI21xp5_ASAP7_75t_L g4418 ( 
.A1(n_4160),
.A2(n_4119),
.B(n_4172),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_L g4419 ( 
.A(n_4143),
.B(n_4135),
.Y(n_4419)
);

HB1xp67_ASAP7_75t_L g4420 ( 
.A(n_4114),
.Y(n_4420)
);

AND2x4_ASAP7_75t_L g4421 ( 
.A(n_4133),
.B(n_4042),
.Y(n_4421)
);

NAND3xp33_ASAP7_75t_L g4422 ( 
.A(n_4105),
.B(n_117),
.C(n_118),
.Y(n_4422)
);

NOR4xp25_ASAP7_75t_L g4423 ( 
.A(n_4209),
.B(n_120),
.C(n_118),
.D(n_119),
.Y(n_4423)
);

NOR2xp33_ASAP7_75t_L g4424 ( 
.A(n_4120),
.B(n_4132),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4182),
.Y(n_4425)
);

AOI21xp5_ASAP7_75t_L g4426 ( 
.A1(n_4197),
.A2(n_540),
.B(n_539),
.Y(n_4426)
);

AND2x2_ASAP7_75t_L g4427 ( 
.A(n_4237),
.B(n_121),
.Y(n_4427)
);

O2A1O1Ixp33_ASAP7_75t_L g4428 ( 
.A1(n_4134),
.A2(n_124),
.B(n_122),
.C(n_123),
.Y(n_4428)
);

AOI21xp5_ASAP7_75t_SL g4429 ( 
.A1(n_4060),
.A2(n_541),
.B(n_540),
.Y(n_4429)
);

BUFx3_ASAP7_75t_L g4430 ( 
.A(n_4265),
.Y(n_4430)
);

CKINVDCx5p33_ASAP7_75t_R g4431 ( 
.A(n_4360),
.Y(n_4431)
);

NOR2xp67_ASAP7_75t_L g4432 ( 
.A(n_4317),
.B(n_4072),
.Y(n_4432)
);

AO21x2_ASAP7_75t_L g4433 ( 
.A1(n_4254),
.A2(n_4208),
.B(n_4204),
.Y(n_4433)
);

OAI21x1_ASAP7_75t_L g4434 ( 
.A1(n_4374),
.A2(n_4152),
.B(n_4175),
.Y(n_4434)
);

INVx2_ASAP7_75t_L g4435 ( 
.A(n_4268),
.Y(n_4435)
);

OAI221xp5_ASAP7_75t_L g4436 ( 
.A1(n_4304),
.A2(n_4277),
.B1(n_4253),
.B2(n_4246),
.C(n_4382),
.Y(n_4436)
);

OAI21x1_ASAP7_75t_L g4437 ( 
.A1(n_4368),
.A2(n_4263),
.B(n_4283),
.Y(n_4437)
);

AND2x4_ASAP7_75t_L g4438 ( 
.A(n_4336),
.B(n_4127),
.Y(n_4438)
);

AOI22xp5_ASAP7_75t_L g4439 ( 
.A1(n_4295),
.A2(n_4343),
.B1(n_4313),
.B2(n_4410),
.Y(n_4439)
);

AOI22xp5_ASAP7_75t_L g4440 ( 
.A1(n_4408),
.A2(n_4207),
.B1(n_4014),
.B2(n_4093),
.Y(n_4440)
);

A2O1A1Ixp33_ASAP7_75t_L g4441 ( 
.A1(n_4418),
.A2(n_4137),
.B(n_4210),
.C(n_4214),
.Y(n_4441)
);

AOI21xp33_ASAP7_75t_L g4442 ( 
.A1(n_4397),
.A2(n_4075),
.B(n_4199),
.Y(n_4442)
);

AOI22x1_ASAP7_75t_L g4443 ( 
.A1(n_4369),
.A2(n_4318),
.B1(n_4280),
.B2(n_4404),
.Y(n_4443)
);

AO32x2_ASAP7_75t_L g4444 ( 
.A1(n_4269),
.A2(n_4227),
.A3(n_4163),
.B1(n_4084),
.B2(n_4216),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_4286),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_4290),
.Y(n_4446)
);

INVx2_ASAP7_75t_L g4447 ( 
.A(n_4294),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_4342),
.Y(n_4448)
);

AOI21xp5_ASAP7_75t_SL g4449 ( 
.A1(n_4274),
.A2(n_4362),
.B(n_4256),
.Y(n_4449)
);

NOR2xp33_ASAP7_75t_L g4450 ( 
.A(n_4419),
.B(n_4113),
.Y(n_4450)
);

AND2x4_ASAP7_75t_L g4451 ( 
.A(n_4373),
.B(n_4094),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4417),
.B(n_4100),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_4293),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_4296),
.Y(n_4454)
);

AO31x2_ASAP7_75t_L g4455 ( 
.A1(n_4399),
.A2(n_4043),
.A3(n_4034),
.B(n_4225),
.Y(n_4455)
);

NOR2xp33_ASAP7_75t_L g4456 ( 
.A(n_4302),
.B(n_4117),
.Y(n_4456)
);

BUFx2_ASAP7_75t_L g4457 ( 
.A(n_4267),
.Y(n_4457)
);

INVxp67_ASAP7_75t_L g4458 ( 
.A(n_4358),
.Y(n_4458)
);

AND2x4_ASAP7_75t_L g4459 ( 
.A(n_4312),
.B(n_4094),
.Y(n_4459)
);

INVx2_ASAP7_75t_SL g4460 ( 
.A(n_4309),
.Y(n_4460)
);

OA21x2_ASAP7_75t_L g4461 ( 
.A1(n_4372),
.A2(n_4061),
.B(n_4071),
.Y(n_4461)
);

OAI21x1_ASAP7_75t_L g4462 ( 
.A1(n_4241),
.A2(n_4062),
.B(n_122),
.Y(n_4462)
);

OAI21x1_ASAP7_75t_L g4463 ( 
.A1(n_4351),
.A2(n_124),
.B(n_125),
.Y(n_4463)
);

OAI21x1_ASAP7_75t_L g4464 ( 
.A1(n_4354),
.A2(n_126),
.B(n_127),
.Y(n_4464)
);

O2A1O1Ixp33_ASAP7_75t_L g4465 ( 
.A1(n_4395),
.A2(n_129),
.B(n_127),
.C(n_128),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_4325),
.Y(n_4466)
);

INVxp67_ASAP7_75t_SL g4467 ( 
.A(n_4381),
.Y(n_4467)
);

CKINVDCx20_ASAP7_75t_R g4468 ( 
.A(n_4259),
.Y(n_4468)
);

BUFx3_ASAP7_75t_L g4469 ( 
.A(n_4386),
.Y(n_4469)
);

INVx11_ASAP7_75t_L g4470 ( 
.A(n_4335),
.Y(n_4470)
);

AO31x2_ASAP7_75t_L g4471 ( 
.A1(n_4243),
.A2(n_130),
.A3(n_128),
.B(n_129),
.Y(n_4471)
);

OA21x2_ASAP7_75t_L g4472 ( 
.A1(n_4349),
.A2(n_131),
.B(n_132),
.Y(n_4472)
);

NAND2x1p5_ASAP7_75t_L g4473 ( 
.A(n_4405),
.B(n_542),
.Y(n_4473)
);

OAI21x1_ASAP7_75t_L g4474 ( 
.A1(n_4282),
.A2(n_131),
.B(n_133),
.Y(n_4474)
);

OAI21xp5_ASAP7_75t_SL g4475 ( 
.A1(n_4316),
.A2(n_133),
.B(n_134),
.Y(n_4475)
);

OAI21x1_ASAP7_75t_L g4476 ( 
.A1(n_4273),
.A2(n_134),
.B(n_135),
.Y(n_4476)
);

AOI22xp5_ASAP7_75t_L g4477 ( 
.A1(n_4424),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_4477)
);

OAI21xp5_ASAP7_75t_L g4478 ( 
.A1(n_4376),
.A2(n_136),
.B(n_138),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_4328),
.Y(n_4479)
);

CKINVDCx5p33_ASAP7_75t_R g4480 ( 
.A(n_4366),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4337),
.Y(n_4481)
);

OAI21x1_ASAP7_75t_L g4482 ( 
.A1(n_4402),
.A2(n_138),
.B(n_139),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4339),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_L g4484 ( 
.A(n_4425),
.B(n_543),
.Y(n_4484)
);

OAI21x1_ASAP7_75t_L g4485 ( 
.A1(n_4412),
.A2(n_139),
.B(n_140),
.Y(n_4485)
);

A2O1A1Ixp33_ASAP7_75t_L g4486 ( 
.A1(n_4370),
.A2(n_544),
.B(n_545),
.C(n_543),
.Y(n_4486)
);

INVx2_ASAP7_75t_L g4487 ( 
.A(n_4364),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_4348),
.Y(n_4488)
);

OAI21x1_ASAP7_75t_L g4489 ( 
.A1(n_4276),
.A2(n_140),
.B(n_141),
.Y(n_4489)
);

OR2x2_ASAP7_75t_L g4490 ( 
.A(n_4398),
.B(n_546),
.Y(n_4490)
);

NOR2xp33_ASAP7_75t_L g4491 ( 
.A(n_4255),
.B(n_547),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4350),
.Y(n_4492)
);

OAI22xp5_ASAP7_75t_L g4493 ( 
.A1(n_4247),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_4493)
);

OAI21x1_ASAP7_75t_L g4494 ( 
.A1(n_4401),
.A2(n_142),
.B(n_143),
.Y(n_4494)
);

AOI22xp33_ASAP7_75t_SL g4495 ( 
.A1(n_4271),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_4495)
);

OAI222xp33_ASAP7_75t_L g4496 ( 
.A1(n_4346),
.A2(n_148),
.B1(n_150),
.B2(n_146),
.C1(n_147),
.C2(n_149),
.Y(n_4496)
);

OA21x2_ASAP7_75t_L g4497 ( 
.A1(n_4341),
.A2(n_147),
.B(n_148),
.Y(n_4497)
);

OAI21x1_ASAP7_75t_L g4498 ( 
.A1(n_4384),
.A2(n_149),
.B(n_150),
.Y(n_4498)
);

NOR2x1_ASAP7_75t_R g4499 ( 
.A(n_4421),
.B(n_149),
.Y(n_4499)
);

AND2x4_ASAP7_75t_L g4500 ( 
.A(n_4245),
.B(n_548),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4251),
.Y(n_4501)
);

OAI22xp5_ASAP7_75t_L g4502 ( 
.A1(n_4323),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_4502)
);

HB1xp67_ASAP7_75t_L g4503 ( 
.A(n_4250),
.Y(n_4503)
);

AOI22xp33_ASAP7_75t_L g4504 ( 
.A1(n_4261),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_4504)
);

A2O1A1Ixp33_ASAP7_75t_L g4505 ( 
.A1(n_4428),
.A2(n_551),
.B(n_552),
.C(n_550),
.Y(n_4505)
);

BUFx6f_ASAP7_75t_L g4506 ( 
.A(n_4331),
.Y(n_4506)
);

OAI21x1_ASAP7_75t_L g4507 ( 
.A1(n_4396),
.A2(n_152),
.B(n_153),
.Y(n_4507)
);

OAI21xp5_ASAP7_75t_L g4508 ( 
.A1(n_4422),
.A2(n_154),
.B(n_155),
.Y(n_4508)
);

OAI21x1_ASAP7_75t_L g4509 ( 
.A1(n_4264),
.A2(n_154),
.B(n_155),
.Y(n_4509)
);

AOI21x1_ASAP7_75t_L g4510 ( 
.A1(n_4406),
.A2(n_155),
.B(n_156),
.Y(n_4510)
);

CKINVDCx5p33_ASAP7_75t_R g4511 ( 
.A(n_4391),
.Y(n_4511)
);

OAI21x1_ASAP7_75t_L g4512 ( 
.A1(n_4281),
.A2(n_156),
.B(n_157),
.Y(n_4512)
);

INVx2_ASAP7_75t_SL g4513 ( 
.A(n_4400),
.Y(n_4513)
);

INVx2_ASAP7_75t_L g4514 ( 
.A(n_4260),
.Y(n_4514)
);

AND2x4_ASAP7_75t_L g4515 ( 
.A(n_4420),
.B(n_551),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4262),
.Y(n_4516)
);

OAI21x1_ASAP7_75t_L g4517 ( 
.A1(n_4344),
.A2(n_156),
.B(n_157),
.Y(n_4517)
);

AND2x4_ASAP7_75t_L g4518 ( 
.A(n_4311),
.B(n_552),
.Y(n_4518)
);

BUFx3_ASAP7_75t_L g4519 ( 
.A(n_4266),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4272),
.Y(n_4520)
);

INVx2_ASAP7_75t_L g4521 ( 
.A(n_4279),
.Y(n_4521)
);

INVxp67_ASAP7_75t_L g4522 ( 
.A(n_4330),
.Y(n_4522)
);

OA21x2_ASAP7_75t_L g4523 ( 
.A1(n_4367),
.A2(n_157),
.B(n_158),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4359),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_4361),
.Y(n_4525)
);

AOI221xp5_ASAP7_75t_L g4526 ( 
.A1(n_4423),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.C(n_162),
.Y(n_4526)
);

OA21x2_ASAP7_75t_L g4527 ( 
.A1(n_4356),
.A2(n_160),
.B(n_162),
.Y(n_4527)
);

INVx2_ASAP7_75t_SL g4528 ( 
.A(n_4278),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4244),
.Y(n_4529)
);

BUFx6f_ASAP7_75t_L g4530 ( 
.A(n_4409),
.Y(n_4530)
);

AO21x2_ASAP7_75t_L g4531 ( 
.A1(n_4314),
.A2(n_163),
.B(n_164),
.Y(n_4531)
);

INVx2_ASAP7_75t_SL g4532 ( 
.A(n_4275),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4413),
.Y(n_4533)
);

INVx2_ASAP7_75t_SL g4534 ( 
.A(n_4329),
.Y(n_4534)
);

INVxp67_ASAP7_75t_L g4535 ( 
.A(n_4392),
.Y(n_4535)
);

OAI21x1_ASAP7_75t_L g4536 ( 
.A1(n_4326),
.A2(n_163),
.B(n_164),
.Y(n_4536)
);

INVxp67_ASAP7_75t_SL g4537 ( 
.A(n_4248),
.Y(n_4537)
);

OAI22xp5_ASAP7_75t_L g4538 ( 
.A1(n_4270),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_4538)
);

OR2x6_ASAP7_75t_L g4539 ( 
.A(n_4429),
.B(n_554),
.Y(n_4539)
);

AOI21xp5_ASAP7_75t_L g4540 ( 
.A1(n_4379),
.A2(n_555),
.B(n_554),
.Y(n_4540)
);

AND2x4_ASAP7_75t_L g4541 ( 
.A(n_4288),
.B(n_4416),
.Y(n_4541)
);

AO21x2_ASAP7_75t_L g4542 ( 
.A1(n_4347),
.A2(n_165),
.B(n_166),
.Y(n_4542)
);

OAI22xp33_ASAP7_75t_L g4543 ( 
.A1(n_4297),
.A2(n_557),
.B1(n_558),
.B2(n_556),
.Y(n_4543)
);

OAI21xp5_ASAP7_75t_L g4544 ( 
.A1(n_4407),
.A2(n_166),
.B(n_167),
.Y(n_4544)
);

AO21x2_ASAP7_75t_L g4545 ( 
.A1(n_4292),
.A2(n_167),
.B(n_168),
.Y(n_4545)
);

NAND2x1p5_ASAP7_75t_L g4546 ( 
.A(n_4355),
.B(n_556),
.Y(n_4546)
);

OR2x6_ASAP7_75t_L g4547 ( 
.A(n_4258),
.B(n_4403),
.Y(n_4547)
);

BUFx2_ASAP7_75t_L g4548 ( 
.A(n_4335),
.Y(n_4548)
);

INVx2_ASAP7_75t_L g4549 ( 
.A(n_4415),
.Y(n_4549)
);

OAI21x1_ASAP7_75t_L g4550 ( 
.A1(n_4371),
.A2(n_167),
.B(n_168),
.Y(n_4550)
);

OAI21xp5_ASAP7_75t_L g4551 ( 
.A1(n_4363),
.A2(n_4285),
.B(n_4383),
.Y(n_4551)
);

INVxp67_ASAP7_75t_SL g4552 ( 
.A(n_4389),
.Y(n_4552)
);

BUFx2_ASAP7_75t_L g4553 ( 
.A(n_4335),
.Y(n_4553)
);

INVx2_ASAP7_75t_L g4554 ( 
.A(n_4514),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4445),
.Y(n_4555)
);

AOI21x1_ASAP7_75t_L g4556 ( 
.A1(n_4510),
.A2(n_4345),
.B(n_4387),
.Y(n_4556)
);

AOI21x1_ASAP7_75t_L g4557 ( 
.A1(n_4529),
.A2(n_4345),
.B(n_4388),
.Y(n_4557)
);

OA21x2_ASAP7_75t_L g4558 ( 
.A1(n_4494),
.A2(n_4426),
.B(n_4303),
.Y(n_4558)
);

HB1xp67_ASAP7_75t_L g4559 ( 
.A(n_4467),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_4446),
.Y(n_4560)
);

AOI21xp5_ASAP7_75t_L g4561 ( 
.A1(n_4441),
.A2(n_4284),
.B(n_4307),
.Y(n_4561)
);

AOI21xp5_ASAP7_75t_L g4562 ( 
.A1(n_4442),
.A2(n_4393),
.B(n_4257),
.Y(n_4562)
);

AOI21xp5_ASAP7_75t_L g4563 ( 
.A1(n_4551),
.A2(n_4411),
.B(n_4334),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_L g4564 ( 
.A(n_4537),
.B(n_4242),
.Y(n_4564)
);

A2O1A1Ixp33_ASAP7_75t_L g4565 ( 
.A1(n_4436),
.A2(n_4377),
.B(n_4324),
.C(n_4390),
.Y(n_4565)
);

A2O1A1Ixp33_ASAP7_75t_L g4566 ( 
.A1(n_4478),
.A2(n_4414),
.B(n_4375),
.C(n_4380),
.Y(n_4566)
);

INVx1_ASAP7_75t_L g4567 ( 
.A(n_4453),
.Y(n_4567)
);

OAI21x1_ASAP7_75t_L g4568 ( 
.A1(n_4437),
.A2(n_4291),
.B(n_4289),
.Y(n_4568)
);

CKINVDCx8_ASAP7_75t_R g4569 ( 
.A(n_4480),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4454),
.Y(n_4570)
);

AOI21x1_ASAP7_75t_L g4571 ( 
.A1(n_4540),
.A2(n_4365),
.B(n_4320),
.Y(n_4571)
);

OAI22xp5_ASAP7_75t_SL g4572 ( 
.A1(n_4511),
.A2(n_4403),
.B1(n_4258),
.B2(n_4315),
.Y(n_4572)
);

NAND2xp5_ASAP7_75t_L g4573 ( 
.A(n_4535),
.B(n_4252),
.Y(n_4573)
);

NAND2xp5_ASAP7_75t_L g4574 ( 
.A(n_4503),
.B(n_4299),
.Y(n_4574)
);

AO31x2_ASAP7_75t_L g4575 ( 
.A1(n_4549),
.A2(n_4385),
.A3(n_4321),
.B(n_4322),
.Y(n_4575)
);

INVx2_ASAP7_75t_L g4576 ( 
.A(n_4521),
.Y(n_4576)
);

AOI21xp5_ASAP7_75t_L g4577 ( 
.A1(n_4433),
.A2(n_4338),
.B(n_4333),
.Y(n_4577)
);

OAI21x1_ASAP7_75t_L g4578 ( 
.A1(n_4434),
.A2(n_4301),
.B(n_4298),
.Y(n_4578)
);

AO21x2_ASAP7_75t_L g4579 ( 
.A1(n_4531),
.A2(n_4327),
.B(n_4319),
.Y(n_4579)
);

OA21x2_ASAP7_75t_L g4580 ( 
.A1(n_4462),
.A2(n_4394),
.B(n_4340),
.Y(n_4580)
);

OA21x2_ASAP7_75t_L g4581 ( 
.A1(n_4463),
.A2(n_4287),
.B(n_4305),
.Y(n_4581)
);

INVx2_ASAP7_75t_L g4582 ( 
.A(n_4501),
.Y(n_4582)
);

CKINVDCx11_ASAP7_75t_R g4583 ( 
.A(n_4468),
.Y(n_4583)
);

NAND2xp5_ASAP7_75t_L g4584 ( 
.A(n_4458),
.B(n_4332),
.Y(n_4584)
);

INVx6_ASAP7_75t_L g4585 ( 
.A(n_4506),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4466),
.Y(n_4586)
);

AO21x2_ASAP7_75t_L g4587 ( 
.A1(n_4552),
.A2(n_4300),
.B(n_4308),
.Y(n_4587)
);

INVx2_ASAP7_75t_L g4588 ( 
.A(n_4516),
.Y(n_4588)
);

OAI21xp5_ASAP7_75t_L g4589 ( 
.A1(n_4544),
.A2(n_4306),
.B(n_4378),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4479),
.Y(n_4590)
);

INVx2_ASAP7_75t_SL g4591 ( 
.A(n_4430),
.Y(n_4591)
);

INVx2_ASAP7_75t_L g4592 ( 
.A(n_4520),
.Y(n_4592)
);

BUFx2_ASAP7_75t_R g4593 ( 
.A(n_4431),
.Y(n_4593)
);

AND2x4_ASAP7_75t_L g4594 ( 
.A(n_4457),
.B(n_4249),
.Y(n_4594)
);

AND2x2_ASAP7_75t_L g4595 ( 
.A(n_4481),
.B(n_4427),
.Y(n_4595)
);

OAI21xp5_ASAP7_75t_L g4596 ( 
.A1(n_4505),
.A2(n_4357),
.B(n_4310),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4483),
.Y(n_4597)
);

OA21x2_ASAP7_75t_L g4598 ( 
.A1(n_4464),
.A2(n_4352),
.B(n_4353),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4488),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4492),
.Y(n_4600)
);

A2O1A1Ixp33_ASAP7_75t_L g4601 ( 
.A1(n_4439),
.A2(n_4475),
.B(n_4508),
.C(n_4465),
.Y(n_4601)
);

BUFx3_ASAP7_75t_L g4602 ( 
.A(n_4469),
.Y(n_4602)
);

BUFx6f_ASAP7_75t_L g4603 ( 
.A(n_4451),
.Y(n_4603)
);

NAND2xp5_ASAP7_75t_L g4604 ( 
.A(n_4522),
.B(n_557),
.Y(n_4604)
);

BUFx6f_ASAP7_75t_L g4605 ( 
.A(n_4459),
.Y(n_4605)
);

AOI22xp33_ASAP7_75t_SL g4606 ( 
.A1(n_4443),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_4606)
);

OAI21xp5_ASAP7_75t_L g4607 ( 
.A1(n_4486),
.A2(n_171),
.B(n_172),
.Y(n_4607)
);

AOI22xp5_ASAP7_75t_L g4608 ( 
.A1(n_4539),
.A2(n_174),
.B1(n_171),
.B2(n_173),
.Y(n_4608)
);

OAI21xp5_ASAP7_75t_L g4609 ( 
.A1(n_4449),
.A2(n_173),
.B(n_174),
.Y(n_4609)
);

INVx2_ASAP7_75t_L g4610 ( 
.A(n_4524),
.Y(n_4610)
);

BUFx2_ASAP7_75t_L g4611 ( 
.A(n_4548),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4525),
.Y(n_4612)
);

NAND2x1p5_ASAP7_75t_L g4613 ( 
.A(n_4553),
.B(n_558),
.Y(n_4613)
);

AO31x2_ASAP7_75t_L g4614 ( 
.A1(n_4538),
.A2(n_177),
.A3(n_175),
.B(n_176),
.Y(n_4614)
);

NAND2xp5_ASAP7_75t_L g4615 ( 
.A(n_4452),
.B(n_559),
.Y(n_4615)
);

OR2x2_ASAP7_75t_L g4616 ( 
.A(n_4490),
.B(n_559),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4435),
.Y(n_4617)
);

AOI21xp5_ASAP7_75t_L g4618 ( 
.A1(n_4539),
.A2(n_176),
.B(n_177),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4447),
.Y(n_4619)
);

AO31x2_ASAP7_75t_L g4620 ( 
.A1(n_4493),
.A2(n_180),
.A3(n_178),
.B(n_179),
.Y(n_4620)
);

OAI21x1_ASAP7_75t_L g4621 ( 
.A1(n_4482),
.A2(n_179),
.B(n_180),
.Y(n_4621)
);

AND2x2_ASAP7_75t_L g4622 ( 
.A(n_4456),
.B(n_560),
.Y(n_4622)
);

OAI21x1_ASAP7_75t_L g4623 ( 
.A1(n_4485),
.A2(n_179),
.B(n_180),
.Y(n_4623)
);

OAI21x1_ASAP7_75t_SL g4624 ( 
.A1(n_4526),
.A2(n_4461),
.B(n_4440),
.Y(n_4624)
);

INVx3_ASAP7_75t_L g4625 ( 
.A(n_4530),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4448),
.B(n_561),
.Y(n_4626)
);

AOI21xp5_ASAP7_75t_L g4627 ( 
.A1(n_4527),
.A2(n_181),
.B(n_182),
.Y(n_4627)
);

NAND2xp5_ASAP7_75t_SL g4628 ( 
.A(n_4541),
.B(n_561),
.Y(n_4628)
);

OAI21xp5_ASAP7_75t_L g4629 ( 
.A1(n_4509),
.A2(n_181),
.B(n_182),
.Y(n_4629)
);

AOI21x1_ASAP7_75t_L g4630 ( 
.A1(n_4474),
.A2(n_183),
.B(n_184),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_L g4631 ( 
.A(n_4487),
.B(n_562),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4533),
.Y(n_4632)
);

OAI21x1_ASAP7_75t_L g4633 ( 
.A1(n_4476),
.A2(n_184),
.B(n_185),
.Y(n_4633)
);

INVxp67_ASAP7_75t_L g4634 ( 
.A(n_4513),
.Y(n_4634)
);

AO31x2_ASAP7_75t_L g4635 ( 
.A1(n_4502),
.A2(n_188),
.A3(n_186),
.B(n_187),
.Y(n_4635)
);

NOR2x1_ASAP7_75t_SL g4636 ( 
.A(n_4545),
.B(n_562),
.Y(n_4636)
);

OAI21xp5_ASAP7_75t_L g4637 ( 
.A1(n_4495),
.A2(n_4517),
.B(n_4543),
.Y(n_4637)
);

NOR2xp33_ASAP7_75t_L g4638 ( 
.A(n_4450),
.B(n_564),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_4484),
.B(n_565),
.Y(n_4639)
);

OA21x2_ASAP7_75t_L g4640 ( 
.A1(n_4550),
.A2(n_4512),
.B(n_4489),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4455),
.Y(n_4641)
);

NAND2x1p5_ASAP7_75t_L g4642 ( 
.A(n_4438),
.B(n_567),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4498),
.Y(n_4643)
);

BUFx12f_ASAP7_75t_L g4644 ( 
.A(n_4500),
.Y(n_4644)
);

INVx1_ASAP7_75t_SL g4645 ( 
.A(n_4519),
.Y(n_4645)
);

AOI21xp5_ASAP7_75t_L g4646 ( 
.A1(n_4497),
.A2(n_191),
.B(n_192),
.Y(n_4646)
);

CKINVDCx8_ASAP7_75t_R g4647 ( 
.A(n_4547),
.Y(n_4647)
);

AOI21xp5_ASAP7_75t_L g4648 ( 
.A1(n_4523),
.A2(n_192),
.B(n_193),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4507),
.Y(n_4649)
);

INVx1_ASAP7_75t_L g4650 ( 
.A(n_4471),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4491),
.B(n_569),
.Y(n_4651)
);

OR2x2_ASAP7_75t_L g4652 ( 
.A(n_4542),
.B(n_570),
.Y(n_4652)
);

NAND2xp5_ASAP7_75t_L g4653 ( 
.A(n_4515),
.B(n_570),
.Y(n_4653)
);

OAI21x1_ASAP7_75t_L g4654 ( 
.A1(n_4536),
.A2(n_194),
.B(n_195),
.Y(n_4654)
);

NAND2xp5_ASAP7_75t_L g4655 ( 
.A(n_4477),
.B(n_571),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4471),
.Y(n_4656)
);

OAI21x1_ASAP7_75t_L g4657 ( 
.A1(n_4472),
.A2(n_196),
.B(n_197),
.Y(n_4657)
);

OA21x2_ASAP7_75t_L g4658 ( 
.A1(n_4496),
.A2(n_196),
.B(n_198),
.Y(n_4658)
);

NAND2xp5_ASAP7_75t_L g4659 ( 
.A(n_4546),
.B(n_572),
.Y(n_4659)
);

AOI21x1_ASAP7_75t_L g4660 ( 
.A1(n_4432),
.A2(n_198),
.B(n_199),
.Y(n_4660)
);

AND2x2_ASAP7_75t_L g4661 ( 
.A(n_4532),
.B(n_573),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_4473),
.B(n_573),
.Y(n_4662)
);

INVx2_ASAP7_75t_L g4663 ( 
.A(n_4460),
.Y(n_4663)
);

AND2x2_ASAP7_75t_L g4664 ( 
.A(n_4611),
.B(n_4534),
.Y(n_4664)
);

INVx2_ASAP7_75t_L g4665 ( 
.A(n_4582),
.Y(n_4665)
);

INVx1_ASAP7_75t_L g4666 ( 
.A(n_4555),
.Y(n_4666)
);

INVx1_ASAP7_75t_L g4667 ( 
.A(n_4560),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4567),
.Y(n_4668)
);

AO21x2_ASAP7_75t_L g4669 ( 
.A1(n_4577),
.A2(n_4518),
.B(n_4470),
.Y(n_4669)
);

INVxp67_ASAP7_75t_L g4670 ( 
.A(n_4574),
.Y(n_4670)
);

INVx2_ASAP7_75t_L g4671 ( 
.A(n_4588),
.Y(n_4671)
);

INVx2_ASAP7_75t_L g4672 ( 
.A(n_4592),
.Y(n_4672)
);

BUFx3_ASAP7_75t_L g4673 ( 
.A(n_4602),
.Y(n_4673)
);

OA21x2_ASAP7_75t_L g4674 ( 
.A1(n_4568),
.A2(n_4504),
.B(n_4528),
.Y(n_4674)
);

HB1xp67_ASAP7_75t_L g4675 ( 
.A(n_4594),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4570),
.Y(n_4676)
);

OAI321xp33_ASAP7_75t_L g4677 ( 
.A1(n_4609),
.A2(n_4444),
.A3(n_4499),
.B1(n_202),
.B2(n_205),
.C(n_200),
.Y(n_4677)
);

HB1xp67_ASAP7_75t_L g4678 ( 
.A(n_4554),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_4586),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_4610),
.Y(n_4680)
);

CKINVDCx6p67_ASAP7_75t_R g4681 ( 
.A(n_4583),
.Y(n_4681)
);

HB1xp67_ASAP7_75t_L g4682 ( 
.A(n_4576),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_4590),
.Y(n_4683)
);

INVx2_ASAP7_75t_L g4684 ( 
.A(n_4597),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4599),
.Y(n_4685)
);

INVx2_ASAP7_75t_L g4686 ( 
.A(n_4600),
.Y(n_4686)
);

HB1xp67_ASAP7_75t_L g4687 ( 
.A(n_4612),
.Y(n_4687)
);

INVx3_ASAP7_75t_L g4688 ( 
.A(n_4603),
.Y(n_4688)
);

INVx2_ASAP7_75t_L g4689 ( 
.A(n_4617),
.Y(n_4689)
);

AND2x4_ASAP7_75t_L g4690 ( 
.A(n_4619),
.B(n_576),
.Y(n_4690)
);

AND2x2_ASAP7_75t_L g4691 ( 
.A(n_4595),
.B(n_576),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4650),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4656),
.Y(n_4693)
);

NAND2xp5_ASAP7_75t_L g4694 ( 
.A(n_4573),
.B(n_577),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4632),
.Y(n_4695)
);

OR2x2_ASAP7_75t_L g4696 ( 
.A(n_4575),
.B(n_578),
.Y(n_4696)
);

NOR2xp33_ASAP7_75t_L g4697 ( 
.A(n_4647),
.B(n_579),
.Y(n_4697)
);

INVx2_ASAP7_75t_SL g4698 ( 
.A(n_4591),
.Y(n_4698)
);

AND2x2_ASAP7_75t_L g4699 ( 
.A(n_4663),
.B(n_4622),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4641),
.Y(n_4700)
);

CKINVDCx11_ASAP7_75t_R g4701 ( 
.A(n_4569),
.Y(n_4701)
);

NAND2xp5_ASAP7_75t_L g4702 ( 
.A(n_4579),
.B(n_579),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4643),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4649),
.Y(n_4704)
);

OR2x2_ASAP7_75t_L g4705 ( 
.A(n_4580),
.B(n_4616),
.Y(n_4705)
);

INVx1_ASAP7_75t_L g4706 ( 
.A(n_4557),
.Y(n_4706)
);

CKINVDCx20_ASAP7_75t_R g4707 ( 
.A(n_4605),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4626),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4631),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_4657),
.Y(n_4710)
);

BUFx3_ASAP7_75t_L g4711 ( 
.A(n_4585),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4640),
.Y(n_4712)
);

AND2x2_ASAP7_75t_L g4713 ( 
.A(n_4634),
.B(n_581),
.Y(n_4713)
);

OAI21xp33_ASAP7_75t_SL g4714 ( 
.A1(n_4652),
.A2(n_4607),
.B(n_4589),
.Y(n_4714)
);

NAND2xp5_ASAP7_75t_L g4715 ( 
.A(n_4563),
.B(n_581),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_4578),
.Y(n_4716)
);

INVx2_ASAP7_75t_L g4717 ( 
.A(n_4587),
.Y(n_4717)
);

AND2x2_ASAP7_75t_L g4718 ( 
.A(n_4625),
.B(n_582),
.Y(n_4718)
);

AO21x2_ASAP7_75t_L g4719 ( 
.A1(n_4646),
.A2(n_201),
.B(n_204),
.Y(n_4719)
);

INVx2_ASAP7_75t_L g4720 ( 
.A(n_4581),
.Y(n_4720)
);

OR2x2_ASAP7_75t_L g4721 ( 
.A(n_4584),
.B(n_583),
.Y(n_4721)
);

INVx1_ASAP7_75t_SL g4722 ( 
.A(n_4593),
.Y(n_4722)
);

INVx2_ASAP7_75t_L g4723 ( 
.A(n_4556),
.Y(n_4723)
);

AND2x2_ASAP7_75t_L g4724 ( 
.A(n_4605),
.B(n_584),
.Y(n_4724)
);

BUFx2_ASAP7_75t_L g4725 ( 
.A(n_4644),
.Y(n_4725)
);

BUFx6f_ASAP7_75t_L g4726 ( 
.A(n_4661),
.Y(n_4726)
);

INVx2_ASAP7_75t_L g4727 ( 
.A(n_4615),
.Y(n_4727)
);

HB1xp67_ASAP7_75t_L g4728 ( 
.A(n_4558),
.Y(n_4728)
);

INVx2_ASAP7_75t_L g4729 ( 
.A(n_4636),
.Y(n_4729)
);

BUFx3_ASAP7_75t_L g4730 ( 
.A(n_4642),
.Y(n_4730)
);

INVx1_ASAP7_75t_L g4731 ( 
.A(n_4630),
.Y(n_4731)
);

AOI22xp33_ASAP7_75t_L g4732 ( 
.A1(n_4637),
.A2(n_4572),
.B1(n_4624),
.B2(n_4596),
.Y(n_4732)
);

INVx2_ASAP7_75t_L g4733 ( 
.A(n_4660),
.Y(n_4733)
);

INVx1_ASAP7_75t_L g4734 ( 
.A(n_4598),
.Y(n_4734)
);

INVx1_ASAP7_75t_L g4735 ( 
.A(n_4621),
.Y(n_4735)
);

INVx3_ASAP7_75t_L g4736 ( 
.A(n_4613),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4623),
.Y(n_4737)
);

AND2x2_ASAP7_75t_L g4738 ( 
.A(n_4638),
.B(n_585),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4654),
.Y(n_4739)
);

AND2x4_ASAP7_75t_L g4740 ( 
.A(n_4571),
.B(n_586),
.Y(n_4740)
);

OA21x2_ASAP7_75t_L g4741 ( 
.A1(n_4648),
.A2(n_588),
.B(n_587),
.Y(n_4741)
);

INVx2_ASAP7_75t_L g4742 ( 
.A(n_4633),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_4604),
.Y(n_4743)
);

OAI21xp5_ASAP7_75t_L g4744 ( 
.A1(n_4562),
.A2(n_201),
.B(n_204),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4566),
.B(n_4639),
.Y(n_4745)
);

BUFx3_ASAP7_75t_L g4746 ( 
.A(n_4653),
.Y(n_4746)
);

OA21x2_ASAP7_75t_L g4747 ( 
.A1(n_4627),
.A2(n_589),
.B(n_588),
.Y(n_4747)
);

OR2x2_ASAP7_75t_L g4748 ( 
.A(n_4651),
.B(n_589),
.Y(n_4748)
);

INVx3_ASAP7_75t_L g4749 ( 
.A(n_4620),
.Y(n_4749)
);

BUFx6f_ASAP7_75t_L g4750 ( 
.A(n_4628),
.Y(n_4750)
);

AND2x4_ASAP7_75t_SL g4751 ( 
.A(n_4608),
.B(n_590),
.Y(n_4751)
);

AND2x2_ASAP7_75t_L g4752 ( 
.A(n_4662),
.B(n_4659),
.Y(n_4752)
);

AND2x2_ASAP7_75t_L g4753 ( 
.A(n_4629),
.B(n_591),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4635),
.Y(n_4754)
);

INVx1_ASAP7_75t_L g4755 ( 
.A(n_4635),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4614),
.Y(n_4756)
);

INVx1_ASAP7_75t_L g4757 ( 
.A(n_4614),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_4561),
.Y(n_4758)
);

AND2x2_ASAP7_75t_L g4759 ( 
.A(n_4618),
.B(n_593),
.Y(n_4759)
);

HB1xp67_ASAP7_75t_L g4760 ( 
.A(n_4655),
.Y(n_4760)
);

INVx4_ASAP7_75t_L g4761 ( 
.A(n_4658),
.Y(n_4761)
);

INVx3_ASAP7_75t_L g4762 ( 
.A(n_4565),
.Y(n_4762)
);

INVx3_ASAP7_75t_L g4763 ( 
.A(n_4601),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4606),
.Y(n_4764)
);

AO21x1_ASAP7_75t_SL g4765 ( 
.A1(n_4564),
.A2(n_205),
.B(n_206),
.Y(n_4765)
);

AO21x2_ASAP7_75t_L g4766 ( 
.A1(n_4577),
.A2(n_206),
.B(n_207),
.Y(n_4766)
);

CKINVDCx5p33_ASAP7_75t_R g4767 ( 
.A(n_4583),
.Y(n_4767)
);

INVx2_ASAP7_75t_L g4768 ( 
.A(n_4582),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4555),
.Y(n_4769)
);

INVx2_ASAP7_75t_L g4770 ( 
.A(n_4582),
.Y(n_4770)
);

BUFx3_ASAP7_75t_L g4771 ( 
.A(n_4602),
.Y(n_4771)
);

INVx3_ASAP7_75t_L g4772 ( 
.A(n_4602),
.Y(n_4772)
);

INVx1_ASAP7_75t_SL g4773 ( 
.A(n_4645),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4555),
.Y(n_4774)
);

INVx1_ASAP7_75t_L g4775 ( 
.A(n_4555),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4555),
.Y(n_4776)
);

HB1xp67_ASAP7_75t_L g4777 ( 
.A(n_4559),
.Y(n_4777)
);

INVx3_ASAP7_75t_L g4778 ( 
.A(n_4602),
.Y(n_4778)
);

OR2x2_ASAP7_75t_L g4779 ( 
.A(n_4777),
.B(n_207),
.Y(n_4779)
);

NAND2xp5_ASAP7_75t_L g4780 ( 
.A(n_4670),
.B(n_596),
.Y(n_4780)
);

OAI21x1_ASAP7_75t_L g4781 ( 
.A1(n_4723),
.A2(n_207),
.B(n_208),
.Y(n_4781)
);

OAI21x1_ASAP7_75t_L g4782 ( 
.A1(n_4717),
.A2(n_208),
.B(n_209),
.Y(n_4782)
);

INVx2_ASAP7_75t_L g4783 ( 
.A(n_4684),
.Y(n_4783)
);

OAI221xp5_ASAP7_75t_L g4784 ( 
.A1(n_4714),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.C(n_213),
.Y(n_4784)
);

AOI22xp33_ASAP7_75t_L g4785 ( 
.A1(n_4732),
.A2(n_598),
.B1(n_599),
.B2(n_597),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4705),
.B(n_597),
.Y(n_4786)
);

AOI222xp33_ASAP7_75t_L g4787 ( 
.A1(n_4744),
.A2(n_214),
.B1(n_216),
.B2(n_210),
.C1(n_211),
.C2(n_215),
.Y(n_4787)
);

OAI22xp5_ASAP7_75t_L g4788 ( 
.A1(n_4762),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_4788)
);

OAI22xp33_ASAP7_75t_L g4789 ( 
.A1(n_4677),
.A2(n_599),
.B1(n_600),
.B2(n_598),
.Y(n_4789)
);

A2O1A1Ixp33_ASAP7_75t_L g4790 ( 
.A1(n_4715),
.A2(n_603),
.B(n_604),
.C(n_602),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4687),
.Y(n_4791)
);

OA21x2_ASAP7_75t_L g4792 ( 
.A1(n_4734),
.A2(n_217),
.B(n_218),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4686),
.Y(n_4793)
);

AOI221xp5_ASAP7_75t_L g4794 ( 
.A1(n_4745),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.C(n_220),
.Y(n_4794)
);

OAI22xp5_ASAP7_75t_L g4795 ( 
.A1(n_4764),
.A2(n_221),
.B1(n_218),
.B2(n_220),
.Y(n_4795)
);

OAI21xp5_ASAP7_75t_L g4796 ( 
.A1(n_4702),
.A2(n_607),
.B(n_605),
.Y(n_4796)
);

AND2x2_ASAP7_75t_L g4797 ( 
.A(n_4678),
.B(n_221),
.Y(n_4797)
);

OAI22xp33_ASAP7_75t_L g4798 ( 
.A1(n_4761),
.A2(n_609),
.B1(n_613),
.B2(n_608),
.Y(n_4798)
);

OAI221xp5_ASAP7_75t_SL g4799 ( 
.A1(n_4753),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.C(n_224),
.Y(n_4799)
);

AND2x4_ASAP7_75t_L g4800 ( 
.A(n_4664),
.B(n_609),
.Y(n_4800)
);

OAI22xp5_ASAP7_75t_SL g4801 ( 
.A1(n_4722),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_4801)
);

AND2x2_ASAP7_75t_L g4802 ( 
.A(n_4682),
.B(n_225),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_L g4803 ( 
.A(n_4727),
.B(n_614),
.Y(n_4803)
);

OAI211xp5_ASAP7_75t_SL g4804 ( 
.A1(n_4708),
.A2(n_228),
.B(n_226),
.C(n_227),
.Y(n_4804)
);

AOI222xp33_ASAP7_75t_L g4805 ( 
.A1(n_4751),
.A2(n_230),
.B1(n_232),
.B2(n_228),
.C1(n_229),
.C2(n_231),
.Y(n_4805)
);

NAND2xp5_ASAP7_75t_L g4806 ( 
.A(n_4709),
.B(n_614),
.Y(n_4806)
);

OAI211xp5_ASAP7_75t_L g4807 ( 
.A1(n_4759),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_4807)
);

BUFx6f_ASAP7_75t_L g4808 ( 
.A(n_4701),
.Y(n_4808)
);

INVx2_ASAP7_75t_L g4809 ( 
.A(n_4666),
.Y(n_4809)
);

INVx4_ASAP7_75t_L g4810 ( 
.A(n_4767),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4667),
.Y(n_4811)
);

BUFx3_ASAP7_75t_L g4812 ( 
.A(n_4681),
.Y(n_4812)
);

NAND3xp33_ASAP7_75t_L g4813 ( 
.A(n_4758),
.B(n_616),
.C(n_615),
.Y(n_4813)
);

INVx1_ASAP7_75t_L g4814 ( 
.A(n_4668),
.Y(n_4814)
);

OAI221xp5_ASAP7_75t_L g4815 ( 
.A1(n_4729),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.C(n_236),
.Y(n_4815)
);

INVx2_ASAP7_75t_L g4816 ( 
.A(n_4676),
.Y(n_4816)
);

OR2x2_ASAP7_75t_L g4817 ( 
.A(n_4703),
.B(n_233),
.Y(n_4817)
);

AND2x2_ASAP7_75t_L g4818 ( 
.A(n_4699),
.B(n_234),
.Y(n_4818)
);

AOI22xp33_ASAP7_75t_L g4819 ( 
.A1(n_4750),
.A2(n_619),
.B1(n_620),
.B2(n_618),
.Y(n_4819)
);

AOI22xp33_ASAP7_75t_L g4820 ( 
.A1(n_4719),
.A2(n_622),
.B1(n_623),
.B2(n_621),
.Y(n_4820)
);

AOI22xp33_ASAP7_75t_L g4821 ( 
.A1(n_4760),
.A2(n_623),
.B1(n_624),
.B2(n_621),
.Y(n_4821)
);

AOI22xp33_ASAP7_75t_L g4822 ( 
.A1(n_4766),
.A2(n_625),
.B1(n_626),
.B2(n_624),
.Y(n_4822)
);

AO221x1_ASAP7_75t_L g4823 ( 
.A1(n_4749),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.C(n_239),
.Y(n_4823)
);

AOI21xp33_ASAP7_75t_L g4824 ( 
.A1(n_4669),
.A2(n_627),
.B(n_626),
.Y(n_4824)
);

OAI211xp5_ASAP7_75t_L g4825 ( 
.A1(n_4754),
.A2(n_243),
.B(n_241),
.C(n_242),
.Y(n_4825)
);

BUFx5_ASAP7_75t_L g4826 ( 
.A(n_4712),
.Y(n_4826)
);

INVx1_ASAP7_75t_L g4827 ( 
.A(n_4679),
.Y(n_4827)
);

NAND2xp5_ASAP7_75t_L g4828 ( 
.A(n_4743),
.B(n_627),
.Y(n_4828)
);

OAI221xp5_ASAP7_75t_L g4829 ( 
.A1(n_4721),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.C(n_245),
.Y(n_4829)
);

INVx2_ASAP7_75t_L g4830 ( 
.A(n_4683),
.Y(n_4830)
);

OAI22xp5_ASAP7_75t_SL g4831 ( 
.A1(n_4707),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_4831)
);

HB1xp67_ASAP7_75t_L g4832 ( 
.A(n_4728),
.Y(n_4832)
);

AOI22xp33_ASAP7_75t_L g4833 ( 
.A1(n_4752),
.A2(n_630),
.B1(n_631),
.B2(n_629),
.Y(n_4833)
);

NAND2xp5_ASAP7_75t_L g4834 ( 
.A(n_4689),
.B(n_629),
.Y(n_4834)
);

INVx1_ASAP7_75t_L g4835 ( 
.A(n_4685),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_L g4836 ( 
.A(n_4695),
.B(n_630),
.Y(n_4836)
);

BUFx3_ASAP7_75t_L g4837 ( 
.A(n_4673),
.Y(n_4837)
);

AO21x2_ASAP7_75t_L g4838 ( 
.A1(n_4706),
.A2(n_246),
.B(n_247),
.Y(n_4838)
);

OAI22xp5_ASAP7_75t_L g4839 ( 
.A1(n_4736),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_4839)
);

OAI332xp33_ASAP7_75t_L g4840 ( 
.A1(n_4755),
.A2(n_251),
.A3(n_250),
.B1(n_248),
.B2(n_252),
.B3(n_246),
.C1(n_247),
.C2(n_249),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_4769),
.Y(n_4841)
);

OAI21x1_ASAP7_75t_L g4842 ( 
.A1(n_4716),
.A2(n_249),
.B(n_250),
.Y(n_4842)
);

AOI221xp5_ASAP7_75t_SL g4843 ( 
.A1(n_4756),
.A2(n_4757),
.B1(n_4697),
.B2(n_4694),
.C(n_4738),
.Y(n_4843)
);

OR2x2_ASAP7_75t_L g4844 ( 
.A(n_4704),
.B(n_249),
.Y(n_4844)
);

INVx2_ASAP7_75t_L g4845 ( 
.A(n_4774),
.Y(n_4845)
);

AOI22xp33_ASAP7_75t_L g4846 ( 
.A1(n_4740),
.A2(n_633),
.B1(n_634),
.B2(n_632),
.Y(n_4846)
);

NOR2x1_ASAP7_75t_SL g4847 ( 
.A(n_4696),
.B(n_4765),
.Y(n_4847)
);

NAND2xp5_ASAP7_75t_SL g4848 ( 
.A(n_4772),
.B(n_4778),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4775),
.Y(n_4849)
);

OAI21x1_ASAP7_75t_L g4850 ( 
.A1(n_4733),
.A2(n_4731),
.B(n_4693),
.Y(n_4850)
);

BUFx6f_ASAP7_75t_L g4851 ( 
.A(n_4711),
.Y(n_4851)
);

AND2x2_ASAP7_75t_L g4852 ( 
.A(n_4665),
.B(n_251),
.Y(n_4852)
);

OA21x2_ASAP7_75t_L g4853 ( 
.A1(n_4692),
.A2(n_4700),
.B(n_4776),
.Y(n_4853)
);

INVx2_ASAP7_75t_SL g4854 ( 
.A(n_4771),
.Y(n_4854)
);

INVx3_ASAP7_75t_L g4855 ( 
.A(n_4688),
.Y(n_4855)
);

BUFx6f_ASAP7_75t_L g4856 ( 
.A(n_4725),
.Y(n_4856)
);

BUFx4f_ASAP7_75t_L g4857 ( 
.A(n_4724),
.Y(n_4857)
);

AOI22xp33_ASAP7_75t_L g4858 ( 
.A1(n_4746),
.A2(n_637),
.B1(n_638),
.B2(n_636),
.Y(n_4858)
);

INVx2_ASAP7_75t_L g4859 ( 
.A(n_4671),
.Y(n_4859)
);

AND2x2_ASAP7_75t_L g4860 ( 
.A(n_4672),
.B(n_252),
.Y(n_4860)
);

CKINVDCx14_ASAP7_75t_R g4861 ( 
.A(n_4726),
.Y(n_4861)
);

INVx3_ASAP7_75t_L g4862 ( 
.A(n_4698),
.Y(n_4862)
);

AOI221xp5_ASAP7_75t_L g4863 ( 
.A1(n_4710),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.C(n_256),
.Y(n_4863)
);

INVx2_ASAP7_75t_L g4864 ( 
.A(n_4680),
.Y(n_4864)
);

NAND3xp33_ASAP7_75t_L g4865 ( 
.A(n_4739),
.B(n_641),
.C(n_639),
.Y(n_4865)
);

AOI22xp33_ASAP7_75t_L g4866 ( 
.A1(n_4741),
.A2(n_642),
.B1(n_643),
.B2(n_641),
.Y(n_4866)
);

AOI221xp5_ASAP7_75t_L g4867 ( 
.A1(n_4735),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.C(n_256),
.Y(n_4867)
);

INVx1_ASAP7_75t_L g4868 ( 
.A(n_4768),
.Y(n_4868)
);

OR2x2_ASAP7_75t_L g4869 ( 
.A(n_4770),
.B(n_256),
.Y(n_4869)
);

AOI21xp5_ASAP7_75t_L g4870 ( 
.A1(n_4747),
.A2(n_257),
.B(n_258),
.Y(n_4870)
);

AOI22xp33_ASAP7_75t_SL g4871 ( 
.A1(n_4730),
.A2(n_644),
.B1(n_645),
.B2(n_643),
.Y(n_4871)
);

OAI33xp33_ASAP7_75t_L g4872 ( 
.A1(n_4748),
.A2(n_259),
.A3(n_261),
.B1(n_257),
.B2(n_258),
.B3(n_260),
.Y(n_4872)
);

AOI22xp33_ASAP7_75t_L g4873 ( 
.A1(n_4674),
.A2(n_645),
.B1(n_646),
.B2(n_644),
.Y(n_4873)
);

AOI21xp33_ASAP7_75t_L g4874 ( 
.A1(n_4737),
.A2(n_647),
.B(n_646),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4742),
.Y(n_4875)
);

INVx2_ASAP7_75t_SL g4876 ( 
.A(n_4726),
.Y(n_4876)
);

OAI22xp5_ASAP7_75t_SL g4877 ( 
.A1(n_4773),
.A2(n_262),
.B1(n_259),
.B2(n_260),
.Y(n_4877)
);

CKINVDCx5p33_ASAP7_75t_R g4878 ( 
.A(n_4718),
.Y(n_4878)
);

AOI22xp33_ASAP7_75t_L g4879 ( 
.A1(n_4690),
.A2(n_649),
.B1(n_650),
.B2(n_648),
.Y(n_4879)
);

AOI22xp33_ASAP7_75t_L g4880 ( 
.A1(n_4691),
.A2(n_653),
.B1(n_654),
.B2(n_652),
.Y(n_4880)
);

OAI21xp5_ASAP7_75t_SL g4881 ( 
.A1(n_4713),
.A2(n_259),
.B(n_260),
.Y(n_4881)
);

NAND2xp5_ASAP7_75t_L g4882 ( 
.A(n_4670),
.B(n_654),
.Y(n_4882)
);

OA21x2_ASAP7_75t_L g4883 ( 
.A1(n_4720),
.A2(n_262),
.B(n_263),
.Y(n_4883)
);

OAI21x1_ASAP7_75t_L g4884 ( 
.A1(n_4723),
.A2(n_264),
.B(n_265),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4687),
.Y(n_4885)
);

AOI21xp33_ASAP7_75t_L g4886 ( 
.A1(n_4714),
.A2(n_656),
.B(n_655),
.Y(n_4886)
);

AOI22xp33_ASAP7_75t_L g4887 ( 
.A1(n_4763),
.A2(n_657),
.B1(n_658),
.B2(n_655),
.Y(n_4887)
);

NOR2xp33_ASAP7_75t_R g4888 ( 
.A(n_4767),
.B(n_657),
.Y(n_4888)
);

AOI22xp33_ASAP7_75t_L g4889 ( 
.A1(n_4763),
.A2(n_660),
.B1(n_662),
.B2(n_659),
.Y(n_4889)
);

OAI211xp5_ASAP7_75t_L g4890 ( 
.A1(n_4714),
.A2(n_269),
.B(n_267),
.C(n_268),
.Y(n_4890)
);

AOI22xp33_ASAP7_75t_L g4891 ( 
.A1(n_4763),
.A2(n_662),
.B1(n_664),
.B2(n_659),
.Y(n_4891)
);

HB1xp67_ASAP7_75t_L g4892 ( 
.A(n_4777),
.Y(n_4892)
);

OAI211xp5_ASAP7_75t_L g4893 ( 
.A1(n_4714),
.A2(n_269),
.B(n_267),
.C(n_268),
.Y(n_4893)
);

NOR2xp33_ASAP7_75t_L g4894 ( 
.A(n_4763),
.B(n_665),
.Y(n_4894)
);

AO31x2_ASAP7_75t_L g4895 ( 
.A1(n_4717),
.A2(n_272),
.A3(n_270),
.B(n_271),
.Y(n_4895)
);

OAI22xp5_ASAP7_75t_L g4896 ( 
.A1(n_4732),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_4896)
);

NAND2xp5_ASAP7_75t_L g4897 ( 
.A(n_4670),
.B(n_665),
.Y(n_4897)
);

AOI22xp33_ASAP7_75t_L g4898 ( 
.A1(n_4763),
.A2(n_667),
.B1(n_669),
.B2(n_666),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4670),
.B(n_666),
.Y(n_4899)
);

AOI22xp33_ASAP7_75t_L g4900 ( 
.A1(n_4763),
.A2(n_669),
.B1(n_670),
.B2(n_667),
.Y(n_4900)
);

AND2x4_ASAP7_75t_L g4901 ( 
.A(n_4675),
.B(n_670),
.Y(n_4901)
);

OR2x2_ASAP7_75t_L g4902 ( 
.A(n_4777),
.B(n_273),
.Y(n_4902)
);

AND2x2_ASAP7_75t_L g4903 ( 
.A(n_4675),
.B(n_274),
.Y(n_4903)
);

AOI22xp33_ASAP7_75t_L g4904 ( 
.A1(n_4763),
.A2(n_672),
.B1(n_673),
.B2(n_671),
.Y(n_4904)
);

AOI222xp33_ASAP7_75t_L g4905 ( 
.A1(n_4714),
.A2(n_277),
.B1(n_279),
.B2(n_275),
.C1(n_276),
.C2(n_278),
.Y(n_4905)
);

BUFx2_ASAP7_75t_L g4906 ( 
.A(n_4856),
.Y(n_4906)
);

HB1xp67_ASAP7_75t_L g4907 ( 
.A(n_4832),
.Y(n_4907)
);

INVx2_ASAP7_75t_L g4908 ( 
.A(n_4853),
.Y(n_4908)
);

INVx5_ASAP7_75t_L g4909 ( 
.A(n_4808),
.Y(n_4909)
);

INVxp67_ASAP7_75t_L g4910 ( 
.A(n_4786),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4811),
.Y(n_4911)
);

INVx3_ASAP7_75t_L g4912 ( 
.A(n_4856),
.Y(n_4912)
);

AND2x4_ASAP7_75t_L g4913 ( 
.A(n_4848),
.B(n_671),
.Y(n_4913)
);

NAND2xp5_ASAP7_75t_L g4914 ( 
.A(n_4843),
.B(n_672),
.Y(n_4914)
);

OR2x2_ASAP7_75t_L g4915 ( 
.A(n_4892),
.B(n_276),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4814),
.Y(n_4916)
);

BUFx2_ASAP7_75t_L g4917 ( 
.A(n_4861),
.Y(n_4917)
);

AND2x4_ASAP7_75t_L g4918 ( 
.A(n_4876),
.B(n_673),
.Y(n_4918)
);

OR2x2_ASAP7_75t_L g4919 ( 
.A(n_4791),
.B(n_277),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4827),
.Y(n_4920)
);

BUFx12f_ASAP7_75t_L g4921 ( 
.A(n_4808),
.Y(n_4921)
);

INVx1_ASAP7_75t_L g4922 ( 
.A(n_4835),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4841),
.Y(n_4923)
);

INVx2_ASAP7_75t_L g4924 ( 
.A(n_4826),
.Y(n_4924)
);

AND2x2_ASAP7_75t_L g4925 ( 
.A(n_4862),
.B(n_279),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4849),
.Y(n_4926)
);

NAND2xp5_ASAP7_75t_L g4927 ( 
.A(n_4885),
.B(n_674),
.Y(n_4927)
);

OAI22xp33_ASAP7_75t_L g4928 ( 
.A1(n_4784),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_4928)
);

AOI22xp33_ASAP7_75t_L g4929 ( 
.A1(n_4886),
.A2(n_675),
.B1(n_676),
.B2(n_674),
.Y(n_4929)
);

AND2x2_ASAP7_75t_L g4930 ( 
.A(n_4855),
.B(n_280),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4809),
.Y(n_4931)
);

AND2x2_ASAP7_75t_L g4932 ( 
.A(n_4854),
.B(n_283),
.Y(n_4932)
);

INVx2_ASAP7_75t_SL g4933 ( 
.A(n_4812),
.Y(n_4933)
);

INVx2_ASAP7_75t_L g4934 ( 
.A(n_4826),
.Y(n_4934)
);

NAND3xp33_ASAP7_75t_L g4935 ( 
.A(n_4905),
.B(n_283),
.C(n_284),
.Y(n_4935)
);

AND2x4_ASAP7_75t_L g4936 ( 
.A(n_4837),
.B(n_677),
.Y(n_4936)
);

INVx1_ASAP7_75t_SL g4937 ( 
.A(n_4888),
.Y(n_4937)
);

INVx2_ASAP7_75t_L g4938 ( 
.A(n_4826),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4816),
.Y(n_4939)
);

AND2x4_ASAP7_75t_SL g4940 ( 
.A(n_4810),
.B(n_678),
.Y(n_4940)
);

AND2x2_ASAP7_75t_L g4941 ( 
.A(n_4859),
.B(n_284),
.Y(n_4941)
);

OR2x2_ASAP7_75t_L g4942 ( 
.A(n_4868),
.B(n_285),
.Y(n_4942)
);

AND2x2_ASAP7_75t_L g4943 ( 
.A(n_4864),
.B(n_285),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_4830),
.B(n_680),
.Y(n_4944)
);

INVx2_ASAP7_75t_L g4945 ( 
.A(n_4826),
.Y(n_4945)
);

AOI22xp33_ASAP7_75t_SL g4946 ( 
.A1(n_4847),
.A2(n_682),
.B1(n_683),
.B2(n_681),
.Y(n_4946)
);

BUFx3_ASAP7_75t_L g4947 ( 
.A(n_4851),
.Y(n_4947)
);

AOI22xp33_ASAP7_75t_L g4948 ( 
.A1(n_4787),
.A2(n_684),
.B1(n_685),
.B2(n_683),
.Y(n_4948)
);

AND2x2_ASAP7_75t_L g4949 ( 
.A(n_4783),
.B(n_285),
.Y(n_4949)
);

OAI21xp5_ASAP7_75t_SL g4950 ( 
.A1(n_4890),
.A2(n_286),
.B(n_287),
.Y(n_4950)
);

AND2x4_ASAP7_75t_L g4951 ( 
.A(n_4845),
.B(n_4793),
.Y(n_4951)
);

HB1xp67_ASAP7_75t_L g4952 ( 
.A(n_4850),
.Y(n_4952)
);

NOR2xp33_ASAP7_75t_SL g4953 ( 
.A(n_4799),
.B(n_684),
.Y(n_4953)
);

BUFx6f_ASAP7_75t_L g4954 ( 
.A(n_4851),
.Y(n_4954)
);

AND2x4_ASAP7_75t_L g4955 ( 
.A(n_4797),
.B(n_685),
.Y(n_4955)
);

INVxp67_ASAP7_75t_L g4956 ( 
.A(n_4894),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4875),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4869),
.Y(n_4958)
);

CKINVDCx5p33_ASAP7_75t_R g4959 ( 
.A(n_4878),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_4817),
.Y(n_4960)
);

AND2x2_ASAP7_75t_L g4961 ( 
.A(n_4903),
.B(n_288),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4844),
.Y(n_4962)
);

NAND2xp5_ASAP7_75t_L g4963 ( 
.A(n_4802),
.B(n_686),
.Y(n_4963)
);

OR2x2_ASAP7_75t_L g4964 ( 
.A(n_4779),
.B(n_289),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4834),
.Y(n_4965)
);

BUFx3_ASAP7_75t_L g4966 ( 
.A(n_4857),
.Y(n_4966)
);

INVx1_ASAP7_75t_L g4967 ( 
.A(n_4836),
.Y(n_4967)
);

OR2x2_ASAP7_75t_L g4968 ( 
.A(n_4902),
.B(n_289),
.Y(n_4968)
);

NOR2xp33_ASAP7_75t_L g4969 ( 
.A(n_4780),
.B(n_687),
.Y(n_4969)
);

INVx2_ASAP7_75t_L g4970 ( 
.A(n_4852),
.Y(n_4970)
);

BUFx2_ASAP7_75t_L g4971 ( 
.A(n_4901),
.Y(n_4971)
);

INVx2_ASAP7_75t_L g4972 ( 
.A(n_4860),
.Y(n_4972)
);

HB1xp67_ASAP7_75t_L g4973 ( 
.A(n_4883),
.Y(n_4973)
);

NAND2xp5_ASAP7_75t_L g4974 ( 
.A(n_4882),
.B(n_687),
.Y(n_4974)
);

BUFx3_ASAP7_75t_L g4975 ( 
.A(n_4800),
.Y(n_4975)
);

OR2x2_ASAP7_75t_L g4976 ( 
.A(n_4897),
.B(n_290),
.Y(n_4976)
);

INVx2_ASAP7_75t_L g4977 ( 
.A(n_4792),
.Y(n_4977)
);

OR2x2_ASAP7_75t_L g4978 ( 
.A(n_4899),
.B(n_290),
.Y(n_4978)
);

INVxp67_ASAP7_75t_L g4979 ( 
.A(n_4806),
.Y(n_4979)
);

HB1xp67_ASAP7_75t_L g4980 ( 
.A(n_4895),
.Y(n_4980)
);

AND2x2_ASAP7_75t_L g4981 ( 
.A(n_4818),
.B(n_290),
.Y(n_4981)
);

INVx2_ASAP7_75t_L g4982 ( 
.A(n_4895),
.Y(n_4982)
);

NAND2xp5_ASAP7_75t_L g4983 ( 
.A(n_4803),
.B(n_688),
.Y(n_4983)
);

OAI22xp5_ASAP7_75t_L g4984 ( 
.A1(n_4873),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_4984)
);

AND2x2_ASAP7_75t_L g4985 ( 
.A(n_4828),
.B(n_291),
.Y(n_4985)
);

INVx1_ASAP7_75t_L g4986 ( 
.A(n_4782),
.Y(n_4986)
);

INVx1_ASAP7_75t_SL g4987 ( 
.A(n_4801),
.Y(n_4987)
);

OR2x2_ASAP7_75t_L g4988 ( 
.A(n_4881),
.B(n_291),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_4838),
.Y(n_4989)
);

AND2x2_ASAP7_75t_L g4990 ( 
.A(n_4781),
.B(n_292),
.Y(n_4990)
);

INVx1_ASAP7_75t_L g4991 ( 
.A(n_4842),
.Y(n_4991)
);

AND2x2_ASAP7_75t_L g4992 ( 
.A(n_4884),
.B(n_293),
.Y(n_4992)
);

AOI222xp33_ASAP7_75t_L g4993 ( 
.A1(n_4877),
.A2(n_296),
.B1(n_298),
.B2(n_294),
.C1(n_295),
.C2(n_297),
.Y(n_4993)
);

AND2x2_ASAP7_75t_L g4994 ( 
.A(n_4796),
.B(n_4824),
.Y(n_4994)
);

INVx2_ASAP7_75t_L g4995 ( 
.A(n_4823),
.Y(n_4995)
);

INVx4_ASAP7_75t_L g4996 ( 
.A(n_4831),
.Y(n_4996)
);

INVx1_ASAP7_75t_L g4997 ( 
.A(n_4870),
.Y(n_4997)
);

NAND2xp33_ASAP7_75t_R g4998 ( 
.A(n_4840),
.B(n_294),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4865),
.Y(n_4999)
);

AND2x4_ASAP7_75t_L g5000 ( 
.A(n_4813),
.B(n_689),
.Y(n_5000)
);

AND2x2_ASAP7_75t_L g5001 ( 
.A(n_4866),
.B(n_297),
.Y(n_5001)
);

AND2x2_ASAP7_75t_L g5002 ( 
.A(n_4846),
.B(n_298),
.Y(n_5002)
);

AND2x2_ASAP7_75t_L g5003 ( 
.A(n_4790),
.B(n_298),
.Y(n_5003)
);

AND2x2_ASAP7_75t_L g5004 ( 
.A(n_4879),
.B(n_4805),
.Y(n_5004)
);

BUFx3_ASAP7_75t_L g5005 ( 
.A(n_4829),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_4825),
.Y(n_5006)
);

AND2x2_ASAP7_75t_L g5007 ( 
.A(n_4822),
.B(n_299),
.Y(n_5007)
);

NOR2xp67_ASAP7_75t_L g5008 ( 
.A(n_4893),
.B(n_299),
.Y(n_5008)
);

AND2x2_ASAP7_75t_L g5009 ( 
.A(n_4880),
.B(n_299),
.Y(n_5009)
);

OAI22xp5_ASAP7_75t_L g5010 ( 
.A1(n_4785),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4807),
.Y(n_5011)
);

AND2x2_ASAP7_75t_L g5012 ( 
.A(n_4820),
.B(n_300),
.Y(n_5012)
);

AND2x2_ASAP7_75t_L g5013 ( 
.A(n_4871),
.B(n_4874),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4798),
.Y(n_5014)
);

AND2x2_ASAP7_75t_L g5015 ( 
.A(n_4795),
.B(n_300),
.Y(n_5015)
);

HB1xp67_ASAP7_75t_L g5016 ( 
.A(n_4839),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4804),
.Y(n_5017)
);

INVx1_ASAP7_75t_L g5018 ( 
.A(n_4815),
.Y(n_5018)
);

NOR2x1p5_ASAP7_75t_L g5019 ( 
.A(n_4872),
.B(n_301),
.Y(n_5019)
);

INVx2_ASAP7_75t_L g5020 ( 
.A(n_4896),
.Y(n_5020)
);

NOR2xp67_ASAP7_75t_L g5021 ( 
.A(n_4788),
.B(n_4858),
.Y(n_5021)
);

AND2x4_ASAP7_75t_L g5022 ( 
.A(n_4819),
.B(n_690),
.Y(n_5022)
);

NAND2xp5_ASAP7_75t_L g5023 ( 
.A(n_4863),
.B(n_691),
.Y(n_5023)
);

NOR2xp33_ASAP7_75t_L g5024 ( 
.A(n_4789),
.B(n_691),
.Y(n_5024)
);

INVx1_ASAP7_75t_L g5025 ( 
.A(n_4867),
.Y(n_5025)
);

HB1xp67_ASAP7_75t_L g5026 ( 
.A(n_4794),
.Y(n_5026)
);

AND2x2_ASAP7_75t_L g5027 ( 
.A(n_4821),
.B(n_303),
.Y(n_5027)
);

INVx5_ASAP7_75t_L g5028 ( 
.A(n_4833),
.Y(n_5028)
);

AND2x2_ASAP7_75t_L g5029 ( 
.A(n_4887),
.B(n_303),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_4889),
.Y(n_5030)
);

INVx2_ASAP7_75t_L g5031 ( 
.A(n_4891),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_L g5032 ( 
.A(n_4898),
.B(n_4900),
.Y(n_5032)
);

AND2x2_ASAP7_75t_L g5033 ( 
.A(n_4904),
.B(n_303),
.Y(n_5033)
);

INVxp67_ASAP7_75t_SL g5034 ( 
.A(n_4832),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_4811),
.Y(n_5035)
);

INVx2_ASAP7_75t_L g5036 ( 
.A(n_4853),
.Y(n_5036)
);

INVxp67_ASAP7_75t_SL g5037 ( 
.A(n_4832),
.Y(n_5037)
);

INVx1_ASAP7_75t_SL g5038 ( 
.A(n_4888),
.Y(n_5038)
);

CKINVDCx6p67_ASAP7_75t_R g5039 ( 
.A(n_4812),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_4843),
.B(n_692),
.Y(n_5040)
);

NAND2xp5_ASAP7_75t_L g5041 ( 
.A(n_4843),
.B(n_692),
.Y(n_5041)
);

AND2x4_ASAP7_75t_L g5042 ( 
.A(n_4848),
.B(n_694),
.Y(n_5042)
);

INVx1_ASAP7_75t_L g5043 ( 
.A(n_4811),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_4811),
.Y(n_5044)
);

AND2x2_ASAP7_75t_L g5045 ( 
.A(n_4892),
.B(n_305),
.Y(n_5045)
);

AND2x4_ASAP7_75t_L g5046 ( 
.A(n_4848),
.B(n_695),
.Y(n_5046)
);

NOR2x1_ASAP7_75t_L g5047 ( 
.A(n_4837),
.B(n_306),
.Y(n_5047)
);

INVx2_ASAP7_75t_SL g5048 ( 
.A(n_4856),
.Y(n_5048)
);

INVx1_ASAP7_75t_L g5049 ( 
.A(n_4811),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_4843),
.B(n_695),
.Y(n_5050)
);

HB1xp67_ASAP7_75t_L g5051 ( 
.A(n_4832),
.Y(n_5051)
);

NAND2xp5_ASAP7_75t_L g5052 ( 
.A(n_4999),
.B(n_696),
.Y(n_5052)
);

AND2x2_ASAP7_75t_L g5053 ( 
.A(n_4906),
.B(n_306),
.Y(n_5053)
);

HB1xp67_ASAP7_75t_L g5054 ( 
.A(n_4973),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_4911),
.Y(n_5055)
);

AND2x2_ASAP7_75t_L g5056 ( 
.A(n_4917),
.B(n_307),
.Y(n_5056)
);

AND2x2_ASAP7_75t_L g5057 ( 
.A(n_4912),
.B(n_307),
.Y(n_5057)
);

AND2x2_ASAP7_75t_L g5058 ( 
.A(n_4910),
.B(n_307),
.Y(n_5058)
);

NOR2xp33_ASAP7_75t_L g5059 ( 
.A(n_4909),
.B(n_696),
.Y(n_5059)
);

AND2x2_ASAP7_75t_L g5060 ( 
.A(n_5048),
.B(n_308),
.Y(n_5060)
);

NOR2x1_ASAP7_75t_SL g5061 ( 
.A(n_4977),
.B(n_308),
.Y(n_5061)
);

NAND2xp5_ASAP7_75t_L g5062 ( 
.A(n_4997),
.B(n_697),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_L g5063 ( 
.A(n_4979),
.B(n_698),
.Y(n_5063)
);

NAND2x1_ASAP7_75t_SL g5064 ( 
.A(n_5047),
.B(n_4907),
.Y(n_5064)
);

NAND2xp5_ASAP7_75t_L g5065 ( 
.A(n_4986),
.B(n_700),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_4916),
.Y(n_5066)
);

OR2x2_ASAP7_75t_L g5067 ( 
.A(n_4960),
.B(n_308),
.Y(n_5067)
);

AND2x4_ASAP7_75t_L g5068 ( 
.A(n_4933),
.B(n_4958),
.Y(n_5068)
);

NAND2xp5_ASAP7_75t_L g5069 ( 
.A(n_4967),
.B(n_701),
.Y(n_5069)
);

INVx2_ASAP7_75t_L g5070 ( 
.A(n_4908),
.Y(n_5070)
);

OR2x2_ASAP7_75t_L g5071 ( 
.A(n_4962),
.B(n_309),
.Y(n_5071)
);

AND2x4_ASAP7_75t_SL g5072 ( 
.A(n_5039),
.B(n_309),
.Y(n_5072)
);

NAND3xp33_ASAP7_75t_L g5073 ( 
.A(n_4998),
.B(n_309),
.C(n_310),
.Y(n_5073)
);

OR2x2_ASAP7_75t_L g5074 ( 
.A(n_4965),
.B(n_5051),
.Y(n_5074)
);

AND2x4_ASAP7_75t_L g5075 ( 
.A(n_4971),
.B(n_310),
.Y(n_5075)
);

NAND2xp5_ASAP7_75t_L g5076 ( 
.A(n_4991),
.B(n_702),
.Y(n_5076)
);

INVx1_ASAP7_75t_L g5077 ( 
.A(n_4920),
.Y(n_5077)
);

AOI221xp5_ASAP7_75t_L g5078 ( 
.A1(n_5026),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.C(n_314),
.Y(n_5078)
);

INVx5_ASAP7_75t_L g5079 ( 
.A(n_4921),
.Y(n_5079)
);

HB1xp67_ASAP7_75t_L g5080 ( 
.A(n_4980),
.Y(n_5080)
);

AND2x2_ASAP7_75t_L g5081 ( 
.A(n_4970),
.B(n_312),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_4922),
.Y(n_5082)
);

INVx2_ASAP7_75t_L g5083 ( 
.A(n_5036),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4923),
.Y(n_5084)
);

AND2x4_ASAP7_75t_L g5085 ( 
.A(n_4972),
.B(n_312),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_4926),
.Y(n_5086)
);

NAND3xp33_ASAP7_75t_L g5087 ( 
.A(n_4953),
.B(n_313),
.C(n_314),
.Y(n_5087)
);

INVx2_ASAP7_75t_L g5088 ( 
.A(n_4924),
.Y(n_5088)
);

NAND2xp5_ASAP7_75t_L g5089 ( 
.A(n_4914),
.B(n_704),
.Y(n_5089)
);

AND2x2_ASAP7_75t_L g5090 ( 
.A(n_5034),
.B(n_315),
.Y(n_5090)
);

AND2x2_ASAP7_75t_L g5091 ( 
.A(n_5037),
.B(n_316),
.Y(n_5091)
);

NOR2xp33_ASAP7_75t_L g5092 ( 
.A(n_4956),
.B(n_704),
.Y(n_5092)
);

AND2x4_ASAP7_75t_L g5093 ( 
.A(n_4966),
.B(n_317),
.Y(n_5093)
);

NAND2xp5_ASAP7_75t_L g5094 ( 
.A(n_5040),
.B(n_705),
.Y(n_5094)
);

NAND2xp5_ASAP7_75t_L g5095 ( 
.A(n_5041),
.B(n_706),
.Y(n_5095)
);

OR2x2_ASAP7_75t_L g5096 ( 
.A(n_4989),
.B(n_318),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_5035),
.Y(n_5097)
);

INVx2_ASAP7_75t_L g5098 ( 
.A(n_4934),
.Y(n_5098)
);

HB1xp67_ASAP7_75t_L g5099 ( 
.A(n_4982),
.Y(n_5099)
);

AOI221xp5_ASAP7_75t_L g5100 ( 
.A1(n_5005),
.A2(n_320),
.B1(n_318),
.B2(n_319),
.C(n_321),
.Y(n_5100)
);

INVx1_ASAP7_75t_L g5101 ( 
.A(n_5043),
.Y(n_5101)
);

INVx2_ASAP7_75t_L g5102 ( 
.A(n_4938),
.Y(n_5102)
);

INVxp67_ASAP7_75t_SL g5103 ( 
.A(n_4952),
.Y(n_5103)
);

AND2x2_ASAP7_75t_L g5104 ( 
.A(n_4931),
.B(n_319),
.Y(n_5104)
);

INVx2_ASAP7_75t_L g5105 ( 
.A(n_4945),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_5044),
.Y(n_5106)
);

OR2x2_ASAP7_75t_L g5107 ( 
.A(n_4939),
.B(n_319),
.Y(n_5107)
);

NAND2xp5_ASAP7_75t_L g5108 ( 
.A(n_5050),
.B(n_707),
.Y(n_5108)
);

INVx1_ASAP7_75t_L g5109 ( 
.A(n_5049),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_4957),
.Y(n_5110)
);

AND2x4_ASAP7_75t_L g5111 ( 
.A(n_4975),
.B(n_320),
.Y(n_5111)
);

NAND2xp5_ASAP7_75t_L g5112 ( 
.A(n_4994),
.B(n_708),
.Y(n_5112)
);

INVx1_ASAP7_75t_L g5113 ( 
.A(n_4942),
.Y(n_5113)
);

INVx2_ASAP7_75t_L g5114 ( 
.A(n_4949),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_4941),
.Y(n_5115)
);

HB1xp67_ASAP7_75t_SL g5116 ( 
.A(n_4996),
.Y(n_5116)
);

BUFx3_ASAP7_75t_L g5117 ( 
.A(n_4947),
.Y(n_5117)
);

OR2x2_ASAP7_75t_L g5118 ( 
.A(n_4919),
.B(n_321),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_4943),
.Y(n_5119)
);

INVx2_ASAP7_75t_SL g5120 ( 
.A(n_4954),
.Y(n_5120)
);

HB1xp67_ASAP7_75t_L g5121 ( 
.A(n_4915),
.Y(n_5121)
);

OR2x2_ASAP7_75t_L g5122 ( 
.A(n_4927),
.B(n_322),
.Y(n_5122)
);

INVx1_ASAP7_75t_L g5123 ( 
.A(n_4944),
.Y(n_5123)
);

INVx2_ASAP7_75t_L g5124 ( 
.A(n_4930),
.Y(n_5124)
);

NAND4xp25_ASAP7_75t_L g5125 ( 
.A(n_4935),
.B(n_325),
.C(n_323),
.D(n_324),
.Y(n_5125)
);

OAI22xp5_ASAP7_75t_L g5126 ( 
.A1(n_5028),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_5045),
.Y(n_5127)
);

OAI221xp5_ASAP7_75t_SL g5128 ( 
.A1(n_4950),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.C(n_328),
.Y(n_5128)
);

NAND2xp5_ASAP7_75t_L g5129 ( 
.A(n_4995),
.B(n_708),
.Y(n_5129)
);

NAND2xp5_ASAP7_75t_SL g5130 ( 
.A(n_4959),
.B(n_327),
.Y(n_5130)
);

AND2x4_ASAP7_75t_L g5131 ( 
.A(n_4925),
.B(n_328),
.Y(n_5131)
);

AND2x2_ASAP7_75t_L g5132 ( 
.A(n_5014),
.B(n_328),
.Y(n_5132)
);

AND2x2_ASAP7_75t_L g5133 ( 
.A(n_5016),
.B(n_4913),
.Y(n_5133)
);

AND2x2_ASAP7_75t_L g5134 ( 
.A(n_5042),
.B(n_5046),
.Y(n_5134)
);

AND2x2_ASAP7_75t_L g5135 ( 
.A(n_5020),
.B(n_329),
.Y(n_5135)
);

INVx2_ASAP7_75t_L g5136 ( 
.A(n_4918),
.Y(n_5136)
);

INVx1_ASAP7_75t_L g5137 ( 
.A(n_4990),
.Y(n_5137)
);

NAND4xp25_ASAP7_75t_L g5138 ( 
.A(n_5008),
.B(n_332),
.C(n_330),
.D(n_331),
.Y(n_5138)
);

INVx1_ASAP7_75t_L g5139 ( 
.A(n_4992),
.Y(n_5139)
);

AND2x2_ASAP7_75t_L g5140 ( 
.A(n_4955),
.B(n_4932),
.Y(n_5140)
);

OR2x2_ASAP7_75t_L g5141 ( 
.A(n_4976),
.B(n_330),
.Y(n_5141)
);

BUFx2_ASAP7_75t_L g5142 ( 
.A(n_4936),
.Y(n_5142)
);

INVx2_ASAP7_75t_L g5143 ( 
.A(n_4964),
.Y(n_5143)
);

NAND2xp5_ASAP7_75t_L g5144 ( 
.A(n_5018),
.B(n_709),
.Y(n_5144)
);

BUFx6f_ASAP7_75t_L g5145 ( 
.A(n_4968),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_4978),
.Y(n_5146)
);

NOR2xp33_ASAP7_75t_L g5147 ( 
.A(n_4937),
.B(n_709),
.Y(n_5147)
);

INVx2_ASAP7_75t_L g5148 ( 
.A(n_4985),
.Y(n_5148)
);

NAND2xp5_ASAP7_75t_L g5149 ( 
.A(n_4969),
.B(n_710),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_5006),
.Y(n_5150)
);

INVx2_ASAP7_75t_L g5151 ( 
.A(n_4981),
.Y(n_5151)
);

HB1xp67_ASAP7_75t_L g5152 ( 
.A(n_5011),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_4983),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_5030),
.Y(n_5154)
);

AND2x2_ASAP7_75t_L g5155 ( 
.A(n_4961),
.B(n_332),
.Y(n_5155)
);

NAND3xp33_ASAP7_75t_L g5156 ( 
.A(n_5028),
.B(n_332),
.C(n_333),
.Y(n_5156)
);

INVxp67_ASAP7_75t_L g5157 ( 
.A(n_4988),
.Y(n_5157)
);

AND2x2_ASAP7_75t_L g5158 ( 
.A(n_5038),
.B(n_333),
.Y(n_5158)
);

AND2x2_ASAP7_75t_L g5159 ( 
.A(n_5031),
.B(n_333),
.Y(n_5159)
);

NAND2xp5_ASAP7_75t_L g5160 ( 
.A(n_5000),
.B(n_711),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_5013),
.B(n_711),
.Y(n_5161)
);

INVx1_ASAP7_75t_L g5162 ( 
.A(n_4963),
.Y(n_5162)
);

AND2x2_ASAP7_75t_L g5163 ( 
.A(n_4987),
.B(n_334),
.Y(n_5163)
);

NAND2xp5_ASAP7_75t_L g5164 ( 
.A(n_4974),
.B(n_713),
.Y(n_5164)
);

INVx2_ASAP7_75t_L g5165 ( 
.A(n_5017),
.Y(n_5165)
);

NAND3xp33_ASAP7_75t_L g5166 ( 
.A(n_5025),
.B(n_5024),
.C(n_4946),
.Y(n_5166)
);

INVx1_ASAP7_75t_L g5167 ( 
.A(n_5004),
.Y(n_5167)
);

INVx2_ASAP7_75t_L g5168 ( 
.A(n_4940),
.Y(n_5168)
);

INVx5_ASAP7_75t_L g5169 ( 
.A(n_5003),
.Y(n_5169)
);

AND2x4_ASAP7_75t_L g5170 ( 
.A(n_5021),
.B(n_334),
.Y(n_5170)
);

NAND2xp5_ASAP7_75t_L g5171 ( 
.A(n_5019),
.B(n_714),
.Y(n_5171)
);

AND2x2_ASAP7_75t_L g5172 ( 
.A(n_5015),
.B(n_335),
.Y(n_5172)
);

AND2x4_ASAP7_75t_L g5173 ( 
.A(n_5032),
.B(n_335),
.Y(n_5173)
);

AND2x4_ASAP7_75t_L g5174 ( 
.A(n_5029),
.B(n_336),
.Y(n_5174)
);

AND2x2_ASAP7_75t_SL g5175 ( 
.A(n_4948),
.B(n_336),
.Y(n_5175)
);

AND2x2_ASAP7_75t_L g5176 ( 
.A(n_5009),
.B(n_337),
.Y(n_5176)
);

NAND2xp5_ASAP7_75t_L g5177 ( 
.A(n_4928),
.B(n_714),
.Y(n_5177)
);

OR2x2_ASAP7_75t_L g5178 ( 
.A(n_5023),
.B(n_337),
.Y(n_5178)
);

AND2x2_ASAP7_75t_L g5179 ( 
.A(n_5002),
.B(n_337),
.Y(n_5179)
);

AND2x2_ASAP7_75t_L g5180 ( 
.A(n_5027),
.B(n_338),
.Y(n_5180)
);

INVx1_ASAP7_75t_L g5181 ( 
.A(n_5001),
.Y(n_5181)
);

HB1xp67_ASAP7_75t_L g5182 ( 
.A(n_5033),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_5007),
.Y(n_5183)
);

AND2x2_ASAP7_75t_L g5184 ( 
.A(n_5022),
.B(n_338),
.Y(n_5184)
);

NAND2xp5_ASAP7_75t_L g5185 ( 
.A(n_4929),
.B(n_715),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_5012),
.Y(n_5186)
);

OR2x2_ASAP7_75t_L g5187 ( 
.A(n_4984),
.B(n_338),
.Y(n_5187)
);

NAND2xp5_ASAP7_75t_L g5188 ( 
.A(n_5010),
.B(n_715),
.Y(n_5188)
);

NAND2xp5_ASAP7_75t_L g5189 ( 
.A(n_4999),
.B(n_716),
.Y(n_5189)
);

AND2x4_ASAP7_75t_L g5190 ( 
.A(n_4917),
.B(n_339),
.Y(n_5190)
);

HB1xp67_ASAP7_75t_L g5191 ( 
.A(n_4973),
.Y(n_5191)
);

AND2x2_ASAP7_75t_L g5192 ( 
.A(n_4906),
.B(n_339),
.Y(n_5192)
);

INVx1_ASAP7_75t_L g5193 ( 
.A(n_4911),
.Y(n_5193)
);

AND2x2_ASAP7_75t_L g5194 ( 
.A(n_4906),
.B(n_340),
.Y(n_5194)
);

AND2x4_ASAP7_75t_SL g5195 ( 
.A(n_5039),
.B(n_340),
.Y(n_5195)
);

BUFx2_ASAP7_75t_SL g5196 ( 
.A(n_4909),
.Y(n_5196)
);

NOR2xp33_ASAP7_75t_L g5197 ( 
.A(n_4909),
.B(n_716),
.Y(n_5197)
);

HB1xp67_ASAP7_75t_L g5198 ( 
.A(n_4973),
.Y(n_5198)
);

AND2x2_ASAP7_75t_L g5199 ( 
.A(n_4906),
.B(n_341),
.Y(n_5199)
);

AND2x2_ASAP7_75t_L g5200 ( 
.A(n_4906),
.B(n_341),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_4911),
.Y(n_5201)
);

AND2x2_ASAP7_75t_L g5202 ( 
.A(n_4906),
.B(n_342),
.Y(n_5202)
);

INVxp33_ASAP7_75t_L g5203 ( 
.A(n_4917),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_4911),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_4911),
.Y(n_5205)
);

OAI211xp5_ASAP7_75t_L g5206 ( 
.A1(n_4993),
.A2(n_344),
.B(n_342),
.C(n_343),
.Y(n_5206)
);

INVx2_ASAP7_75t_L g5207 ( 
.A(n_4951),
.Y(n_5207)
);

NAND2x1_ASAP7_75t_L g5208 ( 
.A(n_4906),
.B(n_343),
.Y(n_5208)
);

AND2x2_ASAP7_75t_L g5209 ( 
.A(n_4906),
.B(n_344),
.Y(n_5209)
);

AND2x2_ASAP7_75t_L g5210 ( 
.A(n_4906),
.B(n_345),
.Y(n_5210)
);

AND2x2_ASAP7_75t_L g5211 ( 
.A(n_4906),
.B(n_345),
.Y(n_5211)
);

OR2x2_ASAP7_75t_L g5212 ( 
.A(n_4960),
.B(n_346),
.Y(n_5212)
);

AND2x2_ASAP7_75t_L g5213 ( 
.A(n_4906),
.B(n_346),
.Y(n_5213)
);

INVx1_ASAP7_75t_L g5214 ( 
.A(n_4911),
.Y(n_5214)
);

NOR2xp33_ASAP7_75t_L g5215 ( 
.A(n_4909),
.B(n_717),
.Y(n_5215)
);

AND2x4_ASAP7_75t_L g5216 ( 
.A(n_4917),
.B(n_346),
.Y(n_5216)
);

BUFx3_ASAP7_75t_L g5217 ( 
.A(n_4921),
.Y(n_5217)
);

BUFx2_ASAP7_75t_L g5218 ( 
.A(n_4917),
.Y(n_5218)
);

NAND2xp5_ASAP7_75t_L g5219 ( 
.A(n_4999),
.B(n_717),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_4911),
.Y(n_5220)
);

OR2x2_ASAP7_75t_L g5221 ( 
.A(n_4960),
.B(n_347),
.Y(n_5221)
);

NOR2xp67_ASAP7_75t_L g5222 ( 
.A(n_4909),
.B(n_347),
.Y(n_5222)
);

INVx1_ASAP7_75t_L g5223 ( 
.A(n_4911),
.Y(n_5223)
);

INVx1_ASAP7_75t_L g5224 ( 
.A(n_4911),
.Y(n_5224)
);

HB1xp67_ASAP7_75t_L g5225 ( 
.A(n_4973),
.Y(n_5225)
);

NAND2xp5_ASAP7_75t_SL g5226 ( 
.A(n_4999),
.B(n_348),
.Y(n_5226)
);

AND2x2_ASAP7_75t_L g5227 ( 
.A(n_4906),
.B(n_348),
.Y(n_5227)
);

NAND2x1p5_ASAP7_75t_L g5228 ( 
.A(n_4906),
.B(n_349),
.Y(n_5228)
);

INVx2_ASAP7_75t_L g5229 ( 
.A(n_4951),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_4911),
.Y(n_5230)
);

AND2x2_ASAP7_75t_L g5231 ( 
.A(n_4906),
.B(n_350),
.Y(n_5231)
);

INVx1_ASAP7_75t_L g5232 ( 
.A(n_4911),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_4911),
.Y(n_5233)
);

HB1xp67_ASAP7_75t_L g5234 ( 
.A(n_4973),
.Y(n_5234)
);

AOI221xp5_ASAP7_75t_L g5235 ( 
.A1(n_5026),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.C(n_353),
.Y(n_5235)
);

INVx3_ASAP7_75t_L g5236 ( 
.A(n_5217),
.Y(n_5236)
);

INVx1_ASAP7_75t_L g5237 ( 
.A(n_5054),
.Y(n_5237)
);

OAI321xp33_ASAP7_75t_L g5238 ( 
.A1(n_5073),
.A2(n_375),
.A3(n_359),
.B1(n_383),
.B2(n_367),
.C(n_351),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_5191),
.Y(n_5239)
);

BUFx2_ASAP7_75t_L g5240 ( 
.A(n_5064),
.Y(n_5240)
);

INVx1_ASAP7_75t_SL g5241 ( 
.A(n_5196),
.Y(n_5241)
);

AND2x2_ASAP7_75t_L g5242 ( 
.A(n_5218),
.B(n_354),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_5198),
.Y(n_5243)
);

AOI31xp33_ASAP7_75t_SL g5244 ( 
.A1(n_5100),
.A2(n_359),
.A3(n_357),
.B(n_358),
.Y(n_5244)
);

NAND2xp5_ASAP7_75t_L g5245 ( 
.A(n_5165),
.B(n_357),
.Y(n_5245)
);

AOI22xp33_ASAP7_75t_L g5246 ( 
.A1(n_5167),
.A2(n_360),
.B1(n_357),
.B2(n_359),
.Y(n_5246)
);

NAND3xp33_ASAP7_75t_L g5247 ( 
.A(n_5156),
.B(n_360),
.C(n_361),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_5225),
.Y(n_5248)
);

INVx4_ASAP7_75t_L g5249 ( 
.A(n_5079),
.Y(n_5249)
);

OAI31xp33_ASAP7_75t_L g5250 ( 
.A1(n_5206),
.A2(n_363),
.A3(n_364),
.B(n_362),
.Y(n_5250)
);

AO31x2_ASAP7_75t_L g5251 ( 
.A1(n_5126),
.A2(n_364),
.A3(n_361),
.B(n_363),
.Y(n_5251)
);

NOR2xp33_ASAP7_75t_L g5252 ( 
.A(n_5079),
.B(n_5203),
.Y(n_5252)
);

OR2x2_ASAP7_75t_L g5253 ( 
.A(n_5154),
.B(n_365),
.Y(n_5253)
);

AND2x2_ASAP7_75t_L g5254 ( 
.A(n_5152),
.B(n_366),
.Y(n_5254)
);

INVx1_ASAP7_75t_L g5255 ( 
.A(n_5234),
.Y(n_5255)
);

INVxp33_ASAP7_75t_L g5256 ( 
.A(n_5116),
.Y(n_5256)
);

OR2x2_ASAP7_75t_L g5257 ( 
.A(n_5074),
.B(n_367),
.Y(n_5257)
);

INVx2_ASAP7_75t_L g5258 ( 
.A(n_5145),
.Y(n_5258)
);

INVx2_ASAP7_75t_L g5259 ( 
.A(n_5145),
.Y(n_5259)
);

INVx1_ASAP7_75t_L g5260 ( 
.A(n_5055),
.Y(n_5260)
);

NAND2xp5_ASAP7_75t_L g5261 ( 
.A(n_5150),
.B(n_368),
.Y(n_5261)
);

NAND2x1_ASAP7_75t_SL g5262 ( 
.A(n_5222),
.B(n_368),
.Y(n_5262)
);

INVx2_ASAP7_75t_SL g5263 ( 
.A(n_5117),
.Y(n_5263)
);

AO21x2_ASAP7_75t_L g5264 ( 
.A1(n_5080),
.A2(n_369),
.B(n_370),
.Y(n_5264)
);

INVx2_ASAP7_75t_L g5265 ( 
.A(n_5068),
.Y(n_5265)
);

INVx1_ASAP7_75t_L g5266 ( 
.A(n_5066),
.Y(n_5266)
);

INVx2_ASAP7_75t_L g5267 ( 
.A(n_5142),
.Y(n_5267)
);

AOI221xp5_ASAP7_75t_L g5268 ( 
.A1(n_5166),
.A2(n_5170),
.B1(n_5235),
.B2(n_5078),
.C(n_5128),
.Y(n_5268)
);

NAND2xp5_ASAP7_75t_L g5269 ( 
.A(n_5146),
.B(n_371),
.Y(n_5269)
);

NAND2xp5_ASAP7_75t_L g5270 ( 
.A(n_5169),
.B(n_372),
.Y(n_5270)
);

INVxp67_ASAP7_75t_SL g5271 ( 
.A(n_5061),
.Y(n_5271)
);

HB1xp67_ASAP7_75t_L g5272 ( 
.A(n_5121),
.Y(n_5272)
);

AND2x2_ASAP7_75t_L g5273 ( 
.A(n_5207),
.B(n_5229),
.Y(n_5273)
);

NAND2xp5_ASAP7_75t_L g5274 ( 
.A(n_5133),
.B(n_373),
.Y(n_5274)
);

AOI22xp33_ASAP7_75t_L g5275 ( 
.A1(n_5175),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_5275)
);

CKINVDCx16_ASAP7_75t_R g5276 ( 
.A(n_5190),
.Y(n_5276)
);

AOI21xp5_ASAP7_75t_L g5277 ( 
.A1(n_5226),
.A2(n_376),
.B(n_377),
.Y(n_5277)
);

AND2x4_ASAP7_75t_L g5278 ( 
.A(n_5120),
.B(n_377),
.Y(n_5278)
);

OR2x2_ASAP7_75t_L g5279 ( 
.A(n_5143),
.B(n_377),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_5077),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_5082),
.Y(n_5281)
);

AND2x2_ASAP7_75t_L g5282 ( 
.A(n_5157),
.B(n_378),
.Y(n_5282)
);

OAI33xp33_ASAP7_75t_L g5283 ( 
.A1(n_5171),
.A2(n_5138),
.A3(n_5125),
.B1(n_5089),
.B2(n_5094),
.B3(n_5108),
.Y(n_5283)
);

NAND4xp25_ASAP7_75t_L g5284 ( 
.A(n_5087),
.B(n_380),
.C(n_378),
.D(n_379),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_5084),
.Y(n_5285)
);

NAND2xp5_ASAP7_75t_L g5286 ( 
.A(n_5113),
.B(n_379),
.Y(n_5286)
);

AO21x2_ASAP7_75t_L g5287 ( 
.A1(n_5103),
.A2(n_5112),
.B(n_5099),
.Y(n_5287)
);

AND2x2_ASAP7_75t_L g5288 ( 
.A(n_5137),
.B(n_381),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_5086),
.Y(n_5289)
);

NAND2xp5_ASAP7_75t_L g5290 ( 
.A(n_5153),
.B(n_381),
.Y(n_5290)
);

NOR3xp33_ASAP7_75t_L g5291 ( 
.A(n_5185),
.B(n_381),
.C(n_382),
.Y(n_5291)
);

INVxp67_ASAP7_75t_L g5292 ( 
.A(n_5182),
.Y(n_5292)
);

INVx2_ASAP7_75t_SL g5293 ( 
.A(n_5208),
.Y(n_5293)
);

NAND4xp25_ASAP7_75t_SL g5294 ( 
.A(n_5177),
.B(n_384),
.C(n_382),
.D(n_383),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_5097),
.Y(n_5295)
);

INVx2_ASAP7_75t_L g5296 ( 
.A(n_5070),
.Y(n_5296)
);

INVx2_ASAP7_75t_L g5297 ( 
.A(n_5083),
.Y(n_5297)
);

INVx1_ASAP7_75t_L g5298 ( 
.A(n_5101),
.Y(n_5298)
);

AOI21xp5_ASAP7_75t_SL g5299 ( 
.A1(n_5130),
.A2(n_385),
.B(n_386),
.Y(n_5299)
);

INVx2_ASAP7_75t_L g5300 ( 
.A(n_5124),
.Y(n_5300)
);

OAI211xp5_ASAP7_75t_L g5301 ( 
.A1(n_5188),
.A2(n_394),
.B(n_400),
.C(n_385),
.Y(n_5301)
);

NAND2xp5_ASAP7_75t_L g5302 ( 
.A(n_5162),
.B(n_387),
.Y(n_5302)
);

AND2x2_ASAP7_75t_L g5303 ( 
.A(n_5139),
.B(n_387),
.Y(n_5303)
);

NAND4xp25_ASAP7_75t_L g5304 ( 
.A(n_5161),
.B(n_5059),
.C(n_5215),
.D(n_5197),
.Y(n_5304)
);

INVxp67_ASAP7_75t_SL g5305 ( 
.A(n_5228),
.Y(n_5305)
);

INVx1_ASAP7_75t_L g5306 ( 
.A(n_5106),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_5109),
.Y(n_5307)
);

AOI211xp5_ASAP7_75t_L g5308 ( 
.A1(n_5187),
.A2(n_390),
.B(n_388),
.C(n_389),
.Y(n_5308)
);

INVx1_ASAP7_75t_L g5309 ( 
.A(n_5193),
.Y(n_5309)
);

AOI22xp33_ASAP7_75t_L g5310 ( 
.A1(n_5178),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_5310)
);

AOI22xp5_ASAP7_75t_L g5311 ( 
.A1(n_5123),
.A2(n_391),
.B1(n_389),
.B2(n_390),
.Y(n_5311)
);

NAND4xp25_ASAP7_75t_L g5312 ( 
.A(n_5092),
.B(n_393),
.C(n_391),
.D(n_392),
.Y(n_5312)
);

AND2x2_ASAP7_75t_L g5313 ( 
.A(n_5148),
.B(n_392),
.Y(n_5313)
);

AOI22xp33_ASAP7_75t_L g5314 ( 
.A1(n_5181),
.A2(n_5173),
.B1(n_5186),
.B2(n_5183),
.Y(n_5314)
);

INVx2_ASAP7_75t_L g5315 ( 
.A(n_5114),
.Y(n_5315)
);

INVx4_ASAP7_75t_L g5316 ( 
.A(n_5072),
.Y(n_5316)
);

BUFx12f_ASAP7_75t_L g5317 ( 
.A(n_5158),
.Y(n_5317)
);

NAND2xp5_ASAP7_75t_L g5318 ( 
.A(n_5095),
.B(n_394),
.Y(n_5318)
);

INVx2_ASAP7_75t_SL g5319 ( 
.A(n_5216),
.Y(n_5319)
);

INVx1_ASAP7_75t_L g5320 ( 
.A(n_5201),
.Y(n_5320)
);

AND2x2_ASAP7_75t_L g5321 ( 
.A(n_5151),
.B(n_396),
.Y(n_5321)
);

INVx1_ASAP7_75t_L g5322 ( 
.A(n_5204),
.Y(n_5322)
);

NAND2xp5_ASAP7_75t_L g5323 ( 
.A(n_5115),
.B(n_396),
.Y(n_5323)
);

AND2x2_ASAP7_75t_L g5324 ( 
.A(n_5127),
.B(n_396),
.Y(n_5324)
);

AND2x4_ASAP7_75t_L g5325 ( 
.A(n_5168),
.B(n_397),
.Y(n_5325)
);

AOI22xp33_ASAP7_75t_L g5326 ( 
.A1(n_5119),
.A2(n_399),
.B1(n_397),
.B2(n_398),
.Y(n_5326)
);

INVx2_ASAP7_75t_L g5327 ( 
.A(n_5088),
.Y(n_5327)
);

INVx1_ASAP7_75t_L g5328 ( 
.A(n_5205),
.Y(n_5328)
);

INVx2_ASAP7_75t_L g5329 ( 
.A(n_5098),
.Y(n_5329)
);

OAI22xp5_ASAP7_75t_L g5330 ( 
.A1(n_5096),
.A2(n_403),
.B1(n_401),
.B2(n_402),
.Y(n_5330)
);

OAI33xp33_ASAP7_75t_L g5331 ( 
.A1(n_5129),
.A2(n_404),
.A3(n_403),
.B1(n_402),
.B2(n_405),
.B3(n_718),
.Y(n_5331)
);

OAI221xp5_ASAP7_75t_L g5332 ( 
.A1(n_5052),
.A2(n_405),
.B1(n_402),
.B2(n_403),
.C(n_719),
.Y(n_5332)
);

AOI21xp33_ASAP7_75t_L g5333 ( 
.A1(n_5062),
.A2(n_720),
.B(n_721),
.Y(n_5333)
);

AND2x2_ASAP7_75t_L g5334 ( 
.A(n_5136),
.B(n_722),
.Y(n_5334)
);

AND2x2_ASAP7_75t_L g5335 ( 
.A(n_5140),
.B(n_722),
.Y(n_5335)
);

OAI21x1_ASAP7_75t_L g5336 ( 
.A1(n_5102),
.A2(n_5105),
.B(n_5110),
.Y(n_5336)
);

AOI322xp5_ASAP7_75t_L g5337 ( 
.A1(n_5163),
.A2(n_728),
.A3(n_727),
.B1(n_725),
.B2(n_723),
.C1(n_724),
.C2(n_726),
.Y(n_5337)
);

INVx4_ASAP7_75t_L g5338 ( 
.A(n_5195),
.Y(n_5338)
);

NOR3xp33_ASAP7_75t_L g5339 ( 
.A(n_5065),
.B(n_726),
.C(n_727),
.Y(n_5339)
);

OAI322xp33_ASAP7_75t_SL g5340 ( 
.A1(n_5144),
.A2(n_733),
.A3(n_732),
.B1(n_730),
.B2(n_728),
.C1(n_729),
.C2(n_731),
.Y(n_5340)
);

INVx5_ASAP7_75t_L g5341 ( 
.A(n_5056),
.Y(n_5341)
);

AOI222xp33_ASAP7_75t_L g5342 ( 
.A1(n_5160),
.A2(n_732),
.B1(n_734),
.B2(n_730),
.C1(n_731),
.C2(n_733),
.Y(n_5342)
);

OAI21xp5_ASAP7_75t_SL g5343 ( 
.A1(n_5149),
.A2(n_736),
.B(n_735),
.Y(n_5343)
);

INVxp67_ASAP7_75t_L g5344 ( 
.A(n_5076),
.Y(n_5344)
);

AND2x4_ASAP7_75t_L g5345 ( 
.A(n_5075),
.B(n_738),
.Y(n_5345)
);

BUFx2_ASAP7_75t_L g5346 ( 
.A(n_5053),
.Y(n_5346)
);

NAND2xp5_ASAP7_75t_L g5347 ( 
.A(n_5104),
.B(n_739),
.Y(n_5347)
);

OAI33xp33_ASAP7_75t_L g5348 ( 
.A1(n_5189),
.A2(n_744),
.A3(n_746),
.B1(n_740),
.B2(n_743),
.B3(n_745),
.Y(n_5348)
);

INVx1_ASAP7_75t_L g5349 ( 
.A(n_5214),
.Y(n_5349)
);

INVx2_ASAP7_75t_L g5350 ( 
.A(n_5107),
.Y(n_5350)
);

OAI31xp33_ASAP7_75t_L g5351 ( 
.A1(n_5219),
.A2(n_1794),
.A3(n_1795),
.B(n_1793),
.Y(n_5351)
);

NAND3xp33_ASAP7_75t_SL g5352 ( 
.A(n_5141),
.B(n_743),
.C(n_746),
.Y(n_5352)
);

INVx2_ASAP7_75t_L g5353 ( 
.A(n_5220),
.Y(n_5353)
);

AND2x4_ASAP7_75t_L g5354 ( 
.A(n_5192),
.B(n_747),
.Y(n_5354)
);

INVx2_ASAP7_75t_L g5355 ( 
.A(n_5223),
.Y(n_5355)
);

INVx3_ASAP7_75t_L g5356 ( 
.A(n_5111),
.Y(n_5356)
);

NAND2xp5_ASAP7_75t_L g5357 ( 
.A(n_5090),
.B(n_750),
.Y(n_5357)
);

INVx2_ASAP7_75t_L g5358 ( 
.A(n_5224),
.Y(n_5358)
);

AND2x2_ASAP7_75t_L g5359 ( 
.A(n_5134),
.B(n_750),
.Y(n_5359)
);

NAND2xp5_ASAP7_75t_L g5360 ( 
.A(n_5091),
.B(n_751),
.Y(n_5360)
);

NOR2xp33_ASAP7_75t_L g5361 ( 
.A(n_5069),
.B(n_752),
.Y(n_5361)
);

OR2x2_ASAP7_75t_L g5362 ( 
.A(n_5230),
.B(n_753),
.Y(n_5362)
);

INVx2_ASAP7_75t_L g5363 ( 
.A(n_5232),
.Y(n_5363)
);

AND2x4_ASAP7_75t_L g5364 ( 
.A(n_5194),
.B(n_753),
.Y(n_5364)
);

INVx2_ASAP7_75t_SL g5365 ( 
.A(n_5199),
.Y(n_5365)
);

NAND2x1p5_ASAP7_75t_L g5366 ( 
.A(n_5240),
.B(n_5263),
.Y(n_5366)
);

OAI211xp5_ASAP7_75t_L g5367 ( 
.A1(n_5250),
.A2(n_5063),
.B(n_5147),
.C(n_5132),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_5272),
.Y(n_5368)
);

AND2x4_ASAP7_75t_L g5369 ( 
.A(n_5236),
.B(n_5200),
.Y(n_5369)
);

AND2x2_ASAP7_75t_L g5370 ( 
.A(n_5241),
.B(n_5159),
.Y(n_5370)
);

NOR2xp33_ASAP7_75t_L g5371 ( 
.A(n_5249),
.B(n_5067),
.Y(n_5371)
);

INVx1_ASAP7_75t_L g5372 ( 
.A(n_5279),
.Y(n_5372)
);

AND2x2_ASAP7_75t_L g5373 ( 
.A(n_5341),
.B(n_5346),
.Y(n_5373)
);

HB1xp67_ASAP7_75t_L g5374 ( 
.A(n_5341),
.Y(n_5374)
);

INVx4_ASAP7_75t_L g5375 ( 
.A(n_5278),
.Y(n_5375)
);

INVx1_ASAP7_75t_L g5376 ( 
.A(n_5353),
.Y(n_5376)
);

INVx2_ASAP7_75t_SL g5377 ( 
.A(n_5262),
.Y(n_5377)
);

AND2x2_ASAP7_75t_L g5378 ( 
.A(n_5341),
.B(n_5135),
.Y(n_5378)
);

OR2x2_ASAP7_75t_L g5379 ( 
.A(n_5267),
.B(n_5071),
.Y(n_5379)
);

INVx2_ASAP7_75t_L g5380 ( 
.A(n_5316),
.Y(n_5380)
);

INVx1_ASAP7_75t_SL g5381 ( 
.A(n_5317),
.Y(n_5381)
);

OR2x2_ASAP7_75t_L g5382 ( 
.A(n_5292),
.B(n_5212),
.Y(n_5382)
);

HB1xp67_ASAP7_75t_L g5383 ( 
.A(n_5365),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_5355),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_5358),
.Y(n_5385)
);

INVxp67_ASAP7_75t_SL g5386 ( 
.A(n_5271),
.Y(n_5386)
);

HB1xp67_ASAP7_75t_L g5387 ( 
.A(n_5287),
.Y(n_5387)
);

NAND2xp5_ASAP7_75t_L g5388 ( 
.A(n_5293),
.B(n_5202),
.Y(n_5388)
);

AND2x2_ASAP7_75t_L g5389 ( 
.A(n_5276),
.B(n_5209),
.Y(n_5389)
);

INVx2_ASAP7_75t_SL g5390 ( 
.A(n_5338),
.Y(n_5390)
);

INVx2_ASAP7_75t_L g5391 ( 
.A(n_5319),
.Y(n_5391)
);

INVx2_ASAP7_75t_L g5392 ( 
.A(n_5356),
.Y(n_5392)
);

INVx1_ASAP7_75t_SL g5393 ( 
.A(n_5242),
.Y(n_5393)
);

OR2x2_ASAP7_75t_L g5394 ( 
.A(n_5350),
.B(n_5221),
.Y(n_5394)
);

AOI22xp5_ASAP7_75t_L g5395 ( 
.A1(n_5252),
.A2(n_5233),
.B1(n_5210),
.B2(n_5213),
.Y(n_5395)
);

OAI31xp33_ASAP7_75t_L g5396 ( 
.A1(n_5301),
.A2(n_5180),
.A3(n_5176),
.B(n_5179),
.Y(n_5396)
);

AND2x2_ASAP7_75t_L g5397 ( 
.A(n_5258),
.B(n_5211),
.Y(n_5397)
);

OR2x2_ASAP7_75t_L g5398 ( 
.A(n_5259),
.B(n_5122),
.Y(n_5398)
);

OR2x2_ASAP7_75t_L g5399 ( 
.A(n_5315),
.B(n_5118),
.Y(n_5399)
);

AND2x2_ASAP7_75t_L g5400 ( 
.A(n_5265),
.B(n_5227),
.Y(n_5400)
);

INVx1_ASAP7_75t_L g5401 ( 
.A(n_5363),
.Y(n_5401)
);

NAND2xp5_ASAP7_75t_L g5402 ( 
.A(n_5314),
.B(n_5231),
.Y(n_5402)
);

NOR3xp33_ASAP7_75t_L g5403 ( 
.A(n_5238),
.B(n_5164),
.C(n_5058),
.Y(n_5403)
);

INVx6_ASAP7_75t_L g5404 ( 
.A(n_5325),
.Y(n_5404)
);

INVx2_ASAP7_75t_L g5405 ( 
.A(n_5336),
.Y(n_5405)
);

A2O1A1Ixp33_ASAP7_75t_L g5406 ( 
.A1(n_5268),
.A2(n_5172),
.B(n_5184),
.C(n_5174),
.Y(n_5406)
);

INVxp67_ASAP7_75t_L g5407 ( 
.A(n_5305),
.Y(n_5407)
);

INVx1_ASAP7_75t_L g5408 ( 
.A(n_5260),
.Y(n_5408)
);

BUFx3_ASAP7_75t_L g5409 ( 
.A(n_5345),
.Y(n_5409)
);

CKINVDCx5p33_ASAP7_75t_R g5410 ( 
.A(n_5299),
.Y(n_5410)
);

NAND2xp5_ASAP7_75t_L g5411 ( 
.A(n_5264),
.B(n_5085),
.Y(n_5411)
);

INVx1_ASAP7_75t_L g5412 ( 
.A(n_5266),
.Y(n_5412)
);

NOR2xp33_ASAP7_75t_L g5413 ( 
.A(n_5256),
.B(n_5093),
.Y(n_5413)
);

OR2x2_ASAP7_75t_L g5414 ( 
.A(n_5257),
.B(n_5081),
.Y(n_5414)
);

INVx2_ASAP7_75t_SL g5415 ( 
.A(n_5354),
.Y(n_5415)
);

INVx2_ASAP7_75t_L g5416 ( 
.A(n_5273),
.Y(n_5416)
);

AND2x2_ASAP7_75t_L g5417 ( 
.A(n_5344),
.B(n_5060),
.Y(n_5417)
);

AND2x2_ASAP7_75t_L g5418 ( 
.A(n_5300),
.B(n_5057),
.Y(n_5418)
);

BUFx3_ASAP7_75t_L g5419 ( 
.A(n_5364),
.Y(n_5419)
);

NAND2xp5_ASAP7_75t_L g5420 ( 
.A(n_5254),
.B(n_5131),
.Y(n_5420)
);

OR2x2_ASAP7_75t_L g5421 ( 
.A(n_5237),
.B(n_5155),
.Y(n_5421)
);

INVx1_ASAP7_75t_L g5422 ( 
.A(n_5280),
.Y(n_5422)
);

NAND2xp5_ASAP7_75t_L g5423 ( 
.A(n_5339),
.B(n_754),
.Y(n_5423)
);

INVx1_ASAP7_75t_L g5424 ( 
.A(n_5281),
.Y(n_5424)
);

AND2x2_ASAP7_75t_L g5425 ( 
.A(n_5359),
.B(n_755),
.Y(n_5425)
);

INVx1_ASAP7_75t_L g5426 ( 
.A(n_5285),
.Y(n_5426)
);

AND2x2_ASAP7_75t_L g5427 ( 
.A(n_5335),
.B(n_755),
.Y(n_5427)
);

NAND2xp5_ASAP7_75t_L g5428 ( 
.A(n_5282),
.B(n_756),
.Y(n_5428)
);

AOI32xp33_ASAP7_75t_L g5429 ( 
.A1(n_5291),
.A2(n_758),
.A3(n_756),
.B1(n_757),
.B2(n_759),
.Y(n_5429)
);

AND2x2_ASAP7_75t_L g5430 ( 
.A(n_5288),
.B(n_757),
.Y(n_5430)
);

NAND2xp5_ASAP7_75t_L g5431 ( 
.A(n_5343),
.B(n_758),
.Y(n_5431)
);

NAND2xp5_ASAP7_75t_L g5432 ( 
.A(n_5245),
.B(n_759),
.Y(n_5432)
);

INVx1_ASAP7_75t_SL g5433 ( 
.A(n_5270),
.Y(n_5433)
);

AND2x2_ASAP7_75t_L g5434 ( 
.A(n_5303),
.B(n_760),
.Y(n_5434)
);

INVx2_ASAP7_75t_L g5435 ( 
.A(n_5296),
.Y(n_5435)
);

NOR2xp33_ASAP7_75t_L g5436 ( 
.A(n_5283),
.B(n_761),
.Y(n_5436)
);

INVx1_ASAP7_75t_L g5437 ( 
.A(n_5289),
.Y(n_5437)
);

OR2x2_ASAP7_75t_L g5438 ( 
.A(n_5239),
.B(n_1796),
.Y(n_5438)
);

OR2x2_ASAP7_75t_L g5439 ( 
.A(n_5243),
.B(n_761),
.Y(n_5439)
);

AND2x2_ASAP7_75t_L g5440 ( 
.A(n_5324),
.B(n_762),
.Y(n_5440)
);

OR2x2_ASAP7_75t_L g5441 ( 
.A(n_5248),
.B(n_1779),
.Y(n_5441)
);

OR2x2_ASAP7_75t_L g5442 ( 
.A(n_5255),
.B(n_1779),
.Y(n_5442)
);

INVx2_ASAP7_75t_L g5443 ( 
.A(n_5297),
.Y(n_5443)
);

AND2x2_ASAP7_75t_L g5444 ( 
.A(n_5334),
.B(n_763),
.Y(n_5444)
);

AND2x2_ASAP7_75t_L g5445 ( 
.A(n_5327),
.B(n_5329),
.Y(n_5445)
);

OR2x2_ASAP7_75t_L g5446 ( 
.A(n_5286),
.B(n_1781),
.Y(n_5446)
);

INVx2_ASAP7_75t_L g5447 ( 
.A(n_5362),
.Y(n_5447)
);

NOR2xp33_ASAP7_75t_L g5448 ( 
.A(n_5304),
.B(n_764),
.Y(n_5448)
);

NAND2xp5_ASAP7_75t_L g5449 ( 
.A(n_5351),
.B(n_765),
.Y(n_5449)
);

INVx2_ASAP7_75t_L g5450 ( 
.A(n_5253),
.Y(n_5450)
);

OA21x2_ASAP7_75t_L g5451 ( 
.A1(n_5295),
.A2(n_5306),
.B(n_5298),
.Y(n_5451)
);

INVx1_ASAP7_75t_SL g5452 ( 
.A(n_5357),
.Y(n_5452)
);

NOR2xp33_ASAP7_75t_L g5453 ( 
.A(n_5269),
.B(n_766),
.Y(n_5453)
);

INVx2_ASAP7_75t_L g5454 ( 
.A(n_5321),
.Y(n_5454)
);

AND2x4_ASAP7_75t_L g5455 ( 
.A(n_5313),
.B(n_1784),
.Y(n_5455)
);

NAND4xp25_ASAP7_75t_L g5456 ( 
.A(n_5308),
.B(n_768),
.C(n_766),
.D(n_767),
.Y(n_5456)
);

BUFx2_ASAP7_75t_L g5457 ( 
.A(n_5274),
.Y(n_5457)
);

INVx1_ASAP7_75t_L g5458 ( 
.A(n_5307),
.Y(n_5458)
);

AND2x2_ASAP7_75t_L g5459 ( 
.A(n_5323),
.B(n_767),
.Y(n_5459)
);

INVx2_ASAP7_75t_L g5460 ( 
.A(n_5309),
.Y(n_5460)
);

AND2x2_ASAP7_75t_L g5461 ( 
.A(n_5389),
.B(n_5261),
.Y(n_5461)
);

AND2x2_ASAP7_75t_L g5462 ( 
.A(n_5381),
.B(n_5302),
.Y(n_5462)
);

AND2x2_ASAP7_75t_L g5463 ( 
.A(n_5390),
.B(n_5378),
.Y(n_5463)
);

INVx1_ASAP7_75t_L g5464 ( 
.A(n_5374),
.Y(n_5464)
);

HB1xp67_ASAP7_75t_L g5465 ( 
.A(n_5373),
.Y(n_5465)
);

INVx1_ASAP7_75t_L g5466 ( 
.A(n_5399),
.Y(n_5466)
);

AND2x2_ASAP7_75t_L g5467 ( 
.A(n_5370),
.B(n_5290),
.Y(n_5467)
);

NAND2xp5_ASAP7_75t_L g5468 ( 
.A(n_5377),
.B(n_5386),
.Y(n_5468)
);

INVx1_ASAP7_75t_L g5469 ( 
.A(n_5451),
.Y(n_5469)
);

AND2x2_ASAP7_75t_L g5470 ( 
.A(n_5380),
.B(n_5320),
.Y(n_5470)
);

AND2x2_ASAP7_75t_L g5471 ( 
.A(n_5369),
.B(n_5322),
.Y(n_5471)
);

AND2x2_ASAP7_75t_L g5472 ( 
.A(n_5366),
.B(n_5328),
.Y(n_5472)
);

NAND2x1p5_ASAP7_75t_L g5473 ( 
.A(n_5375),
.B(n_5277),
.Y(n_5473)
);

AOI21xp33_ASAP7_75t_SL g5474 ( 
.A1(n_5410),
.A2(n_5247),
.B(n_5342),
.Y(n_5474)
);

OAI21xp33_ASAP7_75t_L g5475 ( 
.A1(n_5407),
.A2(n_5284),
.B(n_5337),
.Y(n_5475)
);

AOI221x1_ASAP7_75t_L g5476 ( 
.A1(n_5436),
.A2(n_5330),
.B1(n_5333),
.B2(n_5312),
.C(n_5352),
.Y(n_5476)
);

INVx1_ASAP7_75t_L g5477 ( 
.A(n_5368),
.Y(n_5477)
);

AND2x2_ASAP7_75t_L g5478 ( 
.A(n_5397),
.B(n_5349),
.Y(n_5478)
);

INVx5_ASAP7_75t_L g5479 ( 
.A(n_5404),
.Y(n_5479)
);

INVx2_ASAP7_75t_L g5480 ( 
.A(n_5409),
.Y(n_5480)
);

NOR2xp33_ASAP7_75t_L g5481 ( 
.A(n_5413),
.B(n_5318),
.Y(n_5481)
);

INVx2_ASAP7_75t_L g5482 ( 
.A(n_5419),
.Y(n_5482)
);

NAND2xp5_ASAP7_75t_L g5483 ( 
.A(n_5415),
.B(n_5361),
.Y(n_5483)
);

NAND2xp5_ASAP7_75t_L g5484 ( 
.A(n_5406),
.B(n_5311),
.Y(n_5484)
);

AND2x2_ASAP7_75t_L g5485 ( 
.A(n_5400),
.B(n_5360),
.Y(n_5485)
);

INVx2_ASAP7_75t_L g5486 ( 
.A(n_5391),
.Y(n_5486)
);

AND2x2_ASAP7_75t_L g5487 ( 
.A(n_5392),
.B(n_5347),
.Y(n_5487)
);

INVx1_ASAP7_75t_L g5488 ( 
.A(n_5394),
.Y(n_5488)
);

AND2x2_ASAP7_75t_L g5489 ( 
.A(n_5417),
.B(n_5251),
.Y(n_5489)
);

OR2x2_ASAP7_75t_L g5490 ( 
.A(n_5433),
.B(n_5251),
.Y(n_5490)
);

AND2x2_ASAP7_75t_L g5491 ( 
.A(n_5418),
.B(n_5310),
.Y(n_5491)
);

AND2x2_ASAP7_75t_L g5492 ( 
.A(n_5383),
.B(n_5454),
.Y(n_5492)
);

NAND2xp5_ASAP7_75t_L g5493 ( 
.A(n_5395),
.B(n_5275),
.Y(n_5493)
);

NAND2xp5_ASAP7_75t_L g5494 ( 
.A(n_5411),
.B(n_5246),
.Y(n_5494)
);

NAND2xp5_ASAP7_75t_L g5495 ( 
.A(n_5452),
.B(n_5326),
.Y(n_5495)
);

NAND2xp5_ASAP7_75t_L g5496 ( 
.A(n_5371),
.B(n_5332),
.Y(n_5496)
);

NAND2xp5_ASAP7_75t_L g5497 ( 
.A(n_5457),
.B(n_5340),
.Y(n_5497)
);

AOI221xp5_ASAP7_75t_L g5498 ( 
.A1(n_5387),
.A2(n_5331),
.B1(n_5294),
.B2(n_5348),
.C(n_5244),
.Y(n_5498)
);

AND2x2_ASAP7_75t_L g5499 ( 
.A(n_5416),
.B(n_768),
.Y(n_5499)
);

INVx2_ASAP7_75t_L g5500 ( 
.A(n_5421),
.Y(n_5500)
);

INVx1_ASAP7_75t_L g5501 ( 
.A(n_5372),
.Y(n_5501)
);

AND2x2_ASAP7_75t_L g5502 ( 
.A(n_5450),
.B(n_769),
.Y(n_5502)
);

OR2x2_ASAP7_75t_L g5503 ( 
.A(n_5379),
.B(n_770),
.Y(n_5503)
);

AND2x4_ASAP7_75t_SL g5504 ( 
.A(n_5455),
.B(n_770),
.Y(n_5504)
);

NAND2xp5_ASAP7_75t_L g5505 ( 
.A(n_5396),
.B(n_771),
.Y(n_5505)
);

AND2x2_ASAP7_75t_L g5506 ( 
.A(n_5447),
.B(n_772),
.Y(n_5506)
);

AND2x2_ASAP7_75t_L g5507 ( 
.A(n_5388),
.B(n_5414),
.Y(n_5507)
);

AND2x2_ASAP7_75t_L g5508 ( 
.A(n_5420),
.B(n_5445),
.Y(n_5508)
);

INVx2_ASAP7_75t_L g5509 ( 
.A(n_5398),
.Y(n_5509)
);

INVx1_ASAP7_75t_L g5510 ( 
.A(n_5382),
.Y(n_5510)
);

AND3x2_ASAP7_75t_L g5511 ( 
.A(n_5448),
.B(n_773),
.C(n_774),
.Y(n_5511)
);

NAND2xp5_ASAP7_75t_L g5512 ( 
.A(n_5402),
.B(n_773),
.Y(n_5512)
);

INVx1_ASAP7_75t_L g5513 ( 
.A(n_5438),
.Y(n_5513)
);

NOR2xp33_ASAP7_75t_L g5514 ( 
.A(n_5367),
.B(n_1776),
.Y(n_5514)
);

AND2x2_ASAP7_75t_L g5515 ( 
.A(n_5459),
.B(n_775),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_5439),
.Y(n_5516)
);

INVx1_ASAP7_75t_L g5517 ( 
.A(n_5441),
.Y(n_5517)
);

AND2x2_ASAP7_75t_L g5518 ( 
.A(n_5425),
.B(n_776),
.Y(n_5518)
);

NAND2xp5_ASAP7_75t_SL g5519 ( 
.A(n_5429),
.B(n_776),
.Y(n_5519)
);

INVx2_ASAP7_75t_L g5520 ( 
.A(n_5405),
.Y(n_5520)
);

INVx1_ASAP7_75t_L g5521 ( 
.A(n_5442),
.Y(n_5521)
);

INVx1_ASAP7_75t_L g5522 ( 
.A(n_5376),
.Y(n_5522)
);

INVx1_ASAP7_75t_L g5523 ( 
.A(n_5384),
.Y(n_5523)
);

HB1xp67_ASAP7_75t_L g5524 ( 
.A(n_5435),
.Y(n_5524)
);

NAND2xp5_ASAP7_75t_L g5525 ( 
.A(n_5403),
.B(n_777),
.Y(n_5525)
);

NAND2xp5_ASAP7_75t_L g5526 ( 
.A(n_5443),
.B(n_777),
.Y(n_5526)
);

NAND2x1_ASAP7_75t_L g5527 ( 
.A(n_5460),
.B(n_779),
.Y(n_5527)
);

AND2x2_ASAP7_75t_L g5528 ( 
.A(n_5427),
.B(n_779),
.Y(n_5528)
);

AND2x2_ASAP7_75t_L g5529 ( 
.A(n_5444),
.B(n_780),
.Y(n_5529)
);

INVx1_ASAP7_75t_L g5530 ( 
.A(n_5385),
.Y(n_5530)
);

NAND2xp5_ASAP7_75t_L g5531 ( 
.A(n_5449),
.B(n_780),
.Y(n_5531)
);

OR2x2_ASAP7_75t_L g5532 ( 
.A(n_5401),
.B(n_781),
.Y(n_5532)
);

OAI21x1_ASAP7_75t_L g5533 ( 
.A1(n_5408),
.A2(n_782),
.B(n_783),
.Y(n_5533)
);

INVx2_ASAP7_75t_L g5534 ( 
.A(n_5446),
.Y(n_5534)
);

AND2x2_ASAP7_75t_L g5535 ( 
.A(n_5430),
.B(n_782),
.Y(n_5535)
);

AND2x4_ASAP7_75t_L g5536 ( 
.A(n_5434),
.B(n_783),
.Y(n_5536)
);

INVx1_ASAP7_75t_L g5537 ( 
.A(n_5412),
.Y(n_5537)
);

INVxp67_ASAP7_75t_L g5538 ( 
.A(n_5453),
.Y(n_5538)
);

OAI21xp33_ASAP7_75t_L g5539 ( 
.A1(n_5456),
.A2(n_784),
.B(n_785),
.Y(n_5539)
);

NOR2xp33_ASAP7_75t_L g5540 ( 
.A(n_5431),
.B(n_1793),
.Y(n_5540)
);

NAND2xp5_ASAP7_75t_L g5541 ( 
.A(n_5440),
.B(n_786),
.Y(n_5541)
);

OAI22xp5_ASAP7_75t_L g5542 ( 
.A1(n_5423),
.A2(n_789),
.B1(n_790),
.B2(n_788),
.Y(n_5542)
);

AND2x2_ASAP7_75t_L g5543 ( 
.A(n_5428),
.B(n_787),
.Y(n_5543)
);

INVxp67_ASAP7_75t_L g5544 ( 
.A(n_5432),
.Y(n_5544)
);

INVx2_ASAP7_75t_L g5545 ( 
.A(n_5422),
.Y(n_5545)
);

INVx1_ASAP7_75t_SL g5546 ( 
.A(n_5424),
.Y(n_5546)
);

AND2x4_ASAP7_75t_L g5547 ( 
.A(n_5426),
.B(n_789),
.Y(n_5547)
);

OAI21xp33_ASAP7_75t_L g5548 ( 
.A1(n_5437),
.A2(n_791),
.B(n_792),
.Y(n_5548)
);

INVx1_ASAP7_75t_L g5549 ( 
.A(n_5458),
.Y(n_5549)
);

AND2x4_ASAP7_75t_L g5550 ( 
.A(n_5390),
.B(n_791),
.Y(n_5550)
);

OR3x2_ASAP7_75t_L g5551 ( 
.A(n_5456),
.B(n_792),
.C(n_793),
.Y(n_5551)
);

NOR2x1_ASAP7_75t_L g5552 ( 
.A(n_5380),
.B(n_793),
.Y(n_5552)
);

OR2x2_ASAP7_75t_L g5553 ( 
.A(n_5393),
.B(n_795),
.Y(n_5553)
);

NAND2xp5_ASAP7_75t_L g5554 ( 
.A(n_5377),
.B(n_795),
.Y(n_5554)
);

OR2x2_ASAP7_75t_L g5555 ( 
.A(n_5393),
.B(n_796),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_5464),
.Y(n_5556)
);

NAND2x1_ASAP7_75t_L g5557 ( 
.A(n_5552),
.B(n_796),
.Y(n_5557)
);

INVx4_ASAP7_75t_L g5558 ( 
.A(n_5479),
.Y(n_5558)
);

AND2x2_ASAP7_75t_L g5559 ( 
.A(n_5463),
.B(n_1786),
.Y(n_5559)
);

NAND2x1p5_ASAP7_75t_L g5560 ( 
.A(n_5479),
.B(n_797),
.Y(n_5560)
);

INVx1_ASAP7_75t_L g5561 ( 
.A(n_5502),
.Y(n_5561)
);

INVx2_ASAP7_75t_L g5562 ( 
.A(n_5479),
.Y(n_5562)
);

AOI22xp5_ASAP7_75t_L g5563 ( 
.A1(n_5514),
.A2(n_801),
.B1(n_798),
.B2(n_799),
.Y(n_5563)
);

AOI322xp5_ASAP7_75t_L g5564 ( 
.A1(n_5484),
.A2(n_807),
.A3(n_806),
.B1(n_803),
.B2(n_801),
.C1(n_802),
.C2(n_804),
.Y(n_5564)
);

OAI32xp33_ASAP7_75t_L g5565 ( 
.A1(n_5497),
.A2(n_806),
.A3(n_802),
.B1(n_803),
.B2(n_808),
.Y(n_5565)
);

INVx1_ASAP7_75t_L g5566 ( 
.A(n_5506),
.Y(n_5566)
);

AOI31xp33_ASAP7_75t_L g5567 ( 
.A1(n_5473),
.A2(n_811),
.A3(n_808),
.B(n_810),
.Y(n_5567)
);

INVx1_ASAP7_75t_L g5568 ( 
.A(n_5509),
.Y(n_5568)
);

INVx1_ASAP7_75t_L g5569 ( 
.A(n_5469),
.Y(n_5569)
);

HB1xp67_ASAP7_75t_L g5570 ( 
.A(n_5465),
.Y(n_5570)
);

INVx1_ASAP7_75t_L g5571 ( 
.A(n_5532),
.Y(n_5571)
);

AOI22xp5_ASAP7_75t_L g5572 ( 
.A1(n_5475),
.A2(n_812),
.B1(n_810),
.B2(n_811),
.Y(n_5572)
);

NAND2xp5_ASAP7_75t_L g5573 ( 
.A(n_5511),
.B(n_812),
.Y(n_5573)
);

INVx1_ASAP7_75t_SL g5574 ( 
.A(n_5504),
.Y(n_5574)
);

NAND2xp5_ASAP7_75t_L g5575 ( 
.A(n_5498),
.B(n_814),
.Y(n_5575)
);

INVx1_ASAP7_75t_L g5576 ( 
.A(n_5499),
.Y(n_5576)
);

INVx1_ASAP7_75t_L g5577 ( 
.A(n_5500),
.Y(n_5577)
);

NAND2xp5_ASAP7_75t_L g5578 ( 
.A(n_5480),
.B(n_814),
.Y(n_5578)
);

INVx1_ASAP7_75t_L g5579 ( 
.A(n_5488),
.Y(n_5579)
);

NAND2xp5_ASAP7_75t_L g5580 ( 
.A(n_5482),
.B(n_816),
.Y(n_5580)
);

INVx1_ASAP7_75t_SL g5581 ( 
.A(n_5472),
.Y(n_5581)
);

NAND2xp5_ASAP7_75t_L g5582 ( 
.A(n_5489),
.B(n_817),
.Y(n_5582)
);

AOI322xp5_ASAP7_75t_L g5583 ( 
.A1(n_5494),
.A2(n_822),
.A3(n_821),
.B1(n_819),
.B2(n_817),
.C1(n_818),
.C2(n_820),
.Y(n_5583)
);

NAND2xp5_ASAP7_75t_SL g5584 ( 
.A(n_5474),
.B(n_819),
.Y(n_5584)
);

INVx1_ASAP7_75t_L g5585 ( 
.A(n_5553),
.Y(n_5585)
);

AOI21xp33_ASAP7_75t_SL g5586 ( 
.A1(n_5519),
.A2(n_1775),
.B(n_1774),
.Y(n_5586)
);

INVx1_ASAP7_75t_L g5587 ( 
.A(n_5555),
.Y(n_5587)
);

AND2x2_ASAP7_75t_L g5588 ( 
.A(n_5462),
.B(n_1776),
.Y(n_5588)
);

INVx1_ASAP7_75t_SL g5589 ( 
.A(n_5550),
.Y(n_5589)
);

OR2x2_ASAP7_75t_L g5590 ( 
.A(n_5468),
.B(n_825),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_5503),
.Y(n_5591)
);

NAND2x1p5_ASAP7_75t_L g5592 ( 
.A(n_5527),
.B(n_828),
.Y(n_5592)
);

INVx1_ASAP7_75t_L g5593 ( 
.A(n_5526),
.Y(n_5593)
);

BUFx2_ASAP7_75t_L g5594 ( 
.A(n_5492),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_5510),
.Y(n_5595)
);

OAI21xp33_ASAP7_75t_SL g5596 ( 
.A1(n_5490),
.A2(n_829),
.B(n_830),
.Y(n_5596)
);

AOI211xp5_ASAP7_75t_L g5597 ( 
.A1(n_5493),
.A2(n_834),
.B(n_832),
.C(n_833),
.Y(n_5597)
);

AND2x2_ASAP7_75t_L g5598 ( 
.A(n_5508),
.B(n_1767),
.Y(n_5598)
);

INVxp67_ASAP7_75t_L g5599 ( 
.A(n_5481),
.Y(n_5599)
);

OAI32xp33_ASAP7_75t_L g5600 ( 
.A1(n_5505),
.A2(n_840),
.A3(n_836),
.B1(n_839),
.B2(n_841),
.Y(n_5600)
);

NAND2xp5_ASAP7_75t_L g5601 ( 
.A(n_5461),
.B(n_841),
.Y(n_5601)
);

INVx2_ASAP7_75t_L g5602 ( 
.A(n_5486),
.Y(n_5602)
);

NAND2xp5_ASAP7_75t_L g5603 ( 
.A(n_5491),
.B(n_842),
.Y(n_5603)
);

INVx1_ASAP7_75t_L g5604 ( 
.A(n_5513),
.Y(n_5604)
);

NAND2xp5_ASAP7_75t_L g5605 ( 
.A(n_5485),
.B(n_5467),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_5516),
.Y(n_5606)
);

INVx2_ASAP7_75t_L g5607 ( 
.A(n_5478),
.Y(n_5607)
);

INVx1_ASAP7_75t_L g5608 ( 
.A(n_5517),
.Y(n_5608)
);

AOI22xp5_ASAP7_75t_L g5609 ( 
.A1(n_5551),
.A2(n_846),
.B1(n_844),
.B2(n_845),
.Y(n_5609)
);

AOI32xp33_ASAP7_75t_L g5610 ( 
.A1(n_5525),
.A2(n_847),
.A3(n_845),
.B1(n_846),
.B2(n_848),
.Y(n_5610)
);

AOI22xp5_ASAP7_75t_L g5611 ( 
.A1(n_5496),
.A2(n_849),
.B1(n_847),
.B2(n_848),
.Y(n_5611)
);

NOR2xp33_ASAP7_75t_L g5612 ( 
.A(n_5538),
.B(n_1768),
.Y(n_5612)
);

OAI31xp33_ASAP7_75t_L g5613 ( 
.A1(n_5539),
.A2(n_852),
.A3(n_850),
.B(n_851),
.Y(n_5613)
);

NAND2xp5_ASAP7_75t_L g5614 ( 
.A(n_5507),
.B(n_850),
.Y(n_5614)
);

AOI21xp5_ASAP7_75t_L g5615 ( 
.A1(n_5476),
.A2(n_851),
.B(n_852),
.Y(n_5615)
);

NAND2xp5_ASAP7_75t_L g5616 ( 
.A(n_5487),
.B(n_853),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_5521),
.Y(n_5617)
);

OA21x2_ASAP7_75t_L g5618 ( 
.A1(n_5512),
.A2(n_854),
.B(n_856),
.Y(n_5618)
);

INVx1_ASAP7_75t_L g5619 ( 
.A(n_5466),
.Y(n_5619)
);

A2O1A1Ixp33_ASAP7_75t_L g5620 ( 
.A1(n_5548),
.A2(n_5540),
.B(n_5495),
.C(n_5542),
.Y(n_5620)
);

AND2x4_ASAP7_75t_L g5621 ( 
.A(n_5471),
.B(n_854),
.Y(n_5621)
);

OAI21xp33_ASAP7_75t_L g5622 ( 
.A1(n_5483),
.A2(n_856),
.B(n_857),
.Y(n_5622)
);

AND2x4_ASAP7_75t_L g5623 ( 
.A(n_5470),
.B(n_858),
.Y(n_5623)
);

NAND2xp5_ASAP7_75t_L g5624 ( 
.A(n_5534),
.B(n_858),
.Y(n_5624)
);

AOI21xp5_ASAP7_75t_L g5625 ( 
.A1(n_5531),
.A2(n_859),
.B(n_860),
.Y(n_5625)
);

NOR2xp33_ASAP7_75t_L g5626 ( 
.A(n_5554),
.B(n_1789),
.Y(n_5626)
);

NAND3xp33_ASAP7_75t_L g5627 ( 
.A(n_5477),
.B(n_859),
.C(n_860),
.Y(n_5627)
);

INVx1_ASAP7_75t_SL g5628 ( 
.A(n_5535),
.Y(n_5628)
);

OAI32xp33_ASAP7_75t_L g5629 ( 
.A1(n_5546),
.A2(n_863),
.A3(n_861),
.B1(n_862),
.B2(n_864),
.Y(n_5629)
);

INVx1_ASAP7_75t_SL g5630 ( 
.A(n_5518),
.Y(n_5630)
);

INVx1_ASAP7_75t_L g5631 ( 
.A(n_5524),
.Y(n_5631)
);

AOI222xp33_ASAP7_75t_L g5632 ( 
.A1(n_5544),
.A2(n_864),
.B1(n_866),
.B2(n_867),
.C1(n_862),
.C2(n_865),
.Y(n_5632)
);

INVx1_ASAP7_75t_L g5633 ( 
.A(n_5541),
.Y(n_5633)
);

INVx1_ASAP7_75t_L g5634 ( 
.A(n_5501),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_5529),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_5543),
.Y(n_5636)
);

INVx2_ASAP7_75t_L g5637 ( 
.A(n_5536),
.Y(n_5637)
);

AOI22xp5_ASAP7_75t_L g5638 ( 
.A1(n_5520),
.A2(n_870),
.B1(n_868),
.B2(n_869),
.Y(n_5638)
);

NOR2xp33_ASAP7_75t_L g5639 ( 
.A(n_5515),
.B(n_1770),
.Y(n_5639)
);

HB1xp67_ASAP7_75t_L g5640 ( 
.A(n_5533),
.Y(n_5640)
);

INVx1_ASAP7_75t_L g5641 ( 
.A(n_5528),
.Y(n_5641)
);

INVx2_ASAP7_75t_L g5642 ( 
.A(n_5547),
.Y(n_5642)
);

NAND3xp33_ASAP7_75t_L g5643 ( 
.A(n_5522),
.B(n_869),
.C(n_870),
.Y(n_5643)
);

NAND2xp5_ASAP7_75t_L g5644 ( 
.A(n_5523),
.B(n_871),
.Y(n_5644)
);

INVx1_ASAP7_75t_L g5645 ( 
.A(n_5537),
.Y(n_5645)
);

AO22x1_ASAP7_75t_L g5646 ( 
.A1(n_5545),
.A2(n_874),
.B1(n_872),
.B2(n_873),
.Y(n_5646)
);

OAI21xp33_ASAP7_75t_L g5647 ( 
.A1(n_5530),
.A2(n_874),
.B(n_875),
.Y(n_5647)
);

NAND2x2_ASAP7_75t_L g5648 ( 
.A(n_5549),
.B(n_875),
.Y(n_5648)
);

OAI22xp33_ASAP7_75t_L g5649 ( 
.A1(n_5497),
.A2(n_878),
.B1(n_876),
.B2(n_877),
.Y(n_5649)
);

INVx1_ASAP7_75t_L g5650 ( 
.A(n_5464),
.Y(n_5650)
);

INVx1_ASAP7_75t_L g5651 ( 
.A(n_5464),
.Y(n_5651)
);

INVx2_ASAP7_75t_L g5652 ( 
.A(n_5479),
.Y(n_5652)
);

INVx1_ASAP7_75t_L g5653 ( 
.A(n_5464),
.Y(n_5653)
);

OAI22xp5_ASAP7_75t_L g5654 ( 
.A1(n_5498),
.A2(n_881),
.B1(n_882),
.B2(n_880),
.Y(n_5654)
);

A2O1A1Ixp33_ASAP7_75t_L g5655 ( 
.A1(n_5615),
.A2(n_883),
.B(n_880),
.C(n_881),
.Y(n_5655)
);

AND2x2_ASAP7_75t_L g5656 ( 
.A(n_5581),
.B(n_885),
.Y(n_5656)
);

NOR2xp33_ASAP7_75t_L g5657 ( 
.A(n_5558),
.B(n_5567),
.Y(n_5657)
);

NAND2xp5_ASAP7_75t_SL g5658 ( 
.A(n_5596),
.B(n_886),
.Y(n_5658)
);

INVx1_ASAP7_75t_L g5659 ( 
.A(n_5560),
.Y(n_5659)
);

O2A1O1Ixp33_ASAP7_75t_L g5660 ( 
.A1(n_5654),
.A2(n_5584),
.B(n_5575),
.C(n_5649),
.Y(n_5660)
);

OR2x2_ASAP7_75t_L g5661 ( 
.A(n_5628),
.B(n_5630),
.Y(n_5661)
);

NAND2xp5_ASAP7_75t_L g5662 ( 
.A(n_5559),
.B(n_887),
.Y(n_5662)
);

AOI322xp5_ASAP7_75t_L g5663 ( 
.A1(n_5620),
.A2(n_894),
.A3(n_893),
.B1(n_891),
.B2(n_889),
.C1(n_890),
.C2(n_892),
.Y(n_5663)
);

INVx1_ASAP7_75t_SL g5664 ( 
.A(n_5592),
.Y(n_5664)
);

AOI22xp5_ASAP7_75t_L g5665 ( 
.A1(n_5572),
.A2(n_893),
.B1(n_891),
.B2(n_892),
.Y(n_5665)
);

OAI22xp5_ASAP7_75t_L g5666 ( 
.A1(n_5609),
.A2(n_897),
.B1(n_895),
.B2(n_896),
.Y(n_5666)
);

NAND2xp5_ASAP7_75t_L g5667 ( 
.A(n_5588),
.B(n_895),
.Y(n_5667)
);

AND2x2_ASAP7_75t_L g5668 ( 
.A(n_5637),
.B(n_899),
.Y(n_5668)
);

NAND2xp5_ASAP7_75t_L g5669 ( 
.A(n_5562),
.B(n_901),
.Y(n_5669)
);

OAI21xp33_ASAP7_75t_SL g5670 ( 
.A1(n_5569),
.A2(n_902),
.B(n_903),
.Y(n_5670)
);

INVx1_ASAP7_75t_L g5671 ( 
.A(n_5635),
.Y(n_5671)
);

INVx1_ASAP7_75t_SL g5672 ( 
.A(n_5573),
.Y(n_5672)
);

OAI32xp33_ASAP7_75t_L g5673 ( 
.A1(n_5640),
.A2(n_906),
.A3(n_908),
.B1(n_905),
.B2(n_907),
.Y(n_5673)
);

NAND2xp5_ASAP7_75t_L g5674 ( 
.A(n_5652),
.B(n_904),
.Y(n_5674)
);

NOR3xp33_ASAP7_75t_L g5675 ( 
.A(n_5599),
.B(n_910),
.C(n_911),
.Y(n_5675)
);

OAI221xp5_ASAP7_75t_L g5676 ( 
.A1(n_5613),
.A2(n_914),
.B1(n_911),
.B2(n_913),
.C(n_915),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_5641),
.Y(n_5677)
);

INVx2_ASAP7_75t_SL g5678 ( 
.A(n_5621),
.Y(n_5678)
);

AOI21xp5_ASAP7_75t_SL g5679 ( 
.A1(n_5618),
.A2(n_916),
.B(n_917),
.Y(n_5679)
);

AOI21xp5_ASAP7_75t_L g5680 ( 
.A1(n_5625),
.A2(n_916),
.B(n_917),
.Y(n_5680)
);

OAI22xp5_ASAP7_75t_L g5681 ( 
.A1(n_5563),
.A2(n_920),
.B1(n_918),
.B2(n_919),
.Y(n_5681)
);

NAND2xp5_ASAP7_75t_L g5682 ( 
.A(n_5598),
.B(n_918),
.Y(n_5682)
);

NAND2xp5_ASAP7_75t_L g5683 ( 
.A(n_5642),
.B(n_920),
.Y(n_5683)
);

AND2x4_ASAP7_75t_L g5684 ( 
.A(n_5631),
.B(n_5607),
.Y(n_5684)
);

INVx2_ASAP7_75t_L g5685 ( 
.A(n_5623),
.Y(n_5685)
);

INVx2_ASAP7_75t_L g5686 ( 
.A(n_5636),
.Y(n_5686)
);

OAI221xp5_ASAP7_75t_L g5687 ( 
.A1(n_5610),
.A2(n_925),
.B1(n_922),
.B2(n_924),
.C(n_926),
.Y(n_5687)
);

OAI31xp33_ASAP7_75t_L g5688 ( 
.A1(n_5627),
.A2(n_926),
.A3(n_924),
.B(n_925),
.Y(n_5688)
);

OAI21xp5_ASAP7_75t_L g5689 ( 
.A1(n_5582),
.A2(n_927),
.B(n_928),
.Y(n_5689)
);

OAI21xp33_ASAP7_75t_SL g5690 ( 
.A1(n_5605),
.A2(n_929),
.B(n_931),
.Y(n_5690)
);

AOI22xp5_ASAP7_75t_L g5691 ( 
.A1(n_5568),
.A2(n_5577),
.B1(n_5561),
.B2(n_5566),
.Y(n_5691)
);

INVx2_ASAP7_75t_SL g5692 ( 
.A(n_5648),
.Y(n_5692)
);

AND2x2_ASAP7_75t_L g5693 ( 
.A(n_5576),
.B(n_933),
.Y(n_5693)
);

INVx1_ASAP7_75t_L g5694 ( 
.A(n_5556),
.Y(n_5694)
);

NAND3xp33_ASAP7_75t_L g5695 ( 
.A(n_5650),
.B(n_5653),
.C(n_5651),
.Y(n_5695)
);

AOI22xp5_ASAP7_75t_L g5696 ( 
.A1(n_5585),
.A2(n_5587),
.B1(n_5595),
.B2(n_5579),
.Y(n_5696)
);

INVx1_ASAP7_75t_L g5697 ( 
.A(n_5591),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_5578),
.Y(n_5698)
);

INVx1_ASAP7_75t_L g5699 ( 
.A(n_5580),
.Y(n_5699)
);

AND2x2_ASAP7_75t_L g5700 ( 
.A(n_5571),
.B(n_934),
.Y(n_5700)
);

AOI21xp5_ASAP7_75t_L g5701 ( 
.A1(n_5603),
.A2(n_935),
.B(n_936),
.Y(n_5701)
);

OAI22xp5_ASAP7_75t_L g5702 ( 
.A1(n_5597),
.A2(n_937),
.B1(n_935),
.B2(n_936),
.Y(n_5702)
);

OAI22xp5_ASAP7_75t_L g5703 ( 
.A1(n_5611),
.A2(n_943),
.B1(n_941),
.B2(n_942),
.Y(n_5703)
);

AND2x2_ASAP7_75t_L g5704 ( 
.A(n_5633),
.B(n_942),
.Y(n_5704)
);

AOI21xp33_ASAP7_75t_SL g5705 ( 
.A1(n_5618),
.A2(n_943),
.B(n_944),
.Y(n_5705)
);

INVx2_ASAP7_75t_L g5706 ( 
.A(n_5590),
.Y(n_5706)
);

INVx1_ASAP7_75t_L g5707 ( 
.A(n_5624),
.Y(n_5707)
);

INVx1_ASAP7_75t_L g5708 ( 
.A(n_5619),
.Y(n_5708)
);

INVx1_ASAP7_75t_L g5709 ( 
.A(n_5616),
.Y(n_5709)
);

INVx2_ASAP7_75t_L g5710 ( 
.A(n_5602),
.Y(n_5710)
);

NOR3xp33_ASAP7_75t_L g5711 ( 
.A(n_5593),
.B(n_5606),
.C(n_5604),
.Y(n_5711)
);

AOI22xp5_ASAP7_75t_L g5712 ( 
.A1(n_5608),
.A2(n_5617),
.B1(n_5632),
.B2(n_5614),
.Y(n_5712)
);

INVx1_ASAP7_75t_L g5713 ( 
.A(n_5644),
.Y(n_5713)
);

AOI22xp5_ASAP7_75t_L g5714 ( 
.A1(n_5622),
.A2(n_5612),
.B1(n_5643),
.B2(n_5601),
.Y(n_5714)
);

NAND2xp5_ASAP7_75t_L g5715 ( 
.A(n_5586),
.B(n_948),
.Y(n_5715)
);

A2O1A1Ixp33_ASAP7_75t_L g5716 ( 
.A1(n_5564),
.A2(n_952),
.B(n_950),
.C(n_951),
.Y(n_5716)
);

OAI211xp5_ASAP7_75t_L g5717 ( 
.A1(n_5583),
.A2(n_5565),
.B(n_5600),
.C(n_5629),
.Y(n_5717)
);

INVx2_ASAP7_75t_L g5718 ( 
.A(n_5634),
.Y(n_5718)
);

AND2x2_ASAP7_75t_L g5719 ( 
.A(n_5639),
.B(n_953),
.Y(n_5719)
);

INVx1_ASAP7_75t_L g5720 ( 
.A(n_5646),
.Y(n_5720)
);

OAI211xp5_ASAP7_75t_L g5721 ( 
.A1(n_5638),
.A2(n_5647),
.B(n_5645),
.C(n_5626),
.Y(n_5721)
);

INVx1_ASAP7_75t_L g5722 ( 
.A(n_5570),
.Y(n_5722)
);

AOI222xp33_ASAP7_75t_L g5723 ( 
.A1(n_5584),
.A2(n_985),
.B1(n_965),
.B2(n_992),
.C1(n_976),
.C2(n_956),
.Y(n_5723)
);

AND2x4_ASAP7_75t_L g5724 ( 
.A(n_5558),
.B(n_958),
.Y(n_5724)
);

AOI22xp33_ASAP7_75t_SL g5725 ( 
.A1(n_5654),
.A2(n_960),
.B1(n_958),
.B2(n_959),
.Y(n_5725)
);

AOI322xp5_ASAP7_75t_L g5726 ( 
.A1(n_5584),
.A2(n_966),
.A3(n_965),
.B1(n_962),
.B2(n_959),
.C1(n_961),
.C2(n_964),
.Y(n_5726)
);

NAND2xp5_ASAP7_75t_L g5727 ( 
.A(n_5574),
.B(n_961),
.Y(n_5727)
);

NAND2x1_ASAP7_75t_SL g5728 ( 
.A(n_5558),
.B(n_962),
.Y(n_5728)
);

OR2x2_ASAP7_75t_L g5729 ( 
.A(n_5589),
.B(n_964),
.Y(n_5729)
);

OAI21xp5_ASAP7_75t_L g5730 ( 
.A1(n_5615),
.A2(n_966),
.B(n_968),
.Y(n_5730)
);

OAI21xp33_ASAP7_75t_SL g5731 ( 
.A1(n_5584),
.A2(n_968),
.B(n_969),
.Y(n_5731)
);

BUFx2_ASAP7_75t_L g5732 ( 
.A(n_5558),
.Y(n_5732)
);

INVx1_ASAP7_75t_L g5733 ( 
.A(n_5570),
.Y(n_5733)
);

AND2x2_ASAP7_75t_L g5734 ( 
.A(n_5594),
.B(n_969),
.Y(n_5734)
);

BUFx2_ASAP7_75t_SL g5735 ( 
.A(n_5558),
.Y(n_5735)
);

OAI211xp5_ASAP7_75t_SL g5736 ( 
.A1(n_5584),
.A2(n_973),
.B(n_970),
.C(n_972),
.Y(n_5736)
);

INVxp33_ASAP7_75t_L g5737 ( 
.A(n_5557),
.Y(n_5737)
);

OAI21xp5_ASAP7_75t_SL g5738 ( 
.A1(n_5615),
.A2(n_1772),
.B(n_1771),
.Y(n_5738)
);

INVx1_ASAP7_75t_L g5739 ( 
.A(n_5570),
.Y(n_5739)
);

NOR2xp33_ASAP7_75t_L g5740 ( 
.A(n_5558),
.B(n_978),
.Y(n_5740)
);

NAND2xp5_ASAP7_75t_SL g5741 ( 
.A(n_5558),
.B(n_979),
.Y(n_5741)
);

OAI22x1_ASAP7_75t_L g5742 ( 
.A1(n_5609),
.A2(n_982),
.B1(n_980),
.B2(n_981),
.Y(n_5742)
);

NOR2xp33_ASAP7_75t_L g5743 ( 
.A(n_5558),
.B(n_980),
.Y(n_5743)
);

NAND2xp5_ASAP7_75t_L g5744 ( 
.A(n_5574),
.B(n_981),
.Y(n_5744)
);

AOI22xp5_ASAP7_75t_L g5745 ( 
.A1(n_5654),
.A2(n_985),
.B1(n_983),
.B2(n_984),
.Y(n_5745)
);

AOI22xp33_ASAP7_75t_SL g5746 ( 
.A1(n_5654),
.A2(n_987),
.B1(n_983),
.B2(n_986),
.Y(n_5746)
);

NAND2xp5_ASAP7_75t_SL g5747 ( 
.A(n_5558),
.B(n_986),
.Y(n_5747)
);

AOI222xp33_ASAP7_75t_L g5748 ( 
.A1(n_5584),
.A2(n_1009),
.B1(n_994),
.B2(n_1018),
.C1(n_1001),
.C2(n_987),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_5570),
.Y(n_5749)
);

INVx1_ASAP7_75t_L g5750 ( 
.A(n_5570),
.Y(n_5750)
);

AND2x2_ASAP7_75t_L g5751 ( 
.A(n_5594),
.B(n_993),
.Y(n_5751)
);

OAI22xp33_ASAP7_75t_L g5752 ( 
.A1(n_5609),
.A2(n_997),
.B1(n_995),
.B2(n_996),
.Y(n_5752)
);

CKINVDCx14_ASAP7_75t_R g5753 ( 
.A(n_5594),
.Y(n_5753)
);

INVx1_ASAP7_75t_L g5754 ( 
.A(n_5570),
.Y(n_5754)
);

INVx1_ASAP7_75t_L g5755 ( 
.A(n_5570),
.Y(n_5755)
);

INVx2_ASAP7_75t_L g5756 ( 
.A(n_5560),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_5570),
.Y(n_5757)
);

AOI22xp33_ASAP7_75t_L g5758 ( 
.A1(n_5584),
.A2(n_1000),
.B1(n_998),
.B2(n_999),
.Y(n_5758)
);

INVx1_ASAP7_75t_SL g5759 ( 
.A(n_5594),
.Y(n_5759)
);

NAND2xp5_ASAP7_75t_L g5760 ( 
.A(n_5574),
.B(n_1002),
.Y(n_5760)
);

INVx2_ASAP7_75t_L g5761 ( 
.A(n_5560),
.Y(n_5761)
);

AOI22xp5_ASAP7_75t_L g5762 ( 
.A1(n_5654),
.A2(n_1005),
.B1(n_1003),
.B2(n_1004),
.Y(n_5762)
);

AOI22xp33_ASAP7_75t_L g5763 ( 
.A1(n_5584),
.A2(n_1007),
.B1(n_1005),
.B2(n_1006),
.Y(n_5763)
);

OR2x2_ASAP7_75t_L g5764 ( 
.A(n_5589),
.B(n_1009),
.Y(n_5764)
);

HB1xp67_ASAP7_75t_L g5765 ( 
.A(n_5570),
.Y(n_5765)
);

OAI22xp5_ASAP7_75t_L g5766 ( 
.A1(n_5609),
.A2(n_1012),
.B1(n_1010),
.B2(n_1011),
.Y(n_5766)
);

INVx1_ASAP7_75t_L g5767 ( 
.A(n_5570),
.Y(n_5767)
);

OAI21xp33_ASAP7_75t_SL g5768 ( 
.A1(n_5584),
.A2(n_1013),
.B(n_1014),
.Y(n_5768)
);

AOI222xp33_ASAP7_75t_L g5769 ( 
.A1(n_5584),
.A2(n_1042),
.B1(n_1026),
.B2(n_1050),
.C1(n_1034),
.C2(n_1013),
.Y(n_5769)
);

O2A1O1Ixp33_ASAP7_75t_L g5770 ( 
.A1(n_5615),
.A2(n_1762),
.B(n_1763),
.C(n_1761),
.Y(n_5770)
);

INVx3_ASAP7_75t_L g5771 ( 
.A(n_5558),
.Y(n_5771)
);

INVx1_ASAP7_75t_SL g5772 ( 
.A(n_5594),
.Y(n_5772)
);

NAND2xp5_ASAP7_75t_L g5773 ( 
.A(n_5574),
.B(n_1014),
.Y(n_5773)
);

AOI21xp5_ASAP7_75t_SL g5774 ( 
.A1(n_5567),
.A2(n_1015),
.B(n_1019),
.Y(n_5774)
);

AOI22xp5_ASAP7_75t_L g5775 ( 
.A1(n_5654),
.A2(n_1020),
.B1(n_1015),
.B2(n_1019),
.Y(n_5775)
);

INVx2_ASAP7_75t_L g5776 ( 
.A(n_5560),
.Y(n_5776)
);

NOR2xp33_ASAP7_75t_L g5777 ( 
.A(n_5558),
.B(n_1020),
.Y(n_5777)
);

INVx1_ASAP7_75t_L g5778 ( 
.A(n_5570),
.Y(n_5778)
);

INVx1_ASAP7_75t_L g5779 ( 
.A(n_5570),
.Y(n_5779)
);

NAND2xp5_ASAP7_75t_L g5780 ( 
.A(n_5574),
.B(n_1023),
.Y(n_5780)
);

NOR2xp33_ASAP7_75t_L g5781 ( 
.A(n_5558),
.B(n_1024),
.Y(n_5781)
);

OAI22xp33_ASAP7_75t_L g5782 ( 
.A1(n_5609),
.A2(n_1028),
.B1(n_1026),
.B2(n_1027),
.Y(n_5782)
);

AOI222xp33_ASAP7_75t_L g5783 ( 
.A1(n_5584),
.A2(n_1054),
.B1(n_1038),
.B2(n_1062),
.C1(n_1046),
.C2(n_1027),
.Y(n_5783)
);

OR2x2_ASAP7_75t_L g5784 ( 
.A(n_5589),
.B(n_1029),
.Y(n_5784)
);

AND2x2_ASAP7_75t_L g5785 ( 
.A(n_5594),
.B(n_1029),
.Y(n_5785)
);

OR2x2_ASAP7_75t_L g5786 ( 
.A(n_5759),
.B(n_1030),
.Y(n_5786)
);

INVx1_ASAP7_75t_L g5787 ( 
.A(n_5765),
.Y(n_5787)
);

NOR2xp33_ASAP7_75t_L g5788 ( 
.A(n_5737),
.B(n_1030),
.Y(n_5788)
);

NAND2xp5_ASAP7_75t_L g5789 ( 
.A(n_5753),
.B(n_1031),
.Y(n_5789)
);

OAI21xp33_ASAP7_75t_L g5790 ( 
.A1(n_5657),
.A2(n_1031),
.B(n_1032),
.Y(n_5790)
);

AND2x2_ASAP7_75t_L g5791 ( 
.A(n_5772),
.B(n_5664),
.Y(n_5791)
);

OAI21xp5_ASAP7_75t_L g5792 ( 
.A1(n_5655),
.A2(n_1038),
.B(n_1037),
.Y(n_5792)
);

HB1xp67_ASAP7_75t_L g5793 ( 
.A(n_5728),
.Y(n_5793)
);

AND2x2_ASAP7_75t_L g5794 ( 
.A(n_5756),
.B(n_1036),
.Y(n_5794)
);

AOI22xp33_ASAP7_75t_L g5795 ( 
.A1(n_5692),
.A2(n_1040),
.B1(n_1037),
.B2(n_1039),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_5661),
.Y(n_5796)
);

INVxp33_ASAP7_75t_L g5797 ( 
.A(n_5774),
.Y(n_5797)
);

AND2x2_ASAP7_75t_L g5798 ( 
.A(n_5761),
.B(n_1041),
.Y(n_5798)
);

AND2x2_ASAP7_75t_L g5799 ( 
.A(n_5776),
.B(n_1043),
.Y(n_5799)
);

AOI21xp33_ASAP7_75t_SL g5800 ( 
.A1(n_5658),
.A2(n_5659),
.B(n_5720),
.Y(n_5800)
);

OAI22xp5_ASAP7_75t_L g5801 ( 
.A1(n_5716),
.A2(n_1048),
.B1(n_1046),
.B2(n_1047),
.Y(n_5801)
);

OAI21xp5_ASAP7_75t_L g5802 ( 
.A1(n_5770),
.A2(n_5690),
.B(n_5660),
.Y(n_5802)
);

AND2x2_ASAP7_75t_L g5803 ( 
.A(n_5678),
.B(n_1048),
.Y(n_5803)
);

NOR3xp33_ASAP7_75t_L g5804 ( 
.A(n_5721),
.B(n_1049),
.C(n_1050),
.Y(n_5804)
);

NAND2xp5_ASAP7_75t_L g5805 ( 
.A(n_5732),
.B(n_1049),
.Y(n_5805)
);

OAI22xp5_ASAP7_75t_L g5806 ( 
.A1(n_5725),
.A2(n_5746),
.B1(n_5762),
.B2(n_5745),
.Y(n_5806)
);

AND2x2_ASAP7_75t_L g5807 ( 
.A(n_5672),
.B(n_1051),
.Y(n_5807)
);

AOI221xp5_ASAP7_75t_L g5808 ( 
.A1(n_5695),
.A2(n_1764),
.B1(n_1766),
.B2(n_1762),
.C(n_1761),
.Y(n_5808)
);

INVx1_ASAP7_75t_L g5809 ( 
.A(n_5734),
.Y(n_5809)
);

INVx1_ASAP7_75t_L g5810 ( 
.A(n_5751),
.Y(n_5810)
);

NOR2xp33_ASAP7_75t_L g5811 ( 
.A(n_5738),
.B(n_1051),
.Y(n_5811)
);

AOI222xp33_ASAP7_75t_L g5812 ( 
.A1(n_5730),
.A2(n_1055),
.B1(n_1057),
.B2(n_1052),
.C1(n_1053),
.C2(n_1056),
.Y(n_5812)
);

AOI22xp33_ASAP7_75t_L g5813 ( 
.A1(n_5735),
.A2(n_1055),
.B1(n_1052),
.B2(n_1053),
.Y(n_5813)
);

NAND2xp5_ASAP7_75t_L g5814 ( 
.A(n_5771),
.B(n_1056),
.Y(n_5814)
);

NAND4xp25_ASAP7_75t_L g5815 ( 
.A(n_5712),
.B(n_1059),
.C(n_1057),
.D(n_1058),
.Y(n_5815)
);

OAI22xp5_ASAP7_75t_L g5816 ( 
.A1(n_5775),
.A2(n_1063),
.B1(n_1059),
.B2(n_1061),
.Y(n_5816)
);

INVx1_ASAP7_75t_SL g5817 ( 
.A(n_5785),
.Y(n_5817)
);

AOI32xp33_ASAP7_75t_L g5818 ( 
.A1(n_5736),
.A2(n_1064),
.A3(n_1061),
.B1(n_1063),
.B2(n_1065),
.Y(n_5818)
);

OAI22xp5_ASAP7_75t_L g5819 ( 
.A1(n_5714),
.A2(n_1067),
.B1(n_1064),
.B2(n_1066),
.Y(n_5819)
);

O2A1O1Ixp33_ASAP7_75t_L g5820 ( 
.A1(n_5705),
.A2(n_1070),
.B(n_1068),
.C(n_1069),
.Y(n_5820)
);

INVx1_ASAP7_75t_SL g5821 ( 
.A(n_5656),
.Y(n_5821)
);

NAND2xp5_ASAP7_75t_L g5822 ( 
.A(n_5722),
.B(n_1071),
.Y(n_5822)
);

INVx1_ASAP7_75t_L g5823 ( 
.A(n_5727),
.Y(n_5823)
);

INVx1_ASAP7_75t_L g5824 ( 
.A(n_5744),
.Y(n_5824)
);

AND2x2_ASAP7_75t_L g5825 ( 
.A(n_5685),
.B(n_1072),
.Y(n_5825)
);

OR2x6_ASAP7_75t_L g5826 ( 
.A(n_5760),
.B(n_1073),
.Y(n_5826)
);

OAI22xp5_ASAP7_75t_L g5827 ( 
.A1(n_5758),
.A2(n_1077),
.B1(n_1074),
.B2(n_1076),
.Y(n_5827)
);

OAI22xp33_ASAP7_75t_L g5828 ( 
.A1(n_5676),
.A2(n_1077),
.B1(n_1074),
.B2(n_1076),
.Y(n_5828)
);

NAND2xp5_ASAP7_75t_L g5829 ( 
.A(n_5733),
.B(n_5739),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_5773),
.Y(n_5830)
);

INVx2_ASAP7_75t_SL g5831 ( 
.A(n_5684),
.Y(n_5831)
);

INVx1_ASAP7_75t_L g5832 ( 
.A(n_5780),
.Y(n_5832)
);

NAND2xp5_ASAP7_75t_L g5833 ( 
.A(n_5749),
.B(n_1078),
.Y(n_5833)
);

OAI21xp33_ASAP7_75t_L g5834 ( 
.A1(n_5691),
.A2(n_1079),
.B(n_1081),
.Y(n_5834)
);

INVx2_ASAP7_75t_L g5835 ( 
.A(n_5724),
.Y(n_5835)
);

NOR2xp33_ASAP7_75t_L g5836 ( 
.A(n_5731),
.B(n_1082),
.Y(n_5836)
);

CKINVDCx5p33_ASAP7_75t_R g5837 ( 
.A(n_5679),
.Y(n_5837)
);

OAI32xp33_ASAP7_75t_L g5838 ( 
.A1(n_5670),
.A2(n_1098),
.A3(n_1106),
.B1(n_1091),
.B2(n_1082),
.Y(n_5838)
);

INVxp67_ASAP7_75t_L g5839 ( 
.A(n_5740),
.Y(n_5839)
);

OAI21xp5_ASAP7_75t_L g5840 ( 
.A1(n_5680),
.A2(n_1085),
.B(n_1084),
.Y(n_5840)
);

OR2x2_ASAP7_75t_L g5841 ( 
.A(n_5750),
.B(n_1083),
.Y(n_5841)
);

OAI32xp33_ASAP7_75t_L g5842 ( 
.A1(n_5768),
.A2(n_1101),
.A3(n_1109),
.B1(n_1094),
.B2(n_1084),
.Y(n_5842)
);

AOI22xp5_ASAP7_75t_L g5843 ( 
.A1(n_5717),
.A2(n_1790),
.B1(n_1795),
.B2(n_1778),
.Y(n_5843)
);

INVx1_ASAP7_75t_L g5844 ( 
.A(n_5729),
.Y(n_5844)
);

OAI22xp33_ASAP7_75t_L g5845 ( 
.A1(n_5665),
.A2(n_1089),
.B1(n_1087),
.B2(n_1088),
.Y(n_5845)
);

NAND2xp5_ASAP7_75t_L g5846 ( 
.A(n_5754),
.B(n_1090),
.Y(n_5846)
);

OAI22xp5_ASAP7_75t_L g5847 ( 
.A1(n_5763),
.A2(n_1093),
.B1(n_1091),
.B2(n_1092),
.Y(n_5847)
);

NOR3xp33_ASAP7_75t_SL g5848 ( 
.A(n_5755),
.B(n_5767),
.C(n_5757),
.Y(n_5848)
);

INVx1_ASAP7_75t_L g5849 ( 
.A(n_5764),
.Y(n_5849)
);

INVx1_ASAP7_75t_L g5850 ( 
.A(n_5784),
.Y(n_5850)
);

NAND3xp33_ASAP7_75t_L g5851 ( 
.A(n_5778),
.B(n_1093),
.C(n_1094),
.Y(n_5851)
);

INVx1_ASAP7_75t_L g5852 ( 
.A(n_5779),
.Y(n_5852)
);

NAND3xp33_ASAP7_75t_L g5853 ( 
.A(n_5711),
.B(n_1095),
.C(n_1096),
.Y(n_5853)
);

INVx2_ASAP7_75t_L g5854 ( 
.A(n_5724),
.Y(n_5854)
);

O2A1O1Ixp33_ASAP7_75t_L g5855 ( 
.A1(n_5673),
.A2(n_1098),
.B(n_1096),
.C(n_1097),
.Y(n_5855)
);

NAND2xp5_ASAP7_75t_L g5856 ( 
.A(n_5668),
.B(n_1099),
.Y(n_5856)
);

INVx1_ASAP7_75t_L g5857 ( 
.A(n_5662),
.Y(n_5857)
);

NOR4xp25_ASAP7_75t_SL g5858 ( 
.A(n_5687),
.B(n_1102),
.C(n_1103),
.D(n_1100),
.Y(n_5858)
);

OAI31xp33_ASAP7_75t_L g5859 ( 
.A1(n_5702),
.A2(n_1102),
.A3(n_1099),
.B(n_1100),
.Y(n_5859)
);

AOI21xp33_ASAP7_75t_L g5860 ( 
.A1(n_5697),
.A2(n_1103),
.B(n_1104),
.Y(n_5860)
);

INVx2_ASAP7_75t_L g5861 ( 
.A(n_5700),
.Y(n_5861)
);

AND2x2_ASAP7_75t_L g5862 ( 
.A(n_5706),
.B(n_1105),
.Y(n_5862)
);

AOI22xp5_ASAP7_75t_L g5863 ( 
.A1(n_5675),
.A2(n_1753),
.B1(n_1755),
.B2(n_1752),
.Y(n_5863)
);

OAI221xp5_ASAP7_75t_SL g5864 ( 
.A1(n_5696),
.A2(n_1110),
.B1(n_1107),
.B2(n_1108),
.C(n_1111),
.Y(n_5864)
);

INVx2_ASAP7_75t_L g5865 ( 
.A(n_5693),
.Y(n_5865)
);

AOI222xp33_ASAP7_75t_L g5866 ( 
.A1(n_5694),
.A2(n_1112),
.B1(n_1114),
.B2(n_1107),
.C1(n_1111),
.C2(n_1113),
.Y(n_5866)
);

A2O1A1Ixp33_ASAP7_75t_L g5867 ( 
.A1(n_5663),
.A2(n_1118),
.B(n_1116),
.C(n_1117),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_5667),
.Y(n_5868)
);

INVx1_ASAP7_75t_L g5869 ( 
.A(n_5682),
.Y(n_5869)
);

AND2x2_ASAP7_75t_L g5870 ( 
.A(n_5686),
.B(n_1116),
.Y(n_5870)
);

NAND2xp5_ASAP7_75t_L g5871 ( 
.A(n_5743),
.B(n_1117),
.Y(n_5871)
);

AND2x4_ASAP7_75t_L g5872 ( 
.A(n_5671),
.B(n_1118),
.Y(n_5872)
);

AOI22xp5_ASAP7_75t_L g5873 ( 
.A1(n_5777),
.A2(n_1122),
.B1(n_1120),
.B2(n_1121),
.Y(n_5873)
);

NOR2xp33_ASAP7_75t_L g5874 ( 
.A(n_5741),
.B(n_1121),
.Y(n_5874)
);

INVx1_ASAP7_75t_L g5875 ( 
.A(n_5669),
.Y(n_5875)
);

NAND2xp5_ASAP7_75t_L g5876 ( 
.A(n_5781),
.B(n_1122),
.Y(n_5876)
);

INVx2_ASAP7_75t_SL g5877 ( 
.A(n_5710),
.Y(n_5877)
);

INVx1_ASAP7_75t_L g5878 ( 
.A(n_5674),
.Y(n_5878)
);

NAND3xp33_ASAP7_75t_SL g5879 ( 
.A(n_5723),
.B(n_1123),
.C(n_1124),
.Y(n_5879)
);

INVx1_ASAP7_75t_SL g5880 ( 
.A(n_5747),
.Y(n_5880)
);

AOI21xp5_ASAP7_75t_L g5881 ( 
.A1(n_5701),
.A2(n_1126),
.B(n_1127),
.Y(n_5881)
);

NAND2xp5_ASAP7_75t_L g5882 ( 
.A(n_5748),
.B(n_1126),
.Y(n_5882)
);

AND2x2_ASAP7_75t_L g5883 ( 
.A(n_5677),
.B(n_1127),
.Y(n_5883)
);

INVx1_ASAP7_75t_L g5884 ( 
.A(n_5683),
.Y(n_5884)
);

OAI32xp33_ASAP7_75t_L g5885 ( 
.A1(n_5708),
.A2(n_1146),
.A3(n_1156),
.B1(n_1137),
.B2(n_1129),
.Y(n_5885)
);

INVx2_ASAP7_75t_L g5886 ( 
.A(n_5704),
.Y(n_5886)
);

AOI22xp5_ASAP7_75t_L g5887 ( 
.A1(n_5709),
.A2(n_1771),
.B1(n_1775),
.B2(n_1769),
.Y(n_5887)
);

AND2x2_ASAP7_75t_L g5888 ( 
.A(n_5689),
.B(n_1130),
.Y(n_5888)
);

AOI322xp5_ASAP7_75t_L g5889 ( 
.A1(n_5752),
.A2(n_5782),
.A3(n_5713),
.B1(n_5707),
.B2(n_5718),
.C1(n_5699),
.C2(n_5698),
.Y(n_5889)
);

INVx1_ASAP7_75t_L g5890 ( 
.A(n_5719),
.Y(n_5890)
);

INVx1_ASAP7_75t_SL g5891 ( 
.A(n_5715),
.Y(n_5891)
);

NAND2xp5_ASAP7_75t_SL g5892 ( 
.A(n_5837),
.B(n_5688),
.Y(n_5892)
);

AOI211xp5_ASAP7_75t_L g5893 ( 
.A1(n_5800),
.A2(n_5766),
.B(n_5666),
.C(n_5703),
.Y(n_5893)
);

AOI22xp5_ASAP7_75t_L g5894 ( 
.A1(n_5804),
.A2(n_5769),
.B1(n_5783),
.B2(n_5742),
.Y(n_5894)
);

NAND3xp33_ASAP7_75t_L g5895 ( 
.A(n_5848),
.B(n_5726),
.C(n_5681),
.Y(n_5895)
);

AOI21xp5_ASAP7_75t_L g5896 ( 
.A1(n_5802),
.A2(n_1130),
.B(n_1131),
.Y(n_5896)
);

OAI21xp5_ASAP7_75t_L g5897 ( 
.A1(n_5793),
.A2(n_1132),
.B(n_1133),
.Y(n_5897)
);

NAND4xp25_ASAP7_75t_L g5898 ( 
.A(n_5791),
.B(n_1138),
.C(n_1134),
.D(n_1136),
.Y(n_5898)
);

OAI222xp33_ASAP7_75t_L g5899 ( 
.A1(n_5880),
.A2(n_1757),
.B1(n_1755),
.B2(n_1758),
.C1(n_1756),
.C2(n_1751),
.Y(n_5899)
);

AOI22xp5_ASAP7_75t_L g5900 ( 
.A1(n_5796),
.A2(n_1144),
.B1(n_1141),
.B2(n_1142),
.Y(n_5900)
);

O2A1O1Ixp5_ASAP7_75t_SL g5901 ( 
.A1(n_5787),
.A2(n_1145),
.B(n_1142),
.C(n_1144),
.Y(n_5901)
);

OAI22xp5_ASAP7_75t_L g5902 ( 
.A1(n_5817),
.A2(n_1151),
.B1(n_1147),
.B2(n_1149),
.Y(n_5902)
);

O2A1O1Ixp33_ASAP7_75t_SL g5903 ( 
.A1(n_5867),
.A2(n_1153),
.B(n_1149),
.C(n_1151),
.Y(n_5903)
);

AO22x1_ASAP7_75t_L g5904 ( 
.A1(n_5835),
.A2(n_1159),
.B1(n_1157),
.B2(n_1158),
.Y(n_5904)
);

AOI322xp5_ASAP7_75t_L g5905 ( 
.A1(n_5879),
.A2(n_1747),
.A3(n_1163),
.B1(n_1160),
.B2(n_1162),
.C1(n_1157),
.C2(n_1158),
.Y(n_5905)
);

INVx1_ASAP7_75t_L g5906 ( 
.A(n_5854),
.Y(n_5906)
);

OAI211xp5_ASAP7_75t_SL g5907 ( 
.A1(n_5889),
.A2(n_1163),
.B(n_1160),
.C(n_1161),
.Y(n_5907)
);

AOI222xp33_ASAP7_75t_L g5908 ( 
.A1(n_5806),
.A2(n_1166),
.B1(n_1168),
.B2(n_1164),
.C1(n_1165),
.C2(n_1167),
.Y(n_5908)
);

AOI22xp5_ASAP7_75t_L g5909 ( 
.A1(n_5801),
.A2(n_1171),
.B1(n_1169),
.B2(n_1170),
.Y(n_5909)
);

NAND3x1_ASAP7_75t_L g5910 ( 
.A(n_5789),
.B(n_1169),
.C(n_1170),
.Y(n_5910)
);

AOI21xp5_ASAP7_75t_L g5911 ( 
.A1(n_5881),
.A2(n_1171),
.B(n_1172),
.Y(n_5911)
);

AOI211xp5_ASAP7_75t_L g5912 ( 
.A1(n_5815),
.A2(n_1747),
.B(n_1748),
.C(n_1746),
.Y(n_5912)
);

A2O1A1Ixp33_ASAP7_75t_L g5913 ( 
.A1(n_5820),
.A2(n_1182),
.B(n_1189),
.C(n_1173),
.Y(n_5913)
);

AOI221xp5_ASAP7_75t_L g5914 ( 
.A1(n_5855),
.A2(n_1176),
.B1(n_1174),
.B2(n_1175),
.C(n_1177),
.Y(n_5914)
);

NAND3xp33_ASAP7_75t_SL g5915 ( 
.A(n_5858),
.B(n_1180),
.C(n_1179),
.Y(n_5915)
);

NOR2xp33_ASAP7_75t_L g5916 ( 
.A(n_5821),
.B(n_1178),
.Y(n_5916)
);

AOI211xp5_ASAP7_75t_L g5917 ( 
.A1(n_5842),
.A2(n_1741),
.B(n_1742),
.C(n_1740),
.Y(n_5917)
);

AOI222xp33_ASAP7_75t_L g5918 ( 
.A1(n_5829),
.A2(n_1184),
.B1(n_1186),
.B2(n_1182),
.C1(n_1183),
.C2(n_1185),
.Y(n_5918)
);

INVx1_ASAP7_75t_L g5919 ( 
.A(n_5803),
.Y(n_5919)
);

NOR3xp33_ASAP7_75t_L g5920 ( 
.A(n_5839),
.B(n_1188),
.C(n_1190),
.Y(n_5920)
);

AOI22xp5_ASAP7_75t_L g5921 ( 
.A1(n_5809),
.A2(n_1193),
.B1(n_1190),
.B2(n_1191),
.Y(n_5921)
);

OAI22xp5_ASAP7_75t_L g5922 ( 
.A1(n_5810),
.A2(n_1196),
.B1(n_1194),
.B2(n_1195),
.Y(n_5922)
);

AOI221xp5_ASAP7_75t_SL g5923 ( 
.A1(n_5852),
.A2(n_1198),
.B1(n_1194),
.B2(n_1196),
.C(n_1199),
.Y(n_5923)
);

INVx1_ASAP7_75t_L g5924 ( 
.A(n_5786),
.Y(n_5924)
);

OAI22xp5_ASAP7_75t_L g5925 ( 
.A1(n_5864),
.A2(n_1201),
.B1(n_1199),
.B2(n_1200),
.Y(n_5925)
);

OAI211xp5_ASAP7_75t_L g5926 ( 
.A1(n_5808),
.A2(n_1206),
.B(n_1202),
.C(n_1203),
.Y(n_5926)
);

AOI211xp5_ASAP7_75t_SL g5927 ( 
.A1(n_5890),
.A2(n_1208),
.B(n_1206),
.C(n_1207),
.Y(n_5927)
);

A2O1A1Ixp33_ASAP7_75t_L g5928 ( 
.A1(n_5818),
.A2(n_1215),
.B(n_1223),
.C(n_1207),
.Y(n_5928)
);

OAI211xp5_ASAP7_75t_SL g5929 ( 
.A1(n_5891),
.A2(n_1210),
.B(n_1208),
.C(n_1209),
.Y(n_5929)
);

OR2x2_ASAP7_75t_L g5930 ( 
.A(n_5861),
.B(n_1210),
.Y(n_5930)
);

AOI221xp5_ASAP7_75t_L g5931 ( 
.A1(n_5838),
.A2(n_1213),
.B1(n_1211),
.B2(n_1212),
.C(n_1214),
.Y(n_5931)
);

OAI211xp5_ASAP7_75t_SL g5932 ( 
.A1(n_5844),
.A2(n_1215),
.B(n_1213),
.C(n_1214),
.Y(n_5932)
);

NOR3xp33_ASAP7_75t_L g5933 ( 
.A(n_5849),
.B(n_1216),
.C(n_1217),
.Y(n_5933)
);

A2O1A1Ixp33_ASAP7_75t_L g5934 ( 
.A1(n_5853),
.A2(n_5811),
.B(n_5859),
.C(n_5834),
.Y(n_5934)
);

AOI22xp33_ASAP7_75t_L g5935 ( 
.A1(n_5865),
.A2(n_1221),
.B1(n_1219),
.B2(n_1220),
.Y(n_5935)
);

NAND3xp33_ASAP7_75t_SL g5936 ( 
.A(n_5812),
.B(n_1222),
.C(n_1221),
.Y(n_5936)
);

NOR2xp33_ASAP7_75t_L g5937 ( 
.A(n_5790),
.B(n_1219),
.Y(n_5937)
);

AO21x1_ASAP7_75t_L g5938 ( 
.A1(n_5836),
.A2(n_1745),
.B(n_1222),
.Y(n_5938)
);

AOI22xp5_ASAP7_75t_L g5939 ( 
.A1(n_5788),
.A2(n_1226),
.B1(n_1223),
.B2(n_1224),
.Y(n_5939)
);

AOI22xp33_ASAP7_75t_L g5940 ( 
.A1(n_5886),
.A2(n_1227),
.B1(n_1224),
.B2(n_1226),
.Y(n_5940)
);

INVx1_ASAP7_75t_L g5941 ( 
.A(n_5825),
.Y(n_5941)
);

INVx1_ASAP7_75t_L g5942 ( 
.A(n_5807),
.Y(n_5942)
);

OAI211xp5_ASAP7_75t_L g5943 ( 
.A1(n_5866),
.A2(n_1230),
.B(n_1227),
.C(n_1229),
.Y(n_5943)
);

OAI221xp5_ASAP7_75t_L g5944 ( 
.A1(n_5792),
.A2(n_1231),
.B1(n_1229),
.B2(n_1230),
.C(n_1232),
.Y(n_5944)
);

OAI211xp5_ASAP7_75t_L g5945 ( 
.A1(n_5840),
.A2(n_1233),
.B(n_1231),
.C(n_1232),
.Y(n_5945)
);

AOI22xp33_ASAP7_75t_SL g5946 ( 
.A1(n_5877),
.A2(n_1236),
.B1(n_1234),
.B2(n_1235),
.Y(n_5946)
);

INVx1_ASAP7_75t_L g5947 ( 
.A(n_5794),
.Y(n_5947)
);

NOR3xp33_ASAP7_75t_SL g5948 ( 
.A(n_5850),
.B(n_1236),
.C(n_1237),
.Y(n_5948)
);

OAI221xp5_ASAP7_75t_L g5949 ( 
.A1(n_5805),
.A2(n_1241),
.B1(n_1239),
.B2(n_1240),
.C(n_1242),
.Y(n_5949)
);

INVx1_ASAP7_75t_L g5950 ( 
.A(n_5798),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5799),
.Y(n_5951)
);

NAND2xp5_ASAP7_75t_SL g5952 ( 
.A(n_5828),
.B(n_1243),
.Y(n_5952)
);

OAI221xp5_ASAP7_75t_L g5953 ( 
.A1(n_5882),
.A2(n_1247),
.B1(n_1245),
.B2(n_1246),
.C(n_1248),
.Y(n_5953)
);

AOI322xp5_ASAP7_75t_L g5954 ( 
.A1(n_5888),
.A2(n_1749),
.A3(n_1738),
.B1(n_1253),
.B2(n_1250),
.C1(n_1252),
.C2(n_1248),
.Y(n_5954)
);

OAI22xp5_ASAP7_75t_L g5955 ( 
.A1(n_5863),
.A2(n_5813),
.B1(n_5851),
.B2(n_5795),
.Y(n_5955)
);

AOI21xp5_ASAP7_75t_L g5956 ( 
.A1(n_5814),
.A2(n_1249),
.B(n_1250),
.Y(n_5956)
);

AOI211xp5_ASAP7_75t_SL g5957 ( 
.A1(n_5823),
.A2(n_1255),
.B(n_1251),
.C(n_1254),
.Y(n_5957)
);

OAI21xp5_ASAP7_75t_SL g5958 ( 
.A1(n_5824),
.A2(n_1254),
.B(n_1255),
.Y(n_5958)
);

AOI21xp33_ASAP7_75t_L g5959 ( 
.A1(n_5830),
.A2(n_1257),
.B(n_1258),
.Y(n_5959)
);

OA21x2_ASAP7_75t_L g5960 ( 
.A1(n_5822),
.A2(n_1259),
.B(n_1261),
.Y(n_5960)
);

AOI22xp5_ASAP7_75t_L g5961 ( 
.A1(n_5832),
.A2(n_1263),
.B1(n_1261),
.B2(n_1262),
.Y(n_5961)
);

AOI21xp5_ASAP7_75t_L g5962 ( 
.A1(n_5819),
.A2(n_1264),
.B(n_1265),
.Y(n_5962)
);

OAI221xp5_ASAP7_75t_SL g5963 ( 
.A1(n_5875),
.A2(n_1739),
.B1(n_1741),
.B2(n_1738),
.C(n_1737),
.Y(n_5963)
);

OAI211xp5_ASAP7_75t_L g5964 ( 
.A1(n_5878),
.A2(n_1267),
.B(n_1265),
.C(n_1266),
.Y(n_5964)
);

OAI221xp5_ASAP7_75t_L g5965 ( 
.A1(n_5833),
.A2(n_1268),
.B1(n_1266),
.B2(n_1267),
.C(n_1269),
.Y(n_5965)
);

AOI211xp5_ASAP7_75t_L g5966 ( 
.A1(n_5845),
.A2(n_1746),
.B(n_1749),
.C(n_1745),
.Y(n_5966)
);

OAI221xp5_ASAP7_75t_L g5967 ( 
.A1(n_5846),
.A2(n_5884),
.B1(n_5869),
.B2(n_5868),
.C(n_5857),
.Y(n_5967)
);

NOR4xp25_ASAP7_75t_SL g5968 ( 
.A(n_5860),
.B(n_1274),
.C(n_1272),
.D(n_1273),
.Y(n_5968)
);

OAI21xp5_ASAP7_75t_SL g5969 ( 
.A1(n_5862),
.A2(n_1274),
.B(n_1275),
.Y(n_5969)
);

NAND2xp5_ASAP7_75t_L g5970 ( 
.A(n_5883),
.B(n_1276),
.Y(n_5970)
);

NOR2x1_ASAP7_75t_L g5971 ( 
.A(n_5826),
.B(n_1278),
.Y(n_5971)
);

OAI221xp5_ASAP7_75t_L g5972 ( 
.A1(n_5816),
.A2(n_1281),
.B1(n_1279),
.B2(n_1280),
.C(n_1282),
.Y(n_5972)
);

NAND2xp5_ASAP7_75t_L g5973 ( 
.A(n_5870),
.B(n_1280),
.Y(n_5973)
);

OAI221xp5_ASAP7_75t_L g5974 ( 
.A1(n_5887),
.A2(n_1285),
.B1(n_1282),
.B2(n_1283),
.C(n_1287),
.Y(n_5974)
);

AOI22xp33_ASAP7_75t_L g5975 ( 
.A1(n_5827),
.A2(n_1287),
.B1(n_1283),
.B2(n_1285),
.Y(n_5975)
);

AOI21xp5_ASAP7_75t_L g5976 ( 
.A1(n_5871),
.A2(n_1288),
.B(n_1289),
.Y(n_5976)
);

AOI211xp5_ASAP7_75t_L g5977 ( 
.A1(n_5885),
.A2(n_1760),
.B(n_1759),
.C(n_1291),
.Y(n_5977)
);

NOR3xp33_ASAP7_75t_L g5978 ( 
.A(n_5847),
.B(n_1288),
.C(n_1290),
.Y(n_5978)
);

AO21x1_ASAP7_75t_L g5979 ( 
.A1(n_5874),
.A2(n_1760),
.B(n_1291),
.Y(n_5979)
);

OAI22xp5_ASAP7_75t_L g5980 ( 
.A1(n_5856),
.A2(n_1294),
.B1(n_1292),
.B2(n_1293),
.Y(n_5980)
);

AOI21xp5_ASAP7_75t_L g5981 ( 
.A1(n_5876),
.A2(n_1292),
.B(n_1294),
.Y(n_5981)
);

AOI211xp5_ASAP7_75t_L g5982 ( 
.A1(n_5841),
.A2(n_1734),
.B(n_1735),
.C(n_1733),
.Y(n_5982)
);

NAND2xp5_ASAP7_75t_L g5983 ( 
.A(n_5872),
.B(n_1295),
.Y(n_5983)
);

NAND3xp33_ASAP7_75t_L g5984 ( 
.A(n_5873),
.B(n_1297),
.C(n_1298),
.Y(n_5984)
);

O2A1O1Ixp5_ASAP7_75t_L g5985 ( 
.A1(n_5797),
.A2(n_1299),
.B(n_1297),
.C(n_1298),
.Y(n_5985)
);

AOI221xp5_ASAP7_75t_L g5986 ( 
.A1(n_5848),
.A2(n_1302),
.B1(n_1300),
.B2(n_1301),
.C(n_1303),
.Y(n_5986)
);

O2A1O1Ixp5_ASAP7_75t_SL g5987 ( 
.A1(n_5787),
.A2(n_1304),
.B(n_1301),
.C(n_1302),
.Y(n_5987)
);

INVx1_ASAP7_75t_L g5988 ( 
.A(n_5831),
.Y(n_5988)
);

NAND4xp25_ASAP7_75t_SL g5989 ( 
.A(n_5843),
.B(n_1308),
.C(n_1306),
.D(n_1307),
.Y(n_5989)
);

INVx2_ASAP7_75t_L g5990 ( 
.A(n_5831),
.Y(n_5990)
);

AOI211x1_ASAP7_75t_L g5991 ( 
.A1(n_5802),
.A2(n_1312),
.B(n_1310),
.C(n_1311),
.Y(n_5991)
);

NAND2xp5_ASAP7_75t_L g5992 ( 
.A(n_5831),
.B(n_1312),
.Y(n_5992)
);

NOR3xp33_ASAP7_75t_L g5993 ( 
.A(n_5800),
.B(n_1313),
.C(n_1314),
.Y(n_5993)
);

O2A1O1Ixp33_ASAP7_75t_L g5994 ( 
.A1(n_5867),
.A2(n_1317),
.B(n_1315),
.C(n_1316),
.Y(n_5994)
);

INVx1_ASAP7_75t_L g5995 ( 
.A(n_5831),
.Y(n_5995)
);

AOI21xp5_ASAP7_75t_L g5996 ( 
.A1(n_5802),
.A2(n_1317),
.B(n_1318),
.Y(n_5996)
);

OAI211xp5_ASAP7_75t_L g5997 ( 
.A1(n_5843),
.A2(n_1321),
.B(n_1319),
.C(n_1320),
.Y(n_5997)
);

OAI21xp5_ASAP7_75t_L g5998 ( 
.A1(n_5848),
.A2(n_1322),
.B(n_1325),
.Y(n_5998)
);

OAI222xp33_ASAP7_75t_L g5999 ( 
.A1(n_5843),
.A2(n_1734),
.B1(n_1732),
.B2(n_1736),
.C1(n_1733),
.C2(n_1731),
.Y(n_5999)
);

O2A1O1Ixp5_ASAP7_75t_L g6000 ( 
.A1(n_5797),
.A2(n_1330),
.B(n_1326),
.C(n_1327),
.Y(n_6000)
);

NOR2xp67_ASAP7_75t_L g6001 ( 
.A(n_5831),
.B(n_1333),
.Y(n_6001)
);

NAND2xp5_ASAP7_75t_L g6002 ( 
.A(n_5831),
.B(n_1333),
.Y(n_6002)
);

OR2x2_ASAP7_75t_L g6003 ( 
.A(n_5831),
.B(n_1334),
.Y(n_6003)
);

NAND2xp5_ASAP7_75t_L g6004 ( 
.A(n_5831),
.B(n_1335),
.Y(n_6004)
);

NAND2xp5_ASAP7_75t_L g6005 ( 
.A(n_6001),
.B(n_1338),
.Y(n_6005)
);

INVx3_ASAP7_75t_L g6006 ( 
.A(n_5990),
.Y(n_6006)
);

AOI221xp5_ASAP7_75t_L g6007 ( 
.A1(n_5907),
.A2(n_1341),
.B1(n_1344),
.B2(n_1340),
.C(n_1343),
.Y(n_6007)
);

AOI221xp5_ASAP7_75t_L g6008 ( 
.A1(n_5895),
.A2(n_1343),
.B1(n_1345),
.B2(n_1341),
.C(n_1344),
.Y(n_6008)
);

OAI21xp5_ASAP7_75t_SL g6009 ( 
.A1(n_5894),
.A2(n_1339),
.B(n_1347),
.Y(n_6009)
);

INVx1_ASAP7_75t_L g6010 ( 
.A(n_5971),
.Y(n_6010)
);

O2A1O1Ixp33_ASAP7_75t_L g6011 ( 
.A1(n_5915),
.A2(n_1355),
.B(n_1365),
.C(n_1339),
.Y(n_6011)
);

AOI21xp5_ASAP7_75t_L g6012 ( 
.A1(n_5892),
.A2(n_1348),
.B(n_1349),
.Y(n_6012)
);

INVx1_ASAP7_75t_L g6013 ( 
.A(n_6003),
.Y(n_6013)
);

AOI22xp33_ASAP7_75t_L g6014 ( 
.A1(n_5993),
.A2(n_1352),
.B1(n_1350),
.B2(n_1351),
.Y(n_6014)
);

NOR3xp33_ASAP7_75t_L g6015 ( 
.A(n_5967),
.B(n_1364),
.C(n_1354),
.Y(n_6015)
);

OAI322xp33_ASAP7_75t_L g6016 ( 
.A1(n_5988),
.A2(n_1361),
.A3(n_1359),
.B1(n_1357),
.B2(n_1355),
.C1(n_1356),
.C2(n_1358),
.Y(n_6016)
);

INVx1_ASAP7_75t_L g6017 ( 
.A(n_5995),
.Y(n_6017)
);

AOI21xp5_ASAP7_75t_L g6018 ( 
.A1(n_5998),
.A2(n_1363),
.B(n_1365),
.Y(n_6018)
);

OAI22xp5_ASAP7_75t_L g6019 ( 
.A1(n_5975),
.A2(n_1368),
.B1(n_1366),
.B2(n_1367),
.Y(n_6019)
);

OAI21xp5_ASAP7_75t_L g6020 ( 
.A1(n_5985),
.A2(n_1368),
.B(n_1369),
.Y(n_6020)
);

INVx2_ASAP7_75t_L g6021 ( 
.A(n_5906),
.Y(n_6021)
);

INVx1_ASAP7_75t_SL g6022 ( 
.A(n_5910),
.Y(n_6022)
);

NOR2x1_ASAP7_75t_L g6023 ( 
.A(n_5898),
.B(n_1370),
.Y(n_6023)
);

NAND2xp5_ASAP7_75t_L g6024 ( 
.A(n_5904),
.B(n_5927),
.Y(n_6024)
);

INVx1_ASAP7_75t_L g6025 ( 
.A(n_5992),
.Y(n_6025)
);

AOI22xp5_ASAP7_75t_L g6026 ( 
.A1(n_5989),
.A2(n_1372),
.B1(n_1370),
.B2(n_1371),
.Y(n_6026)
);

AND2x2_ASAP7_75t_L g6027 ( 
.A(n_5919),
.B(n_1373),
.Y(n_6027)
);

AND2x2_ASAP7_75t_L g6028 ( 
.A(n_5948),
.B(n_1374),
.Y(n_6028)
);

OAI22xp5_ASAP7_75t_L g6029 ( 
.A1(n_5893),
.A2(n_1377),
.B1(n_1375),
.B2(n_1376),
.Y(n_6029)
);

OAI22xp5_ASAP7_75t_L g6030 ( 
.A1(n_5909),
.A2(n_1377),
.B1(n_1375),
.B2(n_1376),
.Y(n_6030)
);

NAND2xp5_ASAP7_75t_L g6031 ( 
.A(n_5957),
.B(n_1378),
.Y(n_6031)
);

HB1xp67_ASAP7_75t_L g6032 ( 
.A(n_5960),
.Y(n_6032)
);

NOR2xp33_ASAP7_75t_L g6033 ( 
.A(n_5938),
.B(n_1379),
.Y(n_6033)
);

OAI221xp5_ASAP7_75t_SL g6034 ( 
.A1(n_5934),
.A2(n_1382),
.B1(n_1379),
.B2(n_1380),
.C(n_1383),
.Y(n_6034)
);

AOI32xp33_ASAP7_75t_L g6035 ( 
.A1(n_5929),
.A2(n_1384),
.A3(n_1382),
.B1(n_1383),
.B2(n_1385),
.Y(n_6035)
);

HB1xp67_ASAP7_75t_L g6036 ( 
.A(n_5960),
.Y(n_6036)
);

AOI22xp33_ASAP7_75t_L g6037 ( 
.A1(n_5936),
.A2(n_1390),
.B1(n_1388),
.B2(n_1389),
.Y(n_6037)
);

AOI322xp5_ASAP7_75t_L g6038 ( 
.A1(n_5986),
.A2(n_1395),
.A3(n_1394),
.B1(n_1392),
.B2(n_1388),
.C1(n_1391),
.C2(n_1393),
.Y(n_6038)
);

O2A1O1Ixp33_ASAP7_75t_L g6039 ( 
.A1(n_5899),
.A2(n_5903),
.B(n_5999),
.C(n_6000),
.Y(n_6039)
);

AOI22xp5_ASAP7_75t_L g6040 ( 
.A1(n_5955),
.A2(n_1398),
.B1(n_1396),
.B2(n_1397),
.Y(n_6040)
);

AOI22xp5_ASAP7_75t_L g6041 ( 
.A1(n_5942),
.A2(n_1399),
.B1(n_1397),
.B2(n_1398),
.Y(n_6041)
);

NOR3x1_ASAP7_75t_L g6042 ( 
.A(n_5943),
.B(n_1400),
.C(n_1401),
.Y(n_6042)
);

OR2x2_ASAP7_75t_L g6043 ( 
.A(n_6002),
.B(n_1400),
.Y(n_6043)
);

OAI22xp5_ASAP7_75t_L g6044 ( 
.A1(n_5928),
.A2(n_1404),
.B1(n_1401),
.B2(n_1403),
.Y(n_6044)
);

NAND2xp5_ASAP7_75t_L g6045 ( 
.A(n_5946),
.B(n_1403),
.Y(n_6045)
);

AOI22x1_ASAP7_75t_L g6046 ( 
.A1(n_5924),
.A2(n_1406),
.B1(n_1404),
.B2(n_1405),
.Y(n_6046)
);

INVx2_ASAP7_75t_L g6047 ( 
.A(n_5930),
.Y(n_6047)
);

AND2x2_ASAP7_75t_L g6048 ( 
.A(n_5947),
.B(n_1407),
.Y(n_6048)
);

OAI31xp33_ASAP7_75t_L g6049 ( 
.A1(n_5932),
.A2(n_5926),
.A3(n_5997),
.B(n_5945),
.Y(n_6049)
);

INVx1_ASAP7_75t_L g6050 ( 
.A(n_6004),
.Y(n_6050)
);

NAND2xp5_ASAP7_75t_SL g6051 ( 
.A(n_5979),
.B(n_1408),
.Y(n_6051)
);

AND2x2_ASAP7_75t_L g6052 ( 
.A(n_5950),
.B(n_5951),
.Y(n_6052)
);

INVx1_ASAP7_75t_L g6053 ( 
.A(n_5983),
.Y(n_6053)
);

INVxp67_ASAP7_75t_L g6054 ( 
.A(n_5916),
.Y(n_6054)
);

OAI221xp5_ASAP7_75t_L g6055 ( 
.A1(n_5914),
.A2(n_5913),
.B1(n_5917),
.B2(n_5994),
.C(n_5953),
.Y(n_6055)
);

AOI21xp5_ASAP7_75t_L g6056 ( 
.A1(n_5911),
.A2(n_1409),
.B(n_1410),
.Y(n_6056)
);

INVx1_ASAP7_75t_L g6057 ( 
.A(n_5970),
.Y(n_6057)
);

AOI221xp5_ASAP7_75t_L g6058 ( 
.A1(n_5925),
.A2(n_1414),
.B1(n_1416),
.B2(n_1413),
.C(n_1415),
.Y(n_6058)
);

AOI21xp5_ASAP7_75t_L g6059 ( 
.A1(n_5952),
.A2(n_1411),
.B(n_1413),
.Y(n_6059)
);

NAND2xp5_ASAP7_75t_SL g6060 ( 
.A(n_5977),
.B(n_1417),
.Y(n_6060)
);

O2A1O1Ixp5_ASAP7_75t_L g6061 ( 
.A1(n_5941),
.A2(n_1419),
.B(n_1417),
.C(n_1418),
.Y(n_6061)
);

AOI322xp5_ASAP7_75t_L g6062 ( 
.A1(n_5923),
.A2(n_1424),
.A3(n_1423),
.B1(n_1421),
.B2(n_1418),
.C1(n_1420),
.C2(n_1422),
.Y(n_6062)
);

AOI22xp5_ASAP7_75t_L g6063 ( 
.A1(n_5978),
.A2(n_1428),
.B1(n_1426),
.B2(n_1427),
.Y(n_6063)
);

INVx2_ASAP7_75t_L g6064 ( 
.A(n_5973),
.Y(n_6064)
);

AOI221xp5_ASAP7_75t_L g6065 ( 
.A1(n_5991),
.A2(n_1430),
.B1(n_1432),
.B2(n_1429),
.C(n_1431),
.Y(n_6065)
);

AND2x2_ASAP7_75t_L g6066 ( 
.A(n_5897),
.B(n_1427),
.Y(n_6066)
);

INVxp33_ASAP7_75t_L g6067 ( 
.A(n_5937),
.Y(n_6067)
);

OAI221xp5_ASAP7_75t_SL g6068 ( 
.A1(n_6049),
.A2(n_5905),
.B1(n_5958),
.B2(n_5931),
.C(n_5969),
.Y(n_6068)
);

AO22x2_ASAP7_75t_L g6069 ( 
.A1(n_6029),
.A2(n_5996),
.B1(n_5896),
.B2(n_5981),
.Y(n_6069)
);

OAI22xp5_ASAP7_75t_L g6070 ( 
.A1(n_6037),
.A2(n_5912),
.B1(n_5984),
.B2(n_5944),
.Y(n_6070)
);

OAI22xp5_ASAP7_75t_L g6071 ( 
.A1(n_6026),
.A2(n_5966),
.B1(n_5968),
.B2(n_5982),
.Y(n_6071)
);

AOI21xp5_ASAP7_75t_L g6072 ( 
.A1(n_6011),
.A2(n_5976),
.B(n_5956),
.Y(n_6072)
);

AOI22xp33_ASAP7_75t_L g6073 ( 
.A1(n_6006),
.A2(n_5933),
.B1(n_5920),
.B2(n_5908),
.Y(n_6073)
);

AND2x2_ASAP7_75t_L g6074 ( 
.A(n_6028),
.B(n_6052),
.Y(n_6074)
);

A2O1A1Ixp33_ASAP7_75t_L g6075 ( 
.A1(n_6035),
.A2(n_6039),
.B(n_6033),
.C(n_6061),
.Y(n_6075)
);

O2A1O1Ixp5_ASAP7_75t_L g6076 ( 
.A1(n_6051),
.A2(n_5964),
.B(n_5962),
.C(n_5963),
.Y(n_6076)
);

CKINVDCx5p33_ASAP7_75t_R g6077 ( 
.A(n_6022),
.Y(n_6077)
);

INVxp67_ASAP7_75t_L g6078 ( 
.A(n_6032),
.Y(n_6078)
);

OAI22xp5_ASAP7_75t_L g6079 ( 
.A1(n_6040),
.A2(n_5974),
.B1(n_5965),
.B2(n_5949),
.Y(n_6079)
);

NOR2x1_ASAP7_75t_L g6080 ( 
.A(n_6010),
.B(n_5902),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_6036),
.Y(n_6081)
);

OAI22xp5_ASAP7_75t_L g6082 ( 
.A1(n_6014),
.A2(n_5935),
.B1(n_5940),
.B2(n_5900),
.Y(n_6082)
);

AOI221x1_ASAP7_75t_L g6083 ( 
.A1(n_6015),
.A2(n_5959),
.B1(n_5980),
.B2(n_5922),
.C(n_5918),
.Y(n_6083)
);

NAND2xp5_ASAP7_75t_L g6084 ( 
.A(n_6062),
.B(n_5954),
.Y(n_6084)
);

AND2x2_ASAP7_75t_L g6085 ( 
.A(n_6023),
.B(n_5939),
.Y(n_6085)
);

NOR2x1_ASAP7_75t_L g6086 ( 
.A(n_6016),
.B(n_5972),
.Y(n_6086)
);

NOR2xp33_ASAP7_75t_R g6087 ( 
.A(n_6013),
.B(n_1433),
.Y(n_6087)
);

AOI22xp33_ASAP7_75t_L g6088 ( 
.A1(n_6017),
.A2(n_5921),
.B1(n_5961),
.B2(n_5901),
.Y(n_6088)
);

OAI221xp5_ASAP7_75t_L g6089 ( 
.A1(n_6009),
.A2(n_5987),
.B1(n_1437),
.B2(n_1435),
.C(n_1436),
.Y(n_6089)
);

INVx2_ASAP7_75t_L g6090 ( 
.A(n_6046),
.Y(n_6090)
);

INVx1_ASAP7_75t_L g6091 ( 
.A(n_6005),
.Y(n_6091)
);

INVx1_ASAP7_75t_L g6092 ( 
.A(n_6024),
.Y(n_6092)
);

OAI22xp33_ASAP7_75t_L g6093 ( 
.A1(n_6031),
.A2(n_1439),
.B1(n_1440),
.B2(n_1438),
.Y(n_6093)
);

INVx1_ASAP7_75t_L g6094 ( 
.A(n_6027),
.Y(n_6094)
);

AOI22xp5_ASAP7_75t_L g6095 ( 
.A1(n_6060),
.A2(n_1443),
.B1(n_1441),
.B2(n_1442),
.Y(n_6095)
);

A2O1A1Ixp33_ASAP7_75t_L g6096 ( 
.A1(n_6007),
.A2(n_1446),
.B(n_1444),
.C(n_1445),
.Y(n_6096)
);

OA21x2_ASAP7_75t_SL g6097 ( 
.A1(n_6067),
.A2(n_1446),
.B(n_1447),
.Y(n_6097)
);

AOI22xp5_ASAP7_75t_L g6098 ( 
.A1(n_6054),
.A2(n_1742),
.B1(n_1743),
.B2(n_1739),
.Y(n_6098)
);

AOI211xp5_ASAP7_75t_L g6099 ( 
.A1(n_6055),
.A2(n_6020),
.B(n_6034),
.C(n_6044),
.Y(n_6099)
);

OAI21xp5_ASAP7_75t_L g6100 ( 
.A1(n_6012),
.A2(n_6018),
.B(n_6059),
.Y(n_6100)
);

NAND2xp5_ASAP7_75t_L g6101 ( 
.A(n_6048),
.B(n_6038),
.Y(n_6101)
);

NAND2xp5_ASAP7_75t_L g6102 ( 
.A(n_6065),
.B(n_1451),
.Y(n_6102)
);

AOI322xp5_ASAP7_75t_L g6103 ( 
.A1(n_6008),
.A2(n_1459),
.A3(n_1458),
.B1(n_1455),
.B2(n_1453),
.C1(n_1454),
.C2(n_1457),
.Y(n_6103)
);

NOR2x1_ASAP7_75t_L g6104 ( 
.A(n_6045),
.B(n_1453),
.Y(n_6104)
);

NAND5xp2_ASAP7_75t_L g6105 ( 
.A(n_6057),
.B(n_1474),
.C(n_1485),
.D(n_1463),
.E(n_1454),
.Y(n_6105)
);

OAI21xp5_ASAP7_75t_L g6106 ( 
.A1(n_6056),
.A2(n_6021),
.B(n_6066),
.Y(n_6106)
);

AND2x2_ASAP7_75t_L g6107 ( 
.A(n_6042),
.B(n_6047),
.Y(n_6107)
);

NOR2xp33_ASAP7_75t_R g6108 ( 
.A(n_6025),
.B(n_1455),
.Y(n_6108)
);

AOI222xp33_ASAP7_75t_L g6109 ( 
.A1(n_6050),
.A2(n_1459),
.B1(n_1461),
.B2(n_1457),
.C1(n_1458),
.C2(n_1460),
.Y(n_6109)
);

AOI22xp5_ASAP7_75t_L g6110 ( 
.A1(n_6077),
.A2(n_6058),
.B1(n_6064),
.B2(n_6053),
.Y(n_6110)
);

O2A1O1Ixp33_ASAP7_75t_SL g6111 ( 
.A1(n_6078),
.A2(n_6043),
.B(n_6030),
.C(n_6019),
.Y(n_6111)
);

AOI31xp33_ASAP7_75t_L g6112 ( 
.A1(n_6080),
.A2(n_6063),
.A3(n_6041),
.B(n_1471),
.Y(n_6112)
);

AO22x2_ASAP7_75t_L g6113 ( 
.A1(n_6081),
.A2(n_1758),
.B1(n_1756),
.B2(n_1462),
.Y(n_6113)
);

NAND2xp5_ASAP7_75t_SL g6114 ( 
.A(n_6087),
.B(n_1460),
.Y(n_6114)
);

AOI321xp33_ASAP7_75t_L g6115 ( 
.A1(n_6099),
.A2(n_1463),
.A3(n_1467),
.B1(n_1461),
.B2(n_1462),
.C(n_1465),
.Y(n_6115)
);

AOI22xp5_ASAP7_75t_L g6116 ( 
.A1(n_6092),
.A2(n_6071),
.B1(n_6107),
.B2(n_6082),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_6074),
.Y(n_6117)
);

AOI22xp33_ASAP7_75t_L g6118 ( 
.A1(n_6090),
.A2(n_1469),
.B1(n_1465),
.B2(n_1468),
.Y(n_6118)
);

OAI21xp33_ASAP7_75t_SL g6119 ( 
.A1(n_6073),
.A2(n_1469),
.B(n_1472),
.Y(n_6119)
);

OAI22xp5_ASAP7_75t_L g6120 ( 
.A1(n_6088),
.A2(n_1479),
.B1(n_1473),
.B2(n_1477),
.Y(n_6120)
);

AOI22xp5_ASAP7_75t_L g6121 ( 
.A1(n_6070),
.A2(n_1480),
.B1(n_1477),
.B2(n_1479),
.Y(n_6121)
);

AND2x2_ASAP7_75t_L g6122 ( 
.A(n_6085),
.B(n_1481),
.Y(n_6122)
);

OAI221xp5_ASAP7_75t_L g6123 ( 
.A1(n_6075),
.A2(n_1744),
.B1(n_1732),
.B2(n_1484),
.C(n_1481),
.Y(n_6123)
);

AOI211xp5_ASAP7_75t_SL g6124 ( 
.A1(n_6068),
.A2(n_1485),
.B(n_1482),
.C(n_1484),
.Y(n_6124)
);

OR2x2_ASAP7_75t_L g6125 ( 
.A(n_6084),
.B(n_1486),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_6069),
.Y(n_6126)
);

NOR2xp33_ASAP7_75t_L g6127 ( 
.A(n_6105),
.B(n_1487),
.Y(n_6127)
);

AOI21xp33_ASAP7_75t_L g6128 ( 
.A1(n_6079),
.A2(n_1487),
.B(n_1488),
.Y(n_6128)
);

OAI21xp5_ASAP7_75t_SL g6129 ( 
.A1(n_6095),
.A2(n_1488),
.B(n_1489),
.Y(n_6129)
);

INVx1_ASAP7_75t_L g6130 ( 
.A(n_6104),
.Y(n_6130)
);

INVx2_ASAP7_75t_L g6131 ( 
.A(n_6094),
.Y(n_6131)
);

INVx1_ASAP7_75t_L g6132 ( 
.A(n_6101),
.Y(n_6132)
);

AOI22xp5_ASAP7_75t_L g6133 ( 
.A1(n_6086),
.A2(n_1494),
.B1(n_1492),
.B2(n_1493),
.Y(n_6133)
);

INVx1_ASAP7_75t_L g6134 ( 
.A(n_6076),
.Y(n_6134)
);

AND2x4_ASAP7_75t_L g6135 ( 
.A(n_6091),
.B(n_1494),
.Y(n_6135)
);

INVx1_ASAP7_75t_L g6136 ( 
.A(n_6102),
.Y(n_6136)
);

OR2x2_ASAP7_75t_L g6137 ( 
.A(n_6125),
.B(n_6096),
.Y(n_6137)
);

AOI221xp5_ASAP7_75t_L g6138 ( 
.A1(n_6132),
.A2(n_6089),
.B1(n_6072),
.B2(n_6106),
.C(n_6100),
.Y(n_6138)
);

OAI22xp33_ASAP7_75t_L g6139 ( 
.A1(n_6124),
.A2(n_6133),
.B1(n_6116),
.B2(n_6112),
.Y(n_6139)
);

INVx1_ASAP7_75t_L g6140 ( 
.A(n_6113),
.Y(n_6140)
);

INVx1_ASAP7_75t_L g6141 ( 
.A(n_6113),
.Y(n_6141)
);

NOR2x1_ASAP7_75t_L g6142 ( 
.A(n_6130),
.B(n_6093),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_6122),
.Y(n_6143)
);

OAI22xp33_ASAP7_75t_L g6144 ( 
.A1(n_6110),
.A2(n_6083),
.B1(n_6098),
.B2(n_6097),
.Y(n_6144)
);

INVx1_ASAP7_75t_L g6145 ( 
.A(n_6135),
.Y(n_6145)
);

INVx1_ASAP7_75t_L g6146 ( 
.A(n_6127),
.Y(n_6146)
);

NOR2x1_ASAP7_75t_L g6147 ( 
.A(n_6114),
.B(n_6108),
.Y(n_6147)
);

INVx2_ASAP7_75t_L g6148 ( 
.A(n_6131),
.Y(n_6148)
);

INVx1_ASAP7_75t_L g6149 ( 
.A(n_6117),
.Y(n_6149)
);

INVx1_ASAP7_75t_L g6150 ( 
.A(n_6126),
.Y(n_6150)
);

AOI22xp5_ASAP7_75t_L g6151 ( 
.A1(n_6134),
.A2(n_6109),
.B1(n_6103),
.B2(n_1497),
.Y(n_6151)
);

INVx1_ASAP7_75t_L g6152 ( 
.A(n_6115),
.Y(n_6152)
);

AO22x2_ASAP7_75t_L g6153 ( 
.A1(n_6120),
.A2(n_1497),
.B1(n_1495),
.B2(n_1496),
.Y(n_6153)
);

NOR2x1_ASAP7_75t_L g6154 ( 
.A(n_6140),
.B(n_6123),
.Y(n_6154)
);

NOR2x1_ASAP7_75t_L g6155 ( 
.A(n_6141),
.B(n_6129),
.Y(n_6155)
);

NAND4xp75_ASAP7_75t_L g6156 ( 
.A(n_6142),
.B(n_6147),
.C(n_6138),
.D(n_6149),
.Y(n_6156)
);

NOR4xp25_ASAP7_75t_L g6157 ( 
.A(n_6144),
.B(n_6111),
.C(n_6119),
.D(n_6136),
.Y(n_6157)
);

AND2x2_ASAP7_75t_SL g6158 ( 
.A(n_6137),
.B(n_6118),
.Y(n_6158)
);

AOI22xp5_ASAP7_75t_L g6159 ( 
.A1(n_6152),
.A2(n_6121),
.B1(n_6128),
.B2(n_1501),
.Y(n_6159)
);

INVx1_ASAP7_75t_L g6160 ( 
.A(n_6153),
.Y(n_6160)
);

NAND2x1p5_ASAP7_75t_L g6161 ( 
.A(n_6143),
.B(n_6145),
.Y(n_6161)
);

NOR2x1_ASAP7_75t_L g6162 ( 
.A(n_6139),
.B(n_1498),
.Y(n_6162)
);

OR2x2_ASAP7_75t_L g6163 ( 
.A(n_6148),
.B(n_1500),
.Y(n_6163)
);

AOI21xp33_ASAP7_75t_L g6164 ( 
.A1(n_6150),
.A2(n_1502),
.B(n_1503),
.Y(n_6164)
);

INVx2_ASAP7_75t_L g6165 ( 
.A(n_6146),
.Y(n_6165)
);

OR2x2_ASAP7_75t_L g6166 ( 
.A(n_6151),
.B(n_1502),
.Y(n_6166)
);

OAI221xp5_ASAP7_75t_L g6167 ( 
.A1(n_6157),
.A2(n_1508),
.B1(n_1506),
.B2(n_1507),
.C(n_1509),
.Y(n_6167)
);

AOI221xp5_ASAP7_75t_L g6168 ( 
.A1(n_6160),
.A2(n_1511),
.B1(n_1509),
.B2(n_1510),
.C(n_1512),
.Y(n_6168)
);

AOI221xp5_ASAP7_75t_L g6169 ( 
.A1(n_6165),
.A2(n_1517),
.B1(n_1514),
.B2(n_1515),
.C(n_1518),
.Y(n_6169)
);

INVx1_ASAP7_75t_L g6170 ( 
.A(n_6163),
.Y(n_6170)
);

AOI22xp5_ASAP7_75t_L g6171 ( 
.A1(n_6156),
.A2(n_6158),
.B1(n_6155),
.B2(n_6154),
.Y(n_6171)
);

AOI21xp5_ASAP7_75t_L g6172 ( 
.A1(n_6162),
.A2(n_1515),
.B(n_1517),
.Y(n_6172)
);

OAI211xp5_ASAP7_75t_L g6173 ( 
.A1(n_6159),
.A2(n_1521),
.B(n_1519),
.C(n_1520),
.Y(n_6173)
);

AOI222xp33_ASAP7_75t_L g6174 ( 
.A1(n_6161),
.A2(n_1524),
.B1(n_1526),
.B2(n_1522),
.C1(n_1523),
.C2(n_1525),
.Y(n_6174)
);

AND2x4_ASAP7_75t_L g6175 ( 
.A(n_6170),
.B(n_6166),
.Y(n_6175)
);

NOR3xp33_ASAP7_75t_L g6176 ( 
.A(n_6167),
.B(n_6173),
.C(n_6171),
.Y(n_6176)
);

AND2x4_ASAP7_75t_L g6177 ( 
.A(n_6175),
.B(n_6172),
.Y(n_6177)
);

AND2x4_ASAP7_75t_L g6178 ( 
.A(n_6177),
.B(n_6176),
.Y(n_6178)
);

NAND3xp33_ASAP7_75t_L g6179 ( 
.A(n_6178),
.B(n_6174),
.C(n_6168),
.Y(n_6179)
);

OAI22xp5_ASAP7_75t_L g6180 ( 
.A1(n_6179),
.A2(n_6164),
.B1(n_6169),
.B2(n_1527),
.Y(n_6180)
);

OAI21xp5_ASAP7_75t_L g6181 ( 
.A1(n_6180),
.A2(n_1523),
.B(n_1526),
.Y(n_6181)
);

OAI21xp5_ASAP7_75t_L g6182 ( 
.A1(n_6181),
.A2(n_1528),
.B(n_1529),
.Y(n_6182)
);

INVx1_ASAP7_75t_L g6183 ( 
.A(n_6182),
.Y(n_6183)
);

AOI222xp33_ASAP7_75t_L g6184 ( 
.A1(n_6183),
.A2(n_1535),
.B1(n_1537),
.B2(n_1530),
.C1(n_1531),
.C2(n_1536),
.Y(n_6184)
);

AO21x2_ASAP7_75t_L g6185 ( 
.A1(n_6184),
.A2(n_1535),
.B(n_1536),
.Y(n_6185)
);

AOI221xp5_ASAP7_75t_L g6186 ( 
.A1(n_6185),
.A2(n_1541),
.B1(n_1539),
.B2(n_1540),
.C(n_1542),
.Y(n_6186)
);

AOI211xp5_ASAP7_75t_L g6187 ( 
.A1(n_6186),
.A2(n_1545),
.B(n_1542),
.C(n_1543),
.Y(n_6187)
);


endmodule