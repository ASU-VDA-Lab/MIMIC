module fake_jpeg_19180_n_244 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_244);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_244;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_47),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_0),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g112 ( 
.A(n_50),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_57),
.Y(n_101)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_20),
.B1(n_18),
.B2(n_29),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_61),
.B1(n_71),
.B2(n_78),
.Y(n_91)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_59),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_31),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_64),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_18),
.B1(n_20),
.B2(n_26),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_65),
.B(n_68),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_40),
.B(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_25),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_29),
.B1(n_34),
.B2(n_28),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_34),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_72),
.B(n_76),
.Y(n_104)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_28),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_36),
.B(n_24),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_1),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_26),
.B1(n_24),
.B2(n_23),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_26),
.B1(n_23),
.B2(n_19),
.Y(n_80)
);

AO22x1_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_38),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_36),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_4),
.B(n_6),
.Y(n_111)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_37),
.B(n_19),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_38),
.B(n_17),
.C(n_2),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_93),
.A2(n_115),
.B1(n_78),
.B2(n_60),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_38),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_93),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_61),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_70),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_84),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_109),
.B(n_52),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_3),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_6),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_111),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_74),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_119),
.B(n_127),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_124),
.B1(n_128),
.B2(n_95),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_49),
.C(n_50),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_95),
.C(n_101),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_82),
.B1(n_74),
.B2(n_54),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_56),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_125),
.A2(n_140),
.B1(n_149),
.B2(n_105),
.Y(n_164)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_131),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_67),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_88),
.B1(n_84),
.B2(n_79),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_57),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_129),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_62),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_148),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_133),
.A2(n_146),
.B1(n_112),
.B2(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_94),
.B(n_15),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_94),
.B(n_7),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_62),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_142),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_88),
.C(n_87),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_97),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_63),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

INVxp67_ASAP7_75t_SL g157 ( 
.A(n_147),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_79),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_145),
.A2(n_123),
.B1(n_121),
.B2(n_90),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_150),
.A2(n_153),
.B1(n_156),
.B2(n_145),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_163),
.C(n_141),
.Y(n_180)
);

AND2x4_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_108),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_164),
.B(n_149),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_110),
.B1(n_104),
.B2(n_96),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_105),
.B1(n_107),
.B2(n_117),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_167),
.B1(n_173),
.B2(n_125),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_99),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_168),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_99),
.C(n_106),
.Y(n_163)
);

OAI32xp33_ASAP7_75t_L g168 ( 
.A1(n_121),
.A2(n_92),
.A3(n_112),
.B1(n_102),
.B2(n_51),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_149),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_171),
.B(n_172),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_51),
.B1(n_81),
.B2(n_73),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

NOR4xp25_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_134),
.C(n_9),
.D(n_10),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_184),
.B1(n_160),
.B2(n_173),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_185),
.Y(n_211)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_180),
.B(n_187),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_164),
.B(n_155),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_142),
.C(n_130),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_188),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_140),
.B1(n_143),
.B2(n_137),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_126),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_131),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_130),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_191),
.B(n_193),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_135),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_194),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_92),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_134),
.C(n_9),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_159),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_195),
.B(n_176),
.Y(n_212)
);

AOI221xp5_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_169),
.B1(n_155),
.B2(n_166),
.C(n_171),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_198),
.B(n_199),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_179),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_189),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_190),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

NOR3xp33_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_152),
.C(n_161),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_210),
.B(n_168),
.Y(n_222)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_181),
.C(n_180),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_222),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_182),
.B(n_177),
.Y(n_216)
);

AOI322xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_155),
.A3(n_169),
.B1(n_184),
.B2(n_153),
.C1(n_178),
.C2(n_188),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_SL g228 ( 
.A(n_218),
.B(n_224),
.C(n_204),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_183),
.C(n_192),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_221),
.C(n_223),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_194),
.C(n_162),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_156),
.C(n_176),
.Y(n_223)
);

AOI31xp67_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_198),
.A3(n_212),
.B(n_199),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_227),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_217),
.A2(n_206),
.B1(n_201),
.B2(n_205),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_228),
.A2(n_215),
.B(n_216),
.Y(n_234)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_214),
.A2(n_203),
.B1(n_202),
.B2(n_197),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_221),
.C(n_223),
.Y(n_233)
);

AO21x1_ASAP7_75t_L g238 ( 
.A1(n_234),
.A2(n_229),
.B(n_232),
.Y(n_238)
);

NAND4xp25_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_161),
.C(n_222),
.D(n_197),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_235),
.A2(n_174),
.B(n_12),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_233),
.B(n_227),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_238),
.A2(n_239),
.B(n_236),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_241),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_242),
.A2(n_12),
.B(n_240),
.C(n_230),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g244 ( 
.A(n_243),
.Y(n_244)
);


endmodule