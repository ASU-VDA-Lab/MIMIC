module fake_jpeg_22552_n_235 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_235);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_235;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_4),
.B(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_28),
.B1(n_24),
.B2(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_1),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.C(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_30),
.B1(n_27),
.B2(n_26),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_50),
.B1(n_52),
.B2(n_28),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_33),
.B(n_20),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_38),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_28),
.B1(n_37),
.B2(n_32),
.Y(n_61)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_27),
.B1(n_18),
.B2(n_20),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_18),
.B1(n_20),
.B2(n_31),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_54),
.A2(n_40),
.B1(n_35),
.B2(n_15),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_60),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_65),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx5_ASAP7_75t_SL g87 ( 
.A(n_59),
.Y(n_87)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_61),
.A2(n_67),
.B1(n_21),
.B2(n_15),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_16),
.Y(n_62)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_36),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_41),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_21),
.B1(n_29),
.B2(n_4),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_75),
.Y(n_99)
);

CKINVDCx9p33_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_18),
.B1(n_25),
.B2(n_17),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_76),
.B1(n_80),
.B2(n_34),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_29),
.Y(n_73)
);

BUFx4f_ASAP7_75t_SL g74 ( 
.A(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_29),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_42),
.B(n_36),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_22),
.B1(n_31),
.B2(n_40),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_29),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_22),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_25),
.B1(n_17),
.B2(n_19),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_25),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_92),
.B1(n_96),
.B2(n_103),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_86),
.Y(n_107)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_14),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_1),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_98),
.C(n_103),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_2),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_104),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_99),
.A2(n_54),
.B1(n_68),
.B2(n_63),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_116),
.B1(n_122),
.B2(n_128),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_85),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_60),
.Y(n_111)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_65),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_117),
.Y(n_155)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_115),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_68),
.B1(n_58),
.B2(n_66),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_120),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_68),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_119),
.A2(n_104),
.B(n_91),
.Y(n_139)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_121),
.B(n_123),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_66),
.B1(n_74),
.B2(n_71),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_78),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_55),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_2),
.Y(n_126)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_70),
.B1(n_59),
.B2(n_56),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_2),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_82),
.C(n_97),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_140),
.C(n_143),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_88),
.C(n_89),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_149),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_130),
.A2(n_92),
.B1(n_98),
.B2(n_97),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_138),
.B1(n_109),
.B2(n_113),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_98),
.B1(n_91),
.B2(n_88),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_145),
.B(n_118),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_100),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_89),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_90),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_147),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_90),
.B(n_59),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_119),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_115),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_21),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_107),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_106),
.A2(n_83),
.B1(n_56),
.B2(n_105),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_127),
.B1(n_120),
.B2(n_83),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_166),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_110),
.Y(n_159)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_106),
.Y(n_161)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_173),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_168),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_143),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_112),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_178)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_109),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_131),
.A2(n_21),
.B1(n_4),
.B2(n_5),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_131),
.A2(n_145),
.B1(n_140),
.B2(n_136),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_21),
.B1(n_5),
.B2(n_7),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_3),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_174),
.A2(n_148),
.B1(n_142),
.B2(n_146),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_157),
.B(n_138),
.Y(n_175)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_182),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_144),
.C(n_150),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_160),
.C(n_156),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_164),
.B1(n_163),
.B2(n_174),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_151),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g184 ( 
.A(n_168),
.Y(n_184)
);

INVx11_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_187),
.C(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_191),
.B(n_198),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_188),
.A2(n_159),
.B(n_171),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_197),
.Y(n_204)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_195),
.Y(n_209)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_170),
.B1(n_166),
.B2(n_161),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_178),
.A2(n_162),
.B1(n_165),
.B2(n_173),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_172),
.B1(n_141),
.B2(n_154),
.Y(n_199)
);

OAI21x1_ASAP7_75t_SL g202 ( 
.A1(n_199),
.A2(n_200),
.B(n_183),
.Y(n_202)
);

INVx2_ASAP7_75t_R g200 ( 
.A(n_181),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_141),
.C(n_151),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_186),
.C(n_7),
.Y(n_207)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_207),
.C(n_211),
.Y(n_213)
);

XNOR2x1_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_182),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_192),
.B(n_194),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_3),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_210),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_7),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_8),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_204),
.B(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_207),
.B(n_190),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_215),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_196),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_195),
.B1(n_196),
.B2(n_199),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_220),
.A2(n_203),
.B(n_197),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_222),
.A2(n_218),
.B(n_213),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_224),
.A2(n_225),
.B(n_221),
.Y(n_228)
);

OAI21x1_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_206),
.B(n_211),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_198),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_229),
.C(n_230),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_193),
.C(n_217),
.Y(n_229)
);

AO22x1_ASAP7_75t_L g232 ( 
.A1(n_228),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_232),
.A2(n_11),
.B(n_12),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_233),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_231),
.Y(n_235)
);


endmodule