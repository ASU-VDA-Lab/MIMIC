module fake_aes_8255_n_706 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_706);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_706;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_638;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_30), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_72), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_33), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_42), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_31), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_35), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_61), .Y(n_85) );
CKINVDCx14_ASAP7_75t_R g86 ( .A(n_6), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_75), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_11), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_54), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_65), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_39), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_68), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_78), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_7), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_29), .Y(n_95) );
INVx1_ASAP7_75t_SL g96 ( .A(n_36), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g97 ( .A(n_10), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_4), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_76), .Y(n_99) );
INVxp33_ASAP7_75t_L g100 ( .A(n_38), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_26), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_51), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_12), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_64), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_25), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_3), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_21), .Y(n_107) );
NOR2xp67_ASAP7_75t_L g108 ( .A(n_52), .B(n_46), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_24), .Y(n_110) );
INVxp33_ASAP7_75t_SL g111 ( .A(n_13), .Y(n_111) );
INVxp33_ASAP7_75t_L g112 ( .A(n_59), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_60), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_48), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_70), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_9), .Y(n_116) );
INVxp33_ASAP7_75t_SL g117 ( .A(n_73), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_71), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_13), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_1), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_50), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_16), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_12), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_49), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_15), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_23), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_41), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_115), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_109), .Y(n_129) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_79), .A2(n_28), .B(n_74), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_86), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_79), .Y(n_132) );
INVx5_ASAP7_75t_L g133 ( .A(n_115), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g134 ( .A1(n_97), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_83), .B(n_2), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_83), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_109), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_91), .Y(n_138) );
AND2x6_ASAP7_75t_L g139 ( .A(n_80), .B(n_32), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_111), .B(n_3), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_89), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_91), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_99), .B(n_4), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_118), .Y(n_144) );
BUFx3_ASAP7_75t_L g145 ( .A(n_127), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_99), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_94), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_114), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_80), .Y(n_149) );
XNOR2xp5_ASAP7_75t_L g150 ( .A(n_107), .B(n_5), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_114), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_88), .B(n_5), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_88), .Y(n_153) );
BUFx2_ASAP7_75t_L g154 ( .A(n_98), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_98), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_103), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_81), .B(n_6), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_84), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_81), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_103), .Y(n_160) );
INVx1_ASAP7_75t_SL g161 ( .A(n_100), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_117), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_106), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_106), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_85), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_85), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_116), .B(n_7), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_92), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_104), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_116), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_119), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_142), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_142), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_152), .B(n_119), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_165), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_165), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_161), .B(n_112), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_154), .B(n_120), .Y(n_178) );
AND2x4_ASAP7_75t_SL g179 ( .A(n_160), .B(n_120), .Y(n_179) );
INVx6_ASAP7_75t_L g180 ( .A(n_133), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_168), .B(n_127), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_154), .B(n_125), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_165), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_165), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_164), .A2(n_125), .B1(n_122), .B2(n_123), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_165), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_152), .Y(n_187) );
BUFx2_ASAP7_75t_L g188 ( .A(n_147), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_142), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_142), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_142), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_141), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_168), .B(n_126), .Y(n_193) );
BUFx2_ASAP7_75t_L g194 ( .A(n_147), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_131), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_152), .B(n_122), .Y(n_196) );
BUFx2_ASAP7_75t_L g197 ( .A(n_131), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_148), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_148), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_148), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_148), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_167), .B(n_123), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_148), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_169), .B(n_126), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_128), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_128), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_130), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_156), .B(n_124), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_169), .B(n_124), .Y(n_209) );
BUFx2_ASAP7_75t_L g210 ( .A(n_170), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_128), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_130), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_171), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_158), .B(n_121), .Y(n_214) );
INVxp67_ASAP7_75t_L g215 ( .A(n_141), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_158), .B(n_121), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_153), .Y(n_217) );
AO22x2_ASAP7_75t_L g218 ( .A1(n_167), .A2(n_113), .B1(n_110), .B2(n_105), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_163), .B(n_113), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_128), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_128), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_136), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_167), .B(n_110), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_153), .B(n_95), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_136), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_145), .B(n_95), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_162), .B(n_105), .Y(n_227) );
INVx2_ASAP7_75t_SL g228 ( .A(n_145), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_138), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_162), .B(n_87), .Y(n_230) );
INVx4_ASAP7_75t_L g231 ( .A(n_139), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_153), .Y(n_232) );
BUFx3_ASAP7_75t_L g233 ( .A(n_139), .Y(n_233) );
NAND2x1p5_ASAP7_75t_L g234 ( .A(n_132), .B(n_102), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_155), .B(n_87), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_178), .B(n_155), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_218), .A2(n_140), .B1(n_134), .B2(n_149), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_218), .A2(n_132), .B1(n_149), .B2(n_139), .Y(n_238) );
INVxp67_ASAP7_75t_SL g239 ( .A(n_234), .Y(n_239) );
NAND2xp33_ASAP7_75t_SL g240 ( .A(n_231), .B(n_144), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_178), .B(n_155), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_217), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_177), .B(n_166), .Y(n_243) );
NOR2xp33_ASAP7_75t_R g244 ( .A(n_192), .B(n_144), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_217), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_178), .B(n_150), .Y(n_246) );
AND3x1_ASAP7_75t_SL g247 ( .A(n_185), .B(n_129), .C(n_137), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_233), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_232), .Y(n_249) );
NOR2xp33_ASAP7_75t_R g250 ( .A(n_192), .B(n_139), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_233), .Y(n_251) );
NOR2xp33_ASAP7_75t_R g252 ( .A(n_188), .B(n_139), .Y(n_252) );
BUFx3_ASAP7_75t_L g253 ( .A(n_231), .Y(n_253) );
BUFx8_ASAP7_75t_SL g254 ( .A(n_210), .Y(n_254) );
BUFx4f_ASAP7_75t_L g255 ( .A(n_182), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_232), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_234), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_234), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_235), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_182), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_182), .B(n_166), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_205), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_231), .Y(n_263) );
NOR2xp33_ASAP7_75t_R g264 ( .A(n_188), .B(n_139), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_228), .B(n_159), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_235), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_228), .B(n_159), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_209), .B(n_157), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g269 ( .A1(n_181), .A2(n_143), .B(n_135), .C(n_146), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_235), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_207), .Y(n_271) );
OR2x6_ASAP7_75t_L g272 ( .A(n_194), .B(n_150), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_187), .Y(n_273) );
BUFx8_ASAP7_75t_L g274 ( .A(n_210), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_194), .Y(n_275) );
NOR3xp33_ASAP7_75t_L g276 ( .A(n_213), .B(n_82), .C(n_93), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_235), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_187), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_218), .A2(n_139), .B1(n_146), .B2(n_151), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_223), .B(n_151), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_187), .Y(n_281) );
O2A1O1Ixp33_ASAP7_75t_L g282 ( .A1(n_193), .A2(n_138), .B(n_102), .C(n_101), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_207), .Y(n_283) );
NOR2xp33_ASAP7_75t_R g284 ( .A(n_195), .B(n_8), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_224), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_223), .B(n_133), .Y(n_286) );
INVx5_ASAP7_75t_L g287 ( .A(n_180), .Y(n_287) );
OR2x6_ASAP7_75t_L g288 ( .A(n_215), .B(n_90), .Y(n_288) );
BUFx12f_ASAP7_75t_L g289 ( .A(n_195), .Y(n_289) );
OR2x6_ASAP7_75t_L g290 ( .A(n_197), .B(n_90), .Y(n_290) );
NOR2xp33_ASAP7_75t_R g291 ( .A(n_197), .B(n_8), .Y(n_291) );
CKINVDCx8_ASAP7_75t_R g292 ( .A(n_213), .Y(n_292) );
INVx6_ASAP7_75t_L g293 ( .A(n_174), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_222), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_205), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_179), .B(n_133), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_206), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_223), .B(n_133), .Y(n_298) );
NAND2x1p5_ASAP7_75t_L g299 ( .A(n_202), .B(n_101), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_223), .B(n_133), .Y(n_300) );
INVx4_ASAP7_75t_L g301 ( .A(n_174), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_222), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_206), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_174), .Y(n_304) );
AOI21x1_ASAP7_75t_L g305 ( .A1(n_245), .A2(n_218), .B(n_175), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_259), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_275), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_270), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_266), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_239), .A2(n_202), .B1(n_196), .B2(n_174), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_255), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_268), .A2(n_196), .B(n_207), .Y(n_312) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_255), .A2(n_230), .B1(n_214), .B2(n_227), .Y(n_313) );
INVx2_ASAP7_75t_SL g314 ( .A(n_257), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_258), .Y(n_315) );
OAI222xp33_ASAP7_75t_L g316 ( .A1(n_272), .A2(n_196), .B1(n_202), .B2(n_204), .C1(n_224), .C2(n_226), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_299), .A2(n_196), .B1(n_179), .B2(n_216), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_236), .B(n_208), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_270), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_277), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_238), .B(n_207), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_260), .A2(n_208), .B1(n_219), .B2(n_229), .Y(n_322) );
INVx2_ASAP7_75t_SL g323 ( .A(n_293), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_304), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_260), .B(n_219), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_236), .B(n_229), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_275), .B(n_225), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_236), .B(n_225), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_285), .Y(n_329) );
OR2x6_ASAP7_75t_L g330 ( .A(n_301), .B(n_212), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_304), .B(n_207), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_293), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_241), .B(n_212), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_241), .B(n_212), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_243), .B(n_212), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_290), .B(n_96), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_261), .B(n_212), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_301), .B(n_108), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_290), .B(n_9), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_293), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_247), .A2(n_175), .B1(n_183), .B2(n_184), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_299), .B(n_133), .Y(n_342) );
INVxp67_ASAP7_75t_L g343 ( .A(n_290), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_288), .B(n_10), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_246), .B(n_130), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_271), .Y(n_346) );
INVx5_ASAP7_75t_L g347 ( .A(n_248), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_289), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_289), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_288), .B(n_130), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_253), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_238), .B(n_11), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_284), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_288), .B(n_14), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_273), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_251), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_284), .Y(n_357) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_271), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_345), .B(n_237), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_349), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g361 ( .A1(n_312), .A2(n_279), .B(n_249), .Y(n_361) );
AOI21x1_ASAP7_75t_L g362 ( .A1(n_350), .A2(n_211), .B(n_220), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_339), .A2(n_272), .B1(n_276), .B2(n_244), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_358), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_314), .B(n_273), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_307), .B(n_272), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_339), .A2(n_244), .B1(n_291), .B2(n_274), .Y(n_367) );
OAI222xp33_ASAP7_75t_L g368 ( .A1(n_339), .A2(n_292), .B1(n_247), .B2(n_291), .C1(n_280), .C2(n_282), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_306), .Y(n_369) );
OAI21x1_ASAP7_75t_L g370 ( .A1(n_321), .A2(n_269), .B(n_286), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_358), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_349), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_309), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_335), .A2(n_271), .B(n_283), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_344), .A2(n_265), .B1(n_267), .B2(n_256), .Y(n_375) );
XOR2xp5_ASAP7_75t_L g376 ( .A(n_317), .B(n_254), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_327), .B(n_278), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_320), .Y(n_378) );
OAI222xp33_ASAP7_75t_L g379 ( .A1(n_344), .A2(n_254), .B1(n_296), .B2(n_274), .C1(n_281), .C2(n_249), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_344), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_348), .Y(n_381) );
NAND2x1p5_ASAP7_75t_L g382 ( .A(n_314), .B(n_248), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_327), .B(n_294), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_325), .A2(n_240), .B1(n_264), .B2(n_252), .Y(n_384) );
O2A1O1Ixp33_ASAP7_75t_L g385 ( .A1(n_316), .A2(n_242), .B(n_256), .C(n_300), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_358), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_325), .A2(n_240), .B1(n_264), .B2(n_252), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_325), .B(n_242), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_352), .A2(n_250), .B1(n_302), .B2(n_294), .Y(n_389) );
A2O1A1Ixp33_ASAP7_75t_L g390 ( .A1(n_345), .A2(n_302), .B(n_298), .C(n_263), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_343), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_364), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_359), .B(n_329), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_363), .A2(n_352), .B1(n_353), .B2(n_354), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_369), .Y(n_395) );
OAI221xp5_ASAP7_75t_SL g396 ( .A1(n_367), .A2(n_313), .B1(n_322), .B2(n_353), .C(n_318), .Y(n_396) );
AO21x2_ASAP7_75t_L g397 ( .A1(n_362), .A2(n_321), .B(n_341), .Y(n_397) );
OAI211xp5_ASAP7_75t_L g398 ( .A1(n_376), .A2(n_336), .B(n_357), .C(n_332), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_364), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_379), .B(n_311), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_359), .B(n_315), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g402 ( .A1(n_375), .A2(n_310), .B1(n_315), .B2(n_338), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_375), .A2(n_358), .B(n_346), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_369), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_368), .A2(n_338), .B1(n_328), .B2(n_311), .C(n_326), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_380), .A2(n_338), .B1(n_250), .B2(n_324), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_383), .B(n_328), .Y(n_407) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_385), .A2(n_337), .B(n_333), .Y(n_408) );
INVxp67_ASAP7_75t_L g409 ( .A(n_366), .Y(n_409) );
BUFx4f_ASAP7_75t_SL g410 ( .A(n_366), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_376), .A2(n_340), .B1(n_323), .B2(n_334), .C(n_319), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_360), .B(n_323), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_383), .B(n_373), .Y(n_413) );
BUFx6f_ASAP7_75t_SL g414 ( .A(n_365), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_373), .A2(n_324), .B1(n_308), .B2(n_319), .Y(n_415) );
AO21x1_ASAP7_75t_L g416 ( .A1(n_361), .A2(n_305), .B(n_331), .Y(n_416) );
AOI22xp33_ASAP7_75t_SL g417 ( .A1(n_372), .A2(n_308), .B1(n_319), .B2(n_340), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_378), .B(n_308), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_378), .A2(n_331), .B1(n_355), .B2(n_330), .Y(n_419) );
OAI22xp33_ASAP7_75t_L g420 ( .A1(n_388), .A2(n_330), .B1(n_305), .B2(n_351), .Y(n_420) );
BUFx2_ASAP7_75t_L g421 ( .A(n_392), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_392), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_395), .B(n_371), .Y(n_423) );
NOR5xp2_ASAP7_75t_SL g424 ( .A(n_405), .B(n_390), .C(n_15), .D(n_16), .E(n_17), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_402), .A2(n_387), .B1(n_384), .B2(n_389), .Y(n_425) );
AND2x4_ASAP7_75t_SL g426 ( .A(n_413), .B(n_365), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_395), .Y(n_427) );
AOI22xp33_ASAP7_75t_SL g428 ( .A1(n_411), .A2(n_391), .B1(n_365), .B2(n_381), .Y(n_428) );
BUFx2_ASAP7_75t_L g429 ( .A(n_392), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_413), .B(n_361), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_404), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_401), .B(n_377), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_405), .A2(n_365), .B1(n_331), .B2(n_330), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_410), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_404), .B(n_370), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_398), .B(n_330), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_393), .B(n_370), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_411), .A2(n_356), .B1(n_351), .B2(n_342), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_407), .B(n_382), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_418), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_399), .Y(n_441) );
NAND4xp25_ASAP7_75t_SL g442 ( .A(n_394), .B(n_14), .C(n_17), .D(n_18), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_407), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_399), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_418), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_400), .B(n_18), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_393), .B(n_382), .Y(n_447) );
BUFx3_ASAP7_75t_L g448 ( .A(n_399), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_416), .Y(n_449) );
OAI22xp33_ASAP7_75t_L g450 ( .A1(n_409), .A2(n_347), .B1(n_356), .B2(n_351), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_396), .B(n_374), .C(n_347), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_412), .A2(n_186), .B1(n_176), .B2(n_183), .C(n_184), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_419), .B(n_386), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_416), .Y(n_454) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_408), .A2(n_186), .B1(n_176), .B2(n_203), .C(n_190), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_427), .Y(n_456) );
INVx4_ASAP7_75t_L g457 ( .A(n_426), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_448), .Y(n_458) );
BUFx3_ASAP7_75t_L g459 ( .A(n_434), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_443), .B(n_397), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_430), .B(n_397), .Y(n_461) );
NAND4xp25_ASAP7_75t_L g462 ( .A(n_446), .B(n_417), .C(n_415), .D(n_403), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_422), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_432), .B(n_414), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_430), .B(n_397), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_427), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_442), .A2(n_425), .B1(n_428), .B2(n_433), .Y(n_467) );
INVxp67_ASAP7_75t_L g468 ( .A(n_439), .Y(n_468) );
NOR2xp67_ASAP7_75t_L g469 ( .A(n_449), .B(n_403), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_431), .Y(n_470) );
NAND2xp33_ASAP7_75t_L g471 ( .A(n_432), .B(n_364), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_426), .A2(n_414), .B1(n_406), .B2(n_420), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_431), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_438), .A2(n_414), .B1(n_386), .B2(n_371), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_440), .B(n_397), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_440), .B(n_408), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_422), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_422), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_447), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_445), .B(n_19), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_445), .B(n_362), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_447), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_435), .B(n_371), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_448), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_426), .A2(n_414), .B1(n_386), .B2(n_347), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_435), .B(n_19), .Y(n_486) );
CKINVDCx16_ASAP7_75t_R g487 ( .A(n_439), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_437), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_441), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_436), .B(n_20), .Y(n_490) );
AOI221xp5_ASAP7_75t_L g491 ( .A1(n_449), .A2(n_454), .B1(n_451), .B2(n_423), .C(n_453), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_423), .B(n_20), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_441), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_444), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_450), .A2(n_220), .B(n_211), .C(n_221), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_444), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_453), .A2(n_347), .B1(n_364), .B2(n_271), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_423), .B(n_21), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_423), .B(n_364), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_421), .B(n_364), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_421), .B(n_221), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_451), .B(n_22), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_429), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_429), .B(n_27), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_456), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_463), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_456), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_463), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_466), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_465), .B(n_475), .Y(n_510) );
INVx3_ASAP7_75t_SL g511 ( .A(n_457), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_479), .B(n_454), .Y(n_512) );
INVx5_ASAP7_75t_L g513 ( .A(n_457), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_482), .B(n_448), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_490), .A2(n_452), .B(n_455), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_465), .B(n_172), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_466), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_470), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_470), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_475), .B(n_172), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_487), .B(n_424), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_483), .B(n_173), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_473), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_487), .B(n_424), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_473), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_483), .B(n_173), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_461), .B(n_488), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_493), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_493), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_496), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_461), .B(n_199), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_459), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_488), .B(n_199), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_486), .B(n_203), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_503), .B(n_201), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_503), .B(n_201), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_496), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_459), .B(n_34), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_477), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_477), .B(n_200), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_478), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_478), .B(n_200), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_492), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_468), .B(n_198), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_492), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_460), .B(n_198), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_464), .B(n_191), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_489), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_481), .B(n_494), .Y(n_549) );
NAND3xp33_ASAP7_75t_L g550 ( .A(n_467), .B(n_189), .C(n_190), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_480), .B(n_37), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_481), .B(n_191), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_489), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_494), .B(n_458), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_460), .B(n_476), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_504), .Y(n_556) );
OAI31xp33_ASAP7_75t_SL g557 ( .A1(n_502), .A2(n_40), .A3(n_43), .B(n_44), .Y(n_557) );
BUFx2_ASAP7_75t_SL g558 ( .A(n_457), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_484), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_504), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_500), .B(n_189), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_484), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_511), .A2(n_472), .B1(n_485), .B2(n_491), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_505), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_505), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_507), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_507), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_509), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_510), .B(n_498), .Y(n_569) );
OA21x2_ASAP7_75t_L g570 ( .A1(n_521), .A2(n_469), .B(n_497), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_513), .A2(n_471), .B(n_474), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_509), .Y(n_572) );
OAI322xp33_ASAP7_75t_L g573 ( .A1(n_555), .A2(n_501), .A3(n_485), .B1(n_497), .B2(n_484), .C1(n_499), .C2(n_500), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_511), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_517), .Y(n_575) );
NAND2xp67_ASAP7_75t_L g576 ( .A(n_524), .B(n_499), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_510), .B(n_462), .Y(n_577) );
NAND4xp25_ASAP7_75t_L g578 ( .A(n_550), .B(n_469), .C(n_501), .D(n_495), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_517), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_527), .B(n_189), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_523), .Y(n_581) );
INVx1_ASAP7_75t_SL g582 ( .A(n_511), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_523), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_558), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_558), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_525), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_554), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_527), .B(n_45), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_525), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_551), .A2(n_189), .B1(n_283), .B2(n_346), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_543), .B(n_189), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_545), .B(n_47), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_532), .B(n_53), .Y(n_593) );
OAI21xp5_ASAP7_75t_SL g594 ( .A1(n_557), .A2(n_346), .B(n_358), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_554), .Y(n_595) );
AOI22x1_ASAP7_75t_L g596 ( .A1(n_556), .A2(n_346), .B1(n_56), .B2(n_57), .Y(n_596) );
OAI32xp33_ASAP7_75t_L g597 ( .A1(n_560), .A2(n_55), .A3(n_58), .B1(n_62), .B2(n_63), .Y(n_597) );
INVx2_ASAP7_75t_SL g598 ( .A(n_513), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_518), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_519), .Y(n_600) );
AOI32xp33_ASAP7_75t_L g601 ( .A1(n_538), .A2(n_66), .A3(n_67), .B1(n_69), .B2(n_77), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_555), .B(n_283), .Y(n_602) );
AOI221xp5_ASAP7_75t_SL g603 ( .A1(n_515), .A2(n_303), .B1(n_297), .B2(n_295), .C(n_262), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_528), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_513), .B(n_283), .Y(n_605) );
OAI21xp33_ASAP7_75t_L g606 ( .A1(n_562), .A2(n_303), .B(n_297), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_513), .A2(n_287), .B(n_248), .Y(n_607) );
AOI21xp33_ASAP7_75t_SL g608 ( .A1(n_514), .A2(n_262), .B(n_295), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_513), .A2(n_287), .B1(n_253), .B2(n_263), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_549), .B(n_287), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_549), .B(n_287), .Y(n_611) );
OAI22xp33_ASAP7_75t_L g612 ( .A1(n_513), .A2(n_248), .B1(n_180), .B2(n_251), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_L g613 ( .A1(n_547), .A2(n_180), .B(n_544), .C(n_534), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_599), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_600), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_577), .B(n_528), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_587), .B(n_516), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_595), .B(n_512), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_564), .B(n_529), .Y(n_619) );
XNOR2xp5_ASAP7_75t_L g620 ( .A(n_576), .B(n_516), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_569), .B(n_562), .Y(n_621) );
OAI21xp33_ASAP7_75t_L g622 ( .A1(n_594), .A2(n_512), .B(n_559), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_574), .B(n_559), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_574), .B(n_520), .Y(n_624) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_613), .A2(n_546), .B(n_531), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_563), .A2(n_531), .B1(n_520), .B2(n_552), .Y(n_626) );
OA22x2_ASAP7_75t_L g627 ( .A1(n_584), .A2(n_537), .B1(n_530), .B2(n_529), .Y(n_627) );
NOR2x1_ASAP7_75t_L g628 ( .A(n_584), .B(n_537), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_565), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_566), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_567), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_568), .B(n_530), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_572), .B(n_548), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_575), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_579), .Y(n_635) );
NOR3xp33_ASAP7_75t_L g636 ( .A(n_563), .B(n_546), .C(n_535), .Y(n_636) );
XNOR2x1_ASAP7_75t_L g637 ( .A(n_582), .B(n_526), .Y(n_637) );
NAND2xp33_ASAP7_75t_SL g638 ( .A(n_598), .B(n_553), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_604), .B(n_548), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_582), .B(n_553), .Y(n_640) );
AO22x2_ASAP7_75t_L g641 ( .A1(n_581), .A2(n_539), .B1(n_506), .B2(n_508), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_583), .B(n_539), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_586), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_585), .B(n_561), .Y(n_644) );
O2A1O1Ixp33_ASAP7_75t_L g645 ( .A1(n_608), .A2(n_533), .B(n_536), .C(n_535), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_589), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_580), .Y(n_647) );
OAI21xp33_ASAP7_75t_SL g648 ( .A1(n_585), .A2(n_552), .B(n_506), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_591), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_570), .B(n_508), .Y(n_650) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_628), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_616), .B(n_570), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_627), .Y(n_653) );
NAND4xp75_ASAP7_75t_L g654 ( .A(n_648), .B(n_603), .C(n_593), .D(n_588), .Y(n_654) );
INVx1_ASAP7_75t_SL g655 ( .A(n_637), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_621), .B(n_611), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_624), .B(n_541), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_627), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_616), .B(n_602), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_617), .B(n_610), .Y(n_660) );
OAI21xp5_ASAP7_75t_SL g661 ( .A1(n_636), .A2(n_601), .B(n_571), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_614), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_641), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_626), .A2(n_573), .B1(n_578), .B2(n_597), .C(n_592), .Y(n_664) );
AOI221xp5_ASAP7_75t_SL g665 ( .A1(n_620), .A2(n_612), .B1(n_606), .B2(n_609), .C(n_526), .Y(n_665) );
INVxp67_ASAP7_75t_L g666 ( .A(n_638), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_615), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_645), .A2(n_596), .B1(n_590), .B2(n_605), .Y(n_668) );
OAI21xp33_ASAP7_75t_L g669 ( .A1(n_622), .A2(n_522), .B(n_561), .Y(n_669) );
NOR2xp33_ASAP7_75t_SL g670 ( .A(n_625), .B(n_609), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_645), .A2(n_541), .B1(n_522), .B2(n_533), .Y(n_671) );
XNOR2xp5_ASAP7_75t_L g672 ( .A(n_644), .B(n_536), .Y(n_672) );
NOR3xp33_ASAP7_75t_L g673 ( .A(n_661), .B(n_625), .C(n_650), .Y(n_673) );
NOR3xp33_ASAP7_75t_SL g674 ( .A(n_654), .B(n_650), .C(n_647), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_662), .Y(n_675) );
AOI31xp33_ASAP7_75t_L g676 ( .A1(n_665), .A2(n_640), .A3(n_623), .B(n_618), .Y(n_676) );
NAND4xp75_ASAP7_75t_L g677 ( .A(n_664), .B(n_649), .C(n_632), .D(n_619), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_657), .Y(n_678) );
NOR2x1p5_ASAP7_75t_L g679 ( .A(n_654), .B(n_632), .Y(n_679) );
INVxp67_ASAP7_75t_L g680 ( .A(n_670), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_653), .A2(n_646), .B1(n_643), .B2(n_631), .C(n_635), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g682 ( .A1(n_666), .A2(n_639), .B1(n_642), .B2(n_633), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_655), .B(n_658), .Y(n_683) );
O2A1O1Ixp33_ASAP7_75t_L g684 ( .A1(n_651), .A2(n_629), .B(n_634), .C(n_630), .Y(n_684) );
AOI21xp33_ASAP7_75t_L g685 ( .A1(n_663), .A2(n_641), .B(n_633), .Y(n_685) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_663), .Y(n_686) );
AOI211xp5_ASAP7_75t_L g687 ( .A1(n_671), .A2(n_607), .B(n_641), .C(n_542), .Y(n_687) );
NOR3xp33_ASAP7_75t_SL g688 ( .A(n_668), .B(n_540), .C(n_542), .Y(n_688) );
OAI21xp33_ASAP7_75t_L g689 ( .A1(n_652), .A2(n_540), .B(n_180), .Y(n_689) );
AOI211xp5_ASAP7_75t_L g690 ( .A1(n_669), .A2(n_672), .B(n_659), .C(n_667), .Y(n_690) );
NOR2x1_ASAP7_75t_L g691 ( .A(n_672), .B(n_656), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_660), .B(n_657), .Y(n_692) );
NOR2x1_ASAP7_75t_L g693 ( .A(n_656), .B(n_654), .Y(n_693) );
AND2x4_ASAP7_75t_L g694 ( .A(n_691), .B(n_688), .Y(n_694) );
AOI21xp33_ASAP7_75t_SL g695 ( .A1(n_676), .A2(n_680), .B(n_673), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_683), .B(n_681), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_693), .A2(n_677), .B1(n_674), .B2(n_679), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_675), .Y(n_698) );
NAND4xp25_ASAP7_75t_L g699 ( .A(n_697), .B(n_690), .C(n_687), .D(n_689), .Y(n_699) );
NOR3xp33_ASAP7_75t_L g700 ( .A(n_695), .B(n_685), .C(n_686), .Y(n_700) );
INVxp33_ASAP7_75t_L g701 ( .A(n_694), .Y(n_701) );
XOR2xp5_ASAP7_75t_L g702 ( .A(n_701), .B(n_696), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_700), .Y(n_703) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_702), .Y(n_704) );
AOI322xp5_ASAP7_75t_L g705 ( .A1(n_704), .A2(n_703), .A3(n_682), .B1(n_685), .B2(n_699), .C1(n_698), .C2(n_678), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_705), .A2(n_684), .B(n_692), .Y(n_706) );
endmodule