module fake_jpeg_27144_n_42 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_42);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_42;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_27),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_9),
.B1(n_17),
.B2(n_16),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_19),
.B(n_0),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_8),
.C(n_15),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_30),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_7),
.B1(n_14),
.B2(n_3),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_20),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_23),
.C(n_24),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_37),
.B1(n_31),
.B2(n_35),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_34),
.B(n_2),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_1),
.A3(n_2),
.B1(n_6),
.B2(n_10),
.C1(n_18),
.C2(n_23),
.Y(n_41)
);

BUFx24_ASAP7_75t_SL g42 ( 
.A(n_41),
.Y(n_42)
);


endmodule