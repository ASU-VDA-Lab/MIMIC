module fake_ariane_669_n_2041 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2041);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2041;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_274;
wire n_337;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1769;
wire n_1632;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_928;
wire n_253;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_84),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_125),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_157),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_101),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_123),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_32),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_110),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_55),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_148),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_172),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_73),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_156),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_129),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_18),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_131),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_120),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_144),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_127),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_138),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_50),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_33),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_149),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_57),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_154),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_146),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_50),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_55),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_193),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_133),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_151),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_75),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_40),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_87),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_68),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_47),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_94),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

BUFx8_ASAP7_75t_SL g242 ( 
.A(n_176),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_59),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_121),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_74),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_29),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_171),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_152),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_6),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_194),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_38),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_24),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_184),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_99),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_98),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_113),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_124),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_136),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_122),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_29),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_0),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_45),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_86),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_15),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_104),
.Y(n_265)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_82),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_45),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_88),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_39),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_13),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_42),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_20),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_85),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_16),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_68),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_166),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_12),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_147),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_164),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_70),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g281 ( 
.A(n_160),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_70),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_196),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_183),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_169),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_78),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_47),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_22),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_49),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_181),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_54),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_10),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_83),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_135),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_117),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_72),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_43),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_27),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_97),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_12),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_57),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_90),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_79),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_66),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_73),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_111),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_159),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_36),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_34),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_48),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_182),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_13),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_9),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_58),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_4),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_81),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_17),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_3),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_62),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_14),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_167),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_2),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_58),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_72),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_52),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_18),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_62),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_60),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_61),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_54),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_37),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_191),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_6),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_177),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_0),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_153),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_126),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_61),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_1),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_71),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_77),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_30),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_71),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_35),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_108),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_19),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_32),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_27),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_37),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_163),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_60),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_145),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_23),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_140),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_65),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_33),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_40),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_30),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_190),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_178),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_187),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_28),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_118),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_39),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_64),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_11),
.Y(n_366)
);

BUFx10_ASAP7_75t_L g367 ( 
.A(n_142),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_26),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_114),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_134),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_109),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_43),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_38),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_22),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_103),
.Y(n_375)
);

BUFx5_ASAP7_75t_L g376 ( 
.A(n_20),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_44),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_179),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_63),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_165),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_36),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_102),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_192),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_49),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_44),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_96),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_199),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_5),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_69),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_132),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_56),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_150),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_139),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_11),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_170),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_180),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_116),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_376),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_242),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_376),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_376),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_376),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_376),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_267),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_376),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_264),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_264),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_377),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_264),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_209),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_235),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_355),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_264),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_355),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_240),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_264),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_296),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_248),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_296),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_296),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_296),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_211),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_296),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_206),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_250),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_339),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_339),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_339),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_339),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_339),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_293),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_365),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_299),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_365),
.Y(n_436)
);

BUFx2_ASAP7_75t_SL g437 ( 
.A(n_254),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_365),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_365),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_365),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_274),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_222),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_277),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_222),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_275),
.Y(n_445)
);

INVxp33_ASAP7_75t_SL g446 ( 
.A(n_211),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_275),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_238),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_317),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_310),
.Y(n_450)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_254),
.Y(n_451)
);

INVxp33_ASAP7_75t_L g452 ( 
.A(n_208),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_310),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_357),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_214),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_340),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_251),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_340),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_221),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_239),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_252),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_221),
.Y(n_462)
);

INVxp33_ASAP7_75t_SL g463 ( 
.A(n_214),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_243),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_255),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_255),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_258),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_258),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_311),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_261),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_311),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_371),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_246),
.Y(n_473)
);

CKINVDCx14_ASAP7_75t_R g474 ( 
.A(n_254),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_371),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_259),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_249),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_223),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_272),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_262),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_223),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_309),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_259),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_287),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_225),
.Y(n_485)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_392),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_257),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_289),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_300),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_301),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_305),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_270),
.Y(n_492)
);

INVxp33_ASAP7_75t_SL g493 ( 
.A(n_225),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_320),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_322),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_257),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_228),
.Y(n_497)
);

BUFx2_ASAP7_75t_SL g498 ( 
.A(n_257),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_323),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_278),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_271),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_331),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_335),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_279),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_280),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_338),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_282),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_342),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_228),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_347),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_229),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_349),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_279),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_278),
.Y(n_514)
);

OA21x2_ASAP7_75t_L g515 ( 
.A1(n_398),
.A2(n_216),
.B(n_202),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_434),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_496),
.B(n_260),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_434),
.Y(n_518)
);

OA21x2_ASAP7_75t_L g519 ( 
.A1(n_398),
.A2(n_220),
.B(n_217),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_422),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_434),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_487),
.A2(n_269),
.B1(n_325),
.B2(n_245),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_434),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_407),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_483),
.B(n_309),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_400),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_412),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_400),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_422),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_407),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_431),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_401),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_496),
.B(n_266),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_413),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_401),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_416),
.B(n_260),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_416),
.B(n_260),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_431),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_402),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_483),
.B(n_226),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_483),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_441),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_402),
.Y(n_543)
);

OA21x2_ASAP7_75t_L g544 ( 
.A1(n_403),
.A2(n_234),
.B(n_230),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_403),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_437),
.B(n_215),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_404),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_404),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_437),
.B(n_498),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_414),
.B(n_451),
.Y(n_550)
);

INVxp33_ASAP7_75t_SL g551 ( 
.A(n_399),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_439),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_410),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_405),
.A2(n_241),
.B(n_237),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_453),
.B(n_278),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_482),
.B(n_356),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_443),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_439),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_474),
.B(n_244),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_405),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_408),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_408),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_500),
.A2(n_236),
.B1(n_362),
.B2(n_229),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_409),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_409),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_411),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_417),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_476),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_486),
.A2(n_358),
.B1(n_362),
.B2(n_236),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_411),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_415),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_504),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_415),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_418),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_498),
.B(n_265),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_504),
.B(n_276),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_514),
.A2(n_368),
.B1(n_373),
.B2(n_372),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_418),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_513),
.B(n_358),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_513),
.B(n_215),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_449),
.A2(n_372),
.B1(n_373),
.B2(n_368),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_419),
.Y(n_582)
);

NAND2x1p5_ASAP7_75t_L g583 ( 
.A(n_459),
.B(n_201),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_419),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_446),
.A2(n_374),
.B1(n_379),
.B2(n_389),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_421),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_421),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_426),
.B(n_367),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_423),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_423),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_425),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_425),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_460),
.B(n_285),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_428),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_428),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_420),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_429),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_429),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_464),
.B(n_295),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_430),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_430),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_454),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_427),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_432),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_524),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_524),
.Y(n_606)
);

AND2x2_ASAP7_75t_SL g607 ( 
.A(n_549),
.B(n_486),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_524),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_517),
.B(n_452),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_524),
.Y(n_610)
);

OAI21xp33_ASAP7_75t_SL g611 ( 
.A1(n_533),
.A2(n_473),
.B(n_384),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_530),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_530),
.Y(n_613)
);

AND2x6_ASAP7_75t_L g614 ( 
.A(n_517),
.B(n_224),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_583),
.B(n_477),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_546),
.B(n_559),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_SL g617 ( 
.A1(n_581),
.A2(n_406),
.B1(n_435),
.B2(n_433),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_527),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_530),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_542),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_520),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_530),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_588),
.B(n_448),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_523),
.Y(n_624)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_541),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_516),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_520),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_516),
.Y(n_628)
);

INVx11_ASAP7_75t_L g629 ( 
.A(n_551),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_518),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_518),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_588),
.B(n_457),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_521),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_523),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_521),
.Y(n_635)
);

INVx5_ASAP7_75t_L g636 ( 
.A(n_520),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_575),
.B(n_461),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_562),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_541),
.B(n_470),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_523),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_541),
.B(n_480),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_562),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_561),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_523),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_561),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_561),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_541),
.Y(n_647)
);

INVx2_ASAP7_75t_SL g648 ( 
.A(n_568),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_580),
.A2(n_493),
.B1(n_463),
.B2(n_455),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_565),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_520),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_566),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_555),
.B(n_492),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_561),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_555),
.B(n_501),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_566),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_520),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_587),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_570),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_570),
.Y(n_660)
);

NAND3xp33_ASAP7_75t_L g661 ( 
.A(n_585),
.B(n_507),
.C(n_505),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_571),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_534),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_587),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_L g665 ( 
.A(n_585),
.B(n_478),
.C(n_424),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_SL g666 ( 
.A(n_553),
.B(n_374),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_587),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_587),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_591),
.Y(n_669)
);

OAI22xp33_ASAP7_75t_L g670 ( 
.A1(n_563),
.A2(n_485),
.B1(n_497),
.B2(n_481),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_591),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_SL g672 ( 
.A(n_567),
.B(n_509),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_571),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_573),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_573),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_591),
.Y(n_676)
);

INVx8_ASAP7_75t_L g677 ( 
.A(n_580),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_578),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_520),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_591),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_601),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_568),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_568),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_601),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_526),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_601),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_557),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_572),
.B(n_462),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_601),
.Y(n_689)
);

AND2x6_ASAP7_75t_L g690 ( 
.A(n_536),
.B(n_224),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_536),
.B(n_477),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_578),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_572),
.B(n_465),
.Y(n_693)
);

AND2x6_ASAP7_75t_L g694 ( 
.A(n_537),
.B(n_224),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_550),
.B(n_511),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_574),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_582),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_582),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_574),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_574),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_583),
.B(n_465),
.Y(n_701)
);

XNOR2xp5_ASAP7_75t_L g702 ( 
.A(n_522),
.B(n_379),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_569),
.A2(n_291),
.B1(n_292),
.B2(n_288),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_580),
.A2(n_353),
.B1(n_364),
.B2(n_351),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_583),
.B(n_466),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_584),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_584),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_589),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_SL g709 ( 
.A(n_596),
.B(n_367),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_589),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_572),
.B(n_466),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_572),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_564),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_537),
.B(n_391),
.C(n_389),
.Y(n_714)
);

BUFx4f_ASAP7_75t_L g715 ( 
.A(n_515),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_525),
.B(n_580),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_556),
.B(n_200),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_584),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_579),
.A2(n_381),
.B1(n_385),
.B2(n_366),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_552),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_525),
.B(n_200),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_526),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_593),
.B(n_467),
.Y(n_723)
);

NAND3xp33_ASAP7_75t_L g724 ( 
.A(n_599),
.B(n_532),
.C(n_528),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_586),
.Y(n_725)
);

AOI21x1_ASAP7_75t_L g726 ( 
.A1(n_528),
.A2(n_468),
.B(n_467),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_525),
.B(n_203),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_532),
.B(n_468),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_535),
.B(n_469),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_525),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_564),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_590),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_563),
.B(n_479),
.Y(n_733)
);

INVxp33_ASAP7_75t_L g734 ( 
.A(n_522),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_579),
.Y(n_735)
);

BUFx16f_ASAP7_75t_R g736 ( 
.A(n_602),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_535),
.B(n_469),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_590),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_586),
.Y(n_739)
);

AOI21x1_ASAP7_75t_L g740 ( 
.A1(n_539),
.A2(n_472),
.B(n_471),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_577),
.B(n_603),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_564),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_577),
.A2(n_394),
.B1(n_298),
.B2(n_304),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_579),
.B(n_203),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_586),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_579),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_595),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_595),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_604),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_540),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_515),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_539),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_543),
.B(n_394),
.C(n_308),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_576),
.Y(n_754)
);

INVx8_ASAP7_75t_L g755 ( 
.A(n_564),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_543),
.B(n_204),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_604),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_597),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_564),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_626),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_630),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_607),
.B(n_545),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_616),
.B(n_545),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_609),
.B(n_479),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_607),
.B(n_547),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_630),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_626),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_653),
.B(n_548),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_628),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_631),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_655),
.A2(n_312),
.B1(n_313),
.B2(n_297),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_628),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_623),
.B(n_548),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_682),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_631),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_609),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_633),
.Y(n_777)
);

BUFx5_ASAP7_75t_L g778 ( 
.A(n_685),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_752),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_752),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_632),
.B(n_560),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_691),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_750),
.B(n_515),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_715),
.B(n_554),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_750),
.B(n_314),
.Y(n_785)
);

BUFx8_ASAP7_75t_L g786 ( 
.A(n_733),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_635),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_638),
.Y(n_788)
);

NOR2xp67_ASAP7_75t_SL g789 ( 
.A(n_618),
.B(n_388),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_635),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_695),
.B(n_315),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_701),
.B(n_705),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_611),
.A2(n_488),
.B(n_489),
.C(n_484),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_715),
.B(n_554),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_696),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_621),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_723),
.B(n_515),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_730),
.B(n_519),
.Y(n_798)
);

OAI221xp5_ASAP7_75t_L g799 ( 
.A1(n_733),
.A2(n_324),
.B1(n_343),
.B2(n_344),
.C(n_346),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_642),
.Y(n_800)
);

AO22x2_ASAP7_75t_L g801 ( 
.A1(n_665),
.A2(n_472),
.B1(n_475),
.B2(n_471),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_715),
.B(n_204),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_672),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_751),
.A2(n_544),
.B(n_519),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_615),
.B(n_318),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_606),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_730),
.B(n_691),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_690),
.B(n_694),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_724),
.A2(n_326),
.B1(n_327),
.B2(n_319),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_620),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_606),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_L g812 ( 
.A(n_639),
.B(n_641),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_SL g813 ( 
.A(n_618),
.B(n_663),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_690),
.B(n_694),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_615),
.B(n_328),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_690),
.B(n_519),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_722),
.A2(n_649),
.B1(n_714),
.B2(n_661),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_690),
.B(n_694),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_690),
.B(n_519),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_615),
.B(n_329),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_690),
.B(n_544),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_687),
.B(n_484),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_694),
.B(n_544),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_694),
.B(n_544),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_606),
.Y(n_825)
);

AND2x2_ASAP7_75t_SL g826 ( 
.A(n_709),
.B(n_316),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_610),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_643),
.B(n_205),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_SL g829 ( 
.A(n_663),
.B(n_330),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_712),
.A2(n_333),
.B1(n_348),
.B2(n_283),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_615),
.B(n_284),
.Y(n_831)
);

OAI22xp33_ASAP7_75t_L g832 ( 
.A1(n_734),
.A2(n_502),
.B1(n_499),
.B2(n_488),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_650),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_621),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_621),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_643),
.B(n_205),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_694),
.B(n_475),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_735),
.B(n_597),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_735),
.B(n_600),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_645),
.B(n_207),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_637),
.B(n_290),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_610),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_716),
.B(n_600),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_746),
.A2(n_281),
.B1(n_273),
.B2(n_210),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_702),
.A2(n_594),
.B1(n_592),
.B2(n_604),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_650),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_645),
.B(n_207),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_716),
.B(n_303),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_717),
.B(n_375),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_716),
.B(n_383),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_652),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_746),
.B(n_721),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_666),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_614),
.B(n_212),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_614),
.B(n_212),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_610),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_646),
.B(n_213),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_646),
.B(n_213),
.Y(n_858)
);

AO22x2_ASAP7_75t_L g859 ( 
.A1(n_741),
.A2(n_499),
.B1(n_512),
.B2(n_510),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_656),
.A2(n_218),
.B1(n_219),
.B2(n_227),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_614),
.B(n_218),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_612),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_612),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_614),
.B(n_219),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_682),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_659),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_629),
.Y(n_867)
);

AO221x1_ASAP7_75t_L g868 ( 
.A1(n_670),
.A2(n_224),
.B1(n_321),
.B2(n_332),
.C(n_336),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_624),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_619),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_659),
.A2(n_662),
.B1(n_673),
.B2(n_660),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_619),
.Y(n_872)
);

INVxp67_ASAP7_75t_SL g873 ( 
.A(n_648),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_619),
.B(n_227),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_654),
.B(n_231),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_654),
.B(n_231),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_662),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_621),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_677),
.B(n_232),
.Y(n_879)
);

OR2x6_ASAP7_75t_L g880 ( 
.A(n_677),
.B(n_489),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_699),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_727),
.B(n_490),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_L g883 ( 
.A(n_658),
.B(n_232),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_658),
.B(n_664),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_699),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_700),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_728),
.A2(n_512),
.B(n_510),
.C(n_490),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_700),
.Y(n_888)
);

BUFx6f_ASAP7_75t_SL g889 ( 
.A(n_736),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_624),
.B(n_233),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_673),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_624),
.B(n_233),
.Y(n_892)
);

BUFx6f_ASAP7_75t_SL g893 ( 
.A(n_629),
.Y(n_893)
);

INVxp67_ASAP7_75t_SL g894 ( 
.A(n_648),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_702),
.A2(n_594),
.B1(n_592),
.B2(n_531),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_634),
.B(n_354),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_SL g897 ( 
.A(n_754),
.B(n_367),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_674),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_675),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_744),
.B(n_491),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_666),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_754),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_743),
.B(n_491),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_621),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_664),
.B(n_360),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_678),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_617),
.B(n_703),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_640),
.B(n_369),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_751),
.A2(n_531),
.B1(n_529),
.B2(n_538),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_751),
.A2(n_529),
.B1(n_538),
.B2(n_558),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_678),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_791),
.A2(n_683),
.B1(n_756),
.B2(n_753),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_788),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_763),
.A2(n_622),
.B(n_605),
.Y(n_914)
);

BUFx4f_ASAP7_75t_L g915 ( 
.A(n_810),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_880),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_784),
.A2(n_668),
.B(n_667),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_763),
.A2(n_644),
.B(n_640),
.C(n_667),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_880),
.B(n_640),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_800),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_907),
.A2(n_692),
.B1(n_698),
.B2(n_697),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_880),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_865),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_833),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_826),
.A2(n_704),
.B1(n_719),
.B2(n_707),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_803),
.B(n_494),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_792),
.B(n_692),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_822),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_773),
.B(n_697),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_776),
.B(n_608),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_826),
.A2(n_747),
.B1(n_758),
.B2(n_738),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_902),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_782),
.B(n_608),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_778),
.B(n_625),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_867),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_778),
.B(n_625),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_773),
.B(n_698),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_846),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_SL g939 ( 
.A1(n_799),
.A2(n_508),
.B1(n_506),
.B2(n_503),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_851),
.Y(n_940)
);

NOR3xp33_ASAP7_75t_L g941 ( 
.A(n_817),
.B(n_737),
.C(n_729),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_786),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_764),
.B(n_613),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_903),
.B(n_494),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_807),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_781),
.B(n_708),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_853),
.B(n_613),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_866),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_795),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_865),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_781),
.B(n_708),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_877),
.B(n_710),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_891),
.Y(n_953)
);

BUFx4f_ASAP7_75t_L g954 ( 
.A(n_893),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_852),
.A2(n_738),
.B1(n_758),
.B2(n_732),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_898),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_796),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_899),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_852),
.A2(n_732),
.B1(n_710),
.B2(n_748),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_893),
.Y(n_960)
);

NOR2xp67_ASAP7_75t_L g961 ( 
.A(n_901),
.B(n_688),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_786),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_R g963 ( 
.A(n_813),
.B(n_726),
.Y(n_963)
);

NAND2xp33_ASAP7_75t_L g964 ( 
.A(n_778),
.B(n_647),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_906),
.Y(n_965)
);

NAND2xp33_ASAP7_75t_L g966 ( 
.A(n_778),
.B(n_647),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_911),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_SL g968 ( 
.A1(n_805),
.A2(n_508),
.B1(n_495),
.B2(n_502),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_796),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_885),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_859),
.A2(n_706),
.B1(n_757),
.B2(n_718),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_859),
.A2(n_706),
.B1(n_757),
.B2(n_718),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_849),
.A2(n_711),
.B1(n_693),
.B2(n_671),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_886),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_760),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_886),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_761),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_762),
.B(n_668),
.Y(n_978)
);

NOR2xp67_ASAP7_75t_L g979 ( 
.A(n_831),
.B(n_726),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_761),
.Y(n_980)
);

NAND2x1p5_ASAP7_75t_L g981 ( 
.A(n_774),
.B(n_713),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_801),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_767),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_769),
.B(n_772),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_762),
.B(n_669),
.Y(n_985)
);

AND2x2_ASAP7_75t_SL g986 ( 
.A(n_897),
.B(n_495),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_765),
.A2(n_681),
.B1(n_669),
.B2(n_671),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_779),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_765),
.B(n_676),
.Y(n_989)
);

OR2x6_ASAP7_75t_L g990 ( 
.A(n_859),
.B(n_755),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_790),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_774),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_796),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_843),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_871),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_783),
.B(n_680),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_841),
.A2(n_689),
.B1(n_681),
.B2(n_684),
.Y(n_997)
);

OR2x4_ASAP7_75t_L g998 ( 
.A(n_805),
.B(n_503),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_834),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_780),
.B(n_684),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_815),
.B(n_686),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_815),
.B(n_506),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_869),
.B(n_686),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_790),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_820),
.B(n_689),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_869),
.B(n_768),
.Y(n_1006)
);

NOR2xp67_ASAP7_75t_L g1007 ( 
.A(n_831),
.B(n_740),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_834),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_820),
.B(n_832),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_881),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_848),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_806),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_888),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_850),
.B(n_713),
.Y(n_1014)
);

OR2x6_ASAP7_75t_L g1015 ( 
.A(n_801),
.B(n_755),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_889),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_811),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_868),
.A2(n_725),
.B1(n_707),
.B2(n_749),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_766),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_770),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_R g1021 ( 
.A(n_829),
.B(n_740),
.Y(n_1021)
);

NOR2x2_ASAP7_75t_L g1022 ( 
.A(n_789),
.B(n_725),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_825),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_768),
.B(n_739),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_841),
.B(n_713),
.Y(n_1025)
);

AOI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_832),
.A2(n_745),
.B(n_739),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_797),
.B(n_745),
.Y(n_1027)
);

INVxp33_ASAP7_75t_L g1028 ( 
.A(n_900),
.Y(n_1028)
);

OR2x2_ASAP7_75t_SL g1029 ( 
.A(n_889),
.B(n_442),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_771),
.B(n_731),
.Y(n_1030)
);

OAI21xp33_ASAP7_75t_SL g1031 ( 
.A1(n_882),
.A2(n_742),
.B(n_731),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_845),
.A2(n_749),
.B1(n_759),
.B2(n_742),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_900),
.B(n_731),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_827),
.B(n_742),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_882),
.B(n_442),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_837),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_842),
.B(n_759),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_856),
.Y(n_1038)
);

NOR3xp33_ASAP7_75t_SL g1039 ( 
.A(n_860),
.B(n_370),
.C(n_369),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_862),
.B(n_759),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_863),
.B(n_755),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_870),
.Y(n_1042)
);

NOR2x1_ASAP7_75t_L g1043 ( 
.A(n_879),
.B(n_341),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_834),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_872),
.B(n_775),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_801),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_845),
.A2(n_273),
.B1(n_755),
.B2(n_444),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_844),
.B(n_627),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_777),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_787),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_830),
.Y(n_1051)
);

AO22x1_ASAP7_75t_L g1052 ( 
.A1(n_808),
.A2(n_390),
.B1(n_370),
.B2(n_380),
.Y(n_1052)
);

OR2x6_ASAP7_75t_L g1053 ( 
.A(n_814),
.B(n_818),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_L g1054 ( 
.A(n_809),
.B(n_361),
.C(n_359),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_793),
.A2(n_378),
.B(n_363),
.C(n_382),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_835),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_895),
.A2(n_445),
.B1(n_458),
.B2(n_456),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_838),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_798),
.B(n_627),
.Y(n_1059)
);

INVx5_ASAP7_75t_L g1060 ( 
.A(n_835),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_895),
.B(n_444),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_884),
.B(n_812),
.Y(n_1062)
);

INVx5_ASAP7_75t_L g1063 ( 
.A(n_835),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_884),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_839),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_887),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_828),
.A2(n_445),
.B1(n_447),
.B2(n_450),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_874),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_828),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_890),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_878),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_873),
.B(n_651),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_836),
.B(n_651),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_883),
.A2(n_840),
.B1(n_836),
.B2(n_847),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1031),
.A2(n_918),
.B(n_914),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_1028),
.B(n_840),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_1009),
.A2(n_857),
.B(n_858),
.C(n_847),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_1051),
.B(n_858),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_949),
.Y(n_1079)
);

INVx4_ASAP7_75t_L g1080 ( 
.A(n_954),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_964),
.A2(n_794),
.B(n_784),
.Y(n_1081)
);

BUFx12f_ASAP7_75t_L g1082 ( 
.A(n_1016),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_929),
.A2(n_876),
.B(n_875),
.C(n_905),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_968),
.B(n_875),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_927),
.B(n_894),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_998),
.B(n_876),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_913),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_928),
.B(n_447),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_986),
.B(n_878),
.Y(n_1089)
);

AO22x1_ASAP7_75t_L g1090 ( 
.A1(n_942),
.A2(n_896),
.B1(n_908),
.B2(n_892),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_928),
.Y(n_1091)
);

INVx4_ASAP7_75t_L g1092 ( 
.A(n_954),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_932),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_935),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_927),
.A2(n_802),
.B(n_878),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_929),
.B(n_904),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_937),
.A2(n_905),
.B1(n_910),
.B2(n_909),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_937),
.A2(n_904),
.B(n_804),
.Y(n_1098)
);

CKINVDCx16_ASAP7_75t_R g1099 ( 
.A(n_960),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_919),
.B(n_904),
.Y(n_1100)
);

INVx4_ASAP7_75t_L g1101 ( 
.A(n_1060),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_946),
.A2(n_855),
.B(n_854),
.C(n_864),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_970),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_946),
.A2(n_951),
.B(n_1054),
.C(n_1068),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_957),
.Y(n_1105)
);

OAI21xp33_ASAP7_75t_L g1106 ( 
.A1(n_951),
.A2(n_861),
.B(n_386),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_932),
.Y(n_1107)
);

AOI22x1_ASAP7_75t_L g1108 ( 
.A1(n_914),
.A2(n_720),
.B1(n_651),
.B2(n_657),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1002),
.B(n_816),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1062),
.A2(n_821),
.B(n_819),
.Y(n_1110)
);

OAI21xp33_ASAP7_75t_SL g1111 ( 
.A1(n_931),
.A2(n_824),
.B(n_823),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_915),
.Y(n_1112)
);

INVxp67_ASAP7_75t_L g1113 ( 
.A(n_915),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1054),
.A2(n_393),
.B(n_395),
.C(n_450),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_995),
.B(n_910),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_974),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_944),
.B(n_926),
.Y(n_1117)
);

OA21x2_ASAP7_75t_L g1118 ( 
.A1(n_1027),
.A2(n_909),
.B(n_432),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_920),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_939),
.A2(n_386),
.B1(n_396),
.B2(n_390),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_1069),
.B(n_651),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_976),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_919),
.B(n_651),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_994),
.B(n_657),
.Y(n_1124)
);

NOR2x1_ASAP7_75t_R g1125 ( 
.A(n_962),
.B(n_380),
.Y(n_1125)
);

AO21x1_ASAP7_75t_L g1126 ( 
.A1(n_941),
.A2(n_436),
.B(n_438),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1058),
.B(n_657),
.Y(n_1127)
);

NAND2x1p5_ASAP7_75t_L g1128 ( 
.A(n_1060),
.B(n_636),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_977),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_916),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_916),
.B(n_456),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1060),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_980),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_1029),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_924),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1046),
.A2(n_720),
.B1(n_679),
.B2(n_657),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_922),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_922),
.B(n_636),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_991),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_921),
.A2(n_397),
.B1(n_387),
.B2(n_720),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_917),
.A2(n_636),
.B(n_440),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1011),
.B(n_679),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1062),
.A2(n_679),
.B(n_720),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_988),
.B(n_636),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1027),
.A2(n_720),
.B(n_679),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_933),
.B(n_636),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1065),
.B(n_952),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1072),
.A2(n_306),
.B(n_247),
.Y(n_1148)
);

NOR2x1_ASAP7_75t_R g1149 ( 
.A(n_1001),
.B(n_1060),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1004),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1001),
.A2(n_307),
.B1(n_253),
.B2(n_256),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1070),
.A2(n_558),
.B(n_2),
.C(n_3),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_938),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_1012),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_984),
.A2(n_1),
.B(n_5),
.C(n_7),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_952),
.B(n_598),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_984),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_1157)
);

BUFx4f_ASAP7_75t_L g1158 ( 
.A(n_990),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_940),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1025),
.A2(n_598),
.B(n_552),
.C(n_352),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_923),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_948),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1010),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_917),
.A2(n_302),
.B(n_350),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_945),
.B(n_263),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_963),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1035),
.B(n_598),
.Y(n_1167)
);

INVx4_ASAP7_75t_L g1168 ( 
.A(n_1063),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_945),
.B(n_598),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1013),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1039),
.Y(n_1171)
);

INVx4_ASAP7_75t_L g1172 ( 
.A(n_1063),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1061),
.B(n_955),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_R g1174 ( 
.A(n_923),
.B(n_268),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_912),
.B(n_286),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1059),
.A2(n_936),
.B(n_934),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1061),
.B(n_959),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_953),
.B(n_552),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1055),
.A2(n_8),
.B(n_10),
.C(n_14),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_1021),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1059),
.A2(n_552),
.B(n_224),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1033),
.B(n_294),
.Y(n_1182)
);

NOR3xp33_ASAP7_75t_L g1183 ( 
.A(n_1005),
.B(n_1043),
.C(n_956),
.Y(n_1183)
);

INVx6_ASAP7_75t_L g1184 ( 
.A(n_1063),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_958),
.B(n_552),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_965),
.B(n_552),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_967),
.Y(n_1187)
);

INVxp33_ASAP7_75t_SL g1188 ( 
.A(n_1074),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_975),
.B(n_16),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1006),
.A2(n_17),
.B(n_19),
.C(n_21),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_950),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_1063),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_933),
.B(n_21),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_990),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1019),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1030),
.A2(n_345),
.B(n_337),
.C(n_334),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_983),
.B(n_24),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1049),
.Y(n_1198)
);

AO32x1_ASAP7_75t_L g1199 ( 
.A1(n_982),
.A2(n_25),
.A3(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1050),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_930),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1048),
.B(n_25),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1066),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1181),
.A2(n_996),
.A3(n_1073),
.B(n_1024),
.Y(n_1204)
);

AOI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1181),
.A2(n_1007),
.B(n_979),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1100),
.B(n_943),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1085),
.A2(n_1003),
.B(n_1024),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1126),
.A2(n_1064),
.A3(n_1045),
.B(n_1020),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1188),
.A2(n_990),
.B1(n_1047),
.B2(n_925),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1098),
.A2(n_973),
.B(n_997),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_SL g1211 ( 
.A1(n_1109),
.A2(n_1015),
.B(n_989),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1084),
.A2(n_961),
.B(n_947),
.C(n_943),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1104),
.A2(n_987),
.B(n_985),
.Y(n_1213)
);

BUFx2_ASAP7_75t_R g1214 ( 
.A(n_1171),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1085),
.A2(n_1003),
.B(n_1037),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1117),
.B(n_1057),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_SL g1217 ( 
.A1(n_1149),
.A2(n_1015),
.B(n_989),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_SL g1218 ( 
.A1(n_1147),
.A2(n_1015),
.B(n_978),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1173),
.B(n_978),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1143),
.A2(n_1108),
.B(n_1176),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1145),
.A2(n_971),
.B(n_972),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1096),
.A2(n_1034),
.B(n_1040),
.Y(n_1222)
);

NAND2x1p5_ASAP7_75t_L g1223 ( 
.A(n_1158),
.B(n_969),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1119),
.Y(n_1224)
);

AND2x2_ASAP7_75t_SL g1225 ( 
.A(n_1158),
.B(n_985),
.Y(n_1225)
);

NOR4xp25_ASAP7_75t_L g1226 ( 
.A(n_1203),
.B(n_1026),
.C(n_1067),
.D(n_1038),
.Y(n_1226)
);

AOI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1090),
.A2(n_1052),
.B(n_1045),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_SL g1228 ( 
.A1(n_1097),
.A2(n_1014),
.B(n_993),
.Y(n_1228)
);

AND2x2_ASAP7_75t_SL g1229 ( 
.A(n_1166),
.B(n_947),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1100),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1091),
.Y(n_1231)
);

OAI21xp33_ASAP7_75t_SL g1232 ( 
.A1(n_1173),
.A2(n_1041),
.B(n_1023),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1177),
.A2(n_1032),
.B1(n_992),
.B2(n_1017),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1075),
.A2(n_1018),
.B(n_981),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1097),
.A2(n_1026),
.B(n_1014),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1095),
.A2(n_1071),
.B(n_1056),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1088),
.B(n_1042),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1164),
.A2(n_1041),
.B(n_1000),
.Y(n_1238)
);

NAND2xp33_ASAP7_75t_R g1239 ( 
.A(n_1174),
.B(n_1000),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1184),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1110),
.A2(n_1053),
.A3(n_1022),
.B(n_1036),
.Y(n_1241)
);

AND3x1_ASAP7_75t_SL g1242 ( 
.A(n_1135),
.B(n_41),
.C(n_42),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1078),
.B(n_1036),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1153),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1094),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1160),
.A2(n_1053),
.A3(n_1044),
.B(n_1008),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1141),
.A2(n_999),
.B(n_993),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1115),
.A2(n_100),
.A3(n_189),
.B(n_188),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1093),
.B(n_41),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1112),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1107),
.B(n_46),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1114),
.A2(n_46),
.B(n_48),
.C(n_51),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1159),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1177),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1156),
.A2(n_1118),
.B(n_1178),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_SL g1256 ( 
.A1(n_1077),
.A2(n_106),
.B(n_186),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1131),
.B(n_53),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1076),
.B(n_56),
.Y(n_1258)
);

AO22x2_ASAP7_75t_L g1259 ( 
.A1(n_1140),
.A2(n_59),
.B1(n_63),
.B2(n_64),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1121),
.B(n_65),
.Y(n_1260)
);

NOR4xp25_ASAP7_75t_L g1261 ( 
.A(n_1203),
.B(n_66),
.C(n_67),
.D(n_69),
.Y(n_1261)
);

INVx4_ASAP7_75t_L g1262 ( 
.A(n_1080),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_SL g1263 ( 
.A1(n_1120),
.A2(n_67),
.B(n_74),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1131),
.B(n_76),
.Y(n_1264)
);

AOI211x1_ASAP7_75t_L g1265 ( 
.A1(n_1189),
.A2(n_80),
.B(n_89),
.C(n_91),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1193),
.B(n_92),
.Y(n_1266)
);

CKINVDCx6p67_ASAP7_75t_R g1267 ( 
.A(n_1082),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1201),
.B(n_195),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1118),
.A2(n_93),
.B(n_95),
.Y(n_1269)
);

INVx5_ASAP7_75t_L g1270 ( 
.A(n_1184),
.Y(n_1270)
);

OA21x2_ASAP7_75t_L g1271 ( 
.A1(n_1115),
.A2(n_1167),
.B(n_1127),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1165),
.B(n_185),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1194),
.A2(n_105),
.A3(n_107),
.B(n_112),
.Y(n_1273)
);

AOI21xp33_ASAP7_75t_L g1274 ( 
.A1(n_1140),
.A2(n_115),
.B(n_119),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1130),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1111),
.A2(n_128),
.B(n_130),
.Y(n_1276)
);

NAND3xp33_ASAP7_75t_L g1277 ( 
.A(n_1179),
.B(n_1190),
.C(n_1155),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1162),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1083),
.A2(n_137),
.B(n_141),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1127),
.A2(n_143),
.B(n_158),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1086),
.A2(n_162),
.B(n_173),
.C(n_174),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1102),
.A2(n_1167),
.B(n_1124),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1187),
.B(n_1137),
.Y(n_1283)
);

NAND3xp33_ASAP7_75t_L g1284 ( 
.A(n_1157),
.B(n_1152),
.C(n_1196),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1191),
.B(n_1154),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_R g1286 ( 
.A(n_1099),
.B(n_1092),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1180),
.B(n_1144),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1124),
.A2(n_1089),
.B(n_1175),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1144),
.B(n_1146),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1161),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1113),
.B(n_1142),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1198),
.B(n_1200),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1103),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1116),
.A2(n_1129),
.A3(n_1139),
.B(n_1133),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1189),
.B(n_1197),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1125),
.Y(n_1296)
);

BUFx2_ASAP7_75t_SL g1297 ( 
.A(n_1092),
.Y(n_1297)
);

AND2x2_ASAP7_75t_SL g1298 ( 
.A(n_1138),
.B(n_1136),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1134),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1163),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1106),
.A2(n_1186),
.B(n_1185),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1185),
.A2(n_1186),
.B(n_1202),
.Y(n_1302)
);

INVx3_ASAP7_75t_SL g1303 ( 
.A(n_1184),
.Y(n_1303)
);

AOI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1183),
.A2(n_1151),
.B1(n_1182),
.B2(n_1123),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1170),
.B(n_1195),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1122),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1169),
.A2(n_1150),
.B(n_1148),
.Y(n_1307)
);

NAND2x1_ASAP7_75t_L g1308 ( 
.A(n_1101),
.B(n_1168),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1128),
.A2(n_1192),
.B(n_1132),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1128),
.A2(n_1101),
.B(n_1168),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1105),
.B(n_1172),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_SL g1312 ( 
.A1(n_1199),
.A2(n_1104),
.B(n_1077),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1188),
.A2(n_937),
.B1(n_946),
.B2(n_929),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1079),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1084),
.A2(n_791),
.B(n_1009),
.C(n_785),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1143),
.A2(n_1108),
.B(n_1181),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1098),
.A2(n_1104),
.B(n_763),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1117),
.B(n_928),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1084),
.A2(n_1104),
.B(n_791),
.C(n_1009),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1087),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1181),
.A2(n_1126),
.A3(n_1097),
.B(n_1110),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1081),
.A2(n_966),
.B(n_964),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1100),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1143),
.A2(n_1108),
.B(n_1181),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1081),
.A2(n_966),
.B(n_964),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1147),
.B(n_927),
.Y(n_1326)
);

NOR2xp67_ASAP7_75t_L g1327 ( 
.A(n_1080),
.B(n_810),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1098),
.A2(n_1104),
.B(n_763),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1117),
.B(n_928),
.Y(n_1329)
);

INVxp67_ASAP7_75t_SL g1330 ( 
.A(n_1109),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1098),
.A2(n_1104),
.B(n_763),
.Y(n_1331)
);

OAI22x1_ASAP7_75t_L g1332 ( 
.A1(n_1084),
.A2(n_1078),
.B1(n_1009),
.B2(n_702),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1143),
.A2(n_1108),
.B(n_1181),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1081),
.A2(n_966),
.B(n_964),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1181),
.A2(n_1126),
.A3(n_1097),
.B(n_1110),
.Y(n_1335)
);

AO21x1_ASAP7_75t_L g1336 ( 
.A1(n_1084),
.A2(n_1009),
.B(n_1104),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1081),
.A2(n_966),
.B(n_964),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1081),
.A2(n_966),
.B(n_964),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1143),
.A2(n_1108),
.B(n_1181),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1143),
.A2(n_1108),
.B(n_1181),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1147),
.B(n_927),
.Y(n_1341)
);

OAI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1263),
.A2(n_1313),
.B1(n_1332),
.B2(n_1254),
.Y(n_1342)
);

INVx8_ASAP7_75t_L g1343 ( 
.A(n_1270),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1316),
.A2(n_1333),
.B(n_1324),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_SL g1345 ( 
.A1(n_1319),
.A2(n_1315),
.B(n_1313),
.C(n_1326),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1292),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1204),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1204),
.Y(n_1348)
);

OR2x6_ASAP7_75t_L g1349 ( 
.A(n_1211),
.B(n_1217),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1204),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1263),
.A2(n_1279),
.B(n_1235),
.C(n_1274),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1294),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_1267),
.Y(n_1353)
);

BUFx8_ASAP7_75t_SL g1354 ( 
.A(n_1245),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1339),
.A2(n_1340),
.B(n_1220),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1279),
.A2(n_1328),
.B(n_1317),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1258),
.A2(n_1336),
.B(n_1252),
.C(n_1260),
.Y(n_1357)
);

AOI221xp5_ASAP7_75t_L g1358 ( 
.A1(n_1261),
.A2(n_1226),
.B1(n_1259),
.B2(n_1254),
.C(n_1277),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1286),
.Y(n_1359)
);

BUFx12f_ASAP7_75t_L g1360 ( 
.A(n_1290),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1271),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1322),
.A2(n_1334),
.B(n_1325),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1271),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1321),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1225),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1294),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1294),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1317),
.A2(n_1331),
.B(n_1328),
.Y(n_1368)
);

AOI221xp5_ASAP7_75t_L g1369 ( 
.A1(n_1261),
.A2(n_1226),
.B1(n_1259),
.B2(n_1277),
.C(n_1284),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1329),
.B(n_1231),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1337),
.A2(n_1338),
.B(n_1269),
.Y(n_1371)
);

A2O1A1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1235),
.A2(n_1274),
.B(n_1284),
.C(n_1272),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1303),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1331),
.B(n_1213),
.Y(n_1374)
);

OR2x6_ASAP7_75t_L g1375 ( 
.A(n_1218),
.B(n_1228),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1247),
.A2(n_1222),
.B(n_1210),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1210),
.A2(n_1236),
.B(n_1234),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1221),
.A2(n_1276),
.B(n_1215),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1209),
.A2(n_1216),
.B1(n_1295),
.B2(n_1341),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1243),
.B(n_1326),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1341),
.A2(n_1213),
.B(n_1282),
.Y(n_1381)
);

OR2x6_ASAP7_75t_L g1382 ( 
.A(n_1288),
.B(n_1219),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1282),
.A2(n_1312),
.B(n_1301),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1207),
.A2(n_1232),
.B(n_1256),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1304),
.A2(n_1212),
.B1(n_1291),
.B2(n_1209),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1283),
.B(n_1275),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1214),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1321),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1219),
.B(n_1223),
.Y(n_1389)
);

OR2x6_ASAP7_75t_L g1390 ( 
.A(n_1223),
.B(n_1287),
.Y(n_1390)
);

OA21x2_ASAP7_75t_L g1391 ( 
.A1(n_1238),
.A2(n_1280),
.B(n_1233),
.Y(n_1391)
);

CKINVDCx8_ASAP7_75t_R g1392 ( 
.A(n_1297),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1240),
.Y(n_1393)
);

BUFx3_ASAP7_75t_L g1394 ( 
.A(n_1250),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1321),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1224),
.Y(n_1396)
);

OR2x6_ASAP7_75t_L g1397 ( 
.A(n_1238),
.B(n_1233),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1309),
.A2(n_1307),
.B(n_1227),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1299),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1239),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_R g1401 ( 
.A(n_1262),
.B(n_1229),
.Y(n_1401)
);

NAND2x1p5_ASAP7_75t_L g1402 ( 
.A(n_1289),
.B(n_1230),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1307),
.A2(n_1310),
.B(n_1302),
.Y(n_1403)
);

AO31x2_ASAP7_75t_L g1404 ( 
.A1(n_1244),
.A2(n_1278),
.A3(n_1320),
.B(n_1253),
.Y(n_1404)
);

NAND2x1p5_ASAP7_75t_L g1405 ( 
.A(n_1323),
.B(n_1298),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1310),
.A2(n_1308),
.B(n_1311),
.Y(n_1406)
);

INVxp67_ASAP7_75t_SL g1407 ( 
.A(n_1237),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1264),
.A2(n_1296),
.B1(n_1266),
.B2(n_1206),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1285),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1323),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1323),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1281),
.A2(n_1251),
.B(n_1249),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1262),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1268),
.A2(n_1305),
.B(n_1306),
.Y(n_1414)
);

AO31x2_ASAP7_75t_L g1415 ( 
.A1(n_1293),
.A2(n_1314),
.A3(n_1300),
.B(n_1335),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1335),
.A2(n_1246),
.B(n_1208),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1335),
.A2(n_1246),
.B(n_1208),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1242),
.A2(n_1327),
.B1(n_1265),
.B2(n_1273),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1208),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1241),
.B(n_1246),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1248),
.A2(n_1241),
.B(n_1273),
.Y(n_1421)
);

OR2x6_ASAP7_75t_L g1422 ( 
.A(n_1273),
.B(n_1248),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1248),
.Y(n_1423)
);

OAI31xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1313),
.A2(n_1203),
.A3(n_1084),
.B(n_1254),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1316),
.A2(n_1333),
.B(n_1324),
.Y(n_1425)
);

O2A1O1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1315),
.A2(n_1319),
.B(n_791),
.C(n_1313),
.Y(n_1426)
);

AOI22x1_ASAP7_75t_L g1427 ( 
.A1(n_1317),
.A2(n_663),
.B1(n_618),
.B2(n_1171),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1204),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1318),
.B(n_1257),
.Y(n_1429)
);

OR2x6_ASAP7_75t_L g1430 ( 
.A(n_1211),
.B(n_1217),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1303),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1294),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1294),
.Y(n_1433)
);

INVx5_ASAP7_75t_L g1434 ( 
.A(n_1270),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1332),
.A2(n_1009),
.B1(n_1084),
.B2(n_1336),
.Y(n_1435)
);

BUFx4f_ASAP7_75t_L g1436 ( 
.A(n_1267),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1315),
.A2(n_1319),
.B(n_1084),
.C(n_1313),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1204),
.Y(n_1438)
);

OA21x2_ASAP7_75t_L g1439 ( 
.A1(n_1316),
.A2(n_1333),
.B(n_1324),
.Y(n_1439)
);

INVxp67_ASAP7_75t_SL g1440 ( 
.A(n_1255),
.Y(n_1440)
);

INVx4_ASAP7_75t_L g1441 ( 
.A(n_1245),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1316),
.A2(n_1333),
.B(n_1324),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1318),
.B(n_1257),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1292),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1270),
.B(n_1194),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1292),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1316),
.A2(n_1333),
.B(n_1324),
.Y(n_1447)
);

AOI221xp5_ASAP7_75t_L g1448 ( 
.A1(n_1315),
.A2(n_791),
.B1(n_670),
.B2(n_1261),
.C(n_1313),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1292),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1316),
.A2(n_1333),
.B(n_1324),
.Y(n_1450)
);

INVx2_ASAP7_75t_SL g1451 ( 
.A(n_1245),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_SL g1452 ( 
.A1(n_1336),
.A2(n_1315),
.B(n_1313),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1270),
.B(n_1194),
.Y(n_1453)
);

AO21x2_ASAP7_75t_L g1454 ( 
.A1(n_1312),
.A2(n_1279),
.B(n_1205),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1259),
.A2(n_1209),
.B1(n_986),
.B2(n_1188),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1322),
.A2(n_1334),
.B(n_1325),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1316),
.A2(n_1333),
.B(n_1324),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1316),
.A2(n_1333),
.B(n_1324),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1315),
.A2(n_791),
.B(n_1319),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1263),
.A2(n_1009),
.B1(n_1313),
.B2(n_1332),
.Y(n_1460)
);

NOR2x1_ASAP7_75t_SL g1461 ( 
.A(n_1313),
.B(n_990),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1322),
.A2(n_1334),
.B(n_1325),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1315),
.B(n_1188),
.Y(n_1463)
);

A2O1A1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1315),
.A2(n_1319),
.B(n_1084),
.C(n_1313),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1332),
.A2(n_1009),
.B1(n_1084),
.B2(n_1336),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1318),
.B(n_1257),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1316),
.A2(n_1333),
.B(n_1324),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1318),
.B(n_1257),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1231),
.Y(n_1469)
);

NAND2xp33_ASAP7_75t_R g1470 ( 
.A(n_1279),
.B(n_1188),
.Y(n_1470)
);

OAI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1315),
.A2(n_791),
.B1(n_1319),
.B2(n_1263),
.C(n_1084),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1270),
.B(n_1194),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1315),
.A2(n_791),
.B(n_1319),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1332),
.A2(n_1009),
.B1(n_1084),
.B2(n_1336),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1330),
.B(n_1318),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1316),
.A2(n_1333),
.B(n_1324),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1332),
.A2(n_1084),
.B1(n_826),
.B2(n_1188),
.Y(n_1477)
);

CKINVDCx11_ASAP7_75t_R g1478 ( 
.A(n_1267),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1275),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1332),
.A2(n_1084),
.B1(n_826),
.B2(n_1188),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1294),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1294),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1330),
.B(n_1318),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1294),
.Y(n_1484)
);

O2A1O1Ixp5_ASAP7_75t_L g1485 ( 
.A1(n_1460),
.A2(n_1342),
.B(n_1473),
.C(n_1459),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1471),
.A2(n_1464),
.B1(n_1437),
.B2(n_1448),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1437),
.A2(n_1464),
.B1(n_1351),
.B2(n_1463),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1407),
.B(n_1380),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1404),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1384),
.A2(n_1356),
.B(n_1362),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1429),
.B(n_1443),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1370),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1466),
.B(n_1468),
.Y(n_1493)
);

A2O1A1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1426),
.A2(n_1424),
.B(n_1351),
.C(n_1463),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_SL g1495 ( 
.A1(n_1372),
.A2(n_1357),
.B(n_1460),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1407),
.B(n_1379),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1479),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1456),
.A2(n_1462),
.B(n_1372),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1373),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1345),
.A2(n_1374),
.B(n_1368),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1394),
.B(n_1445),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1475),
.B(n_1483),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1479),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1441),
.B(n_1409),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1386),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1379),
.B(n_1381),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1404),
.Y(n_1507)
);

O2A1O1Ixp5_ASAP7_75t_L g1508 ( 
.A1(n_1342),
.A2(n_1374),
.B(n_1385),
.C(n_1412),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1469),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1373),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1346),
.B(n_1444),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1445),
.B(n_1453),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1478),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1345),
.A2(n_1368),
.B(n_1440),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1344),
.A2(n_1442),
.B(n_1425),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1360),
.Y(n_1516)
);

INVxp67_ASAP7_75t_L g1517 ( 
.A(n_1431),
.Y(n_1517)
);

AOI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1358),
.A2(n_1369),
.B1(n_1465),
.B2(n_1435),
.C(n_1474),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1435),
.A2(n_1474),
.B1(n_1465),
.B2(n_1477),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1431),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1446),
.B(n_1449),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1368),
.A2(n_1440),
.B(n_1371),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1391),
.A2(n_1452),
.B(n_1422),
.Y(n_1523)
);

A2O1A1Ixp33_ASAP7_75t_L g1524 ( 
.A1(n_1480),
.A2(n_1455),
.B(n_1408),
.C(n_1418),
.Y(n_1524)
);

INVxp67_ASAP7_75t_L g1525 ( 
.A(n_1451),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1396),
.Y(n_1526)
);

AOI211xp5_ASAP7_75t_L g1527 ( 
.A1(n_1470),
.A2(n_1395),
.B(n_1364),
.C(n_1388),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1391),
.A2(n_1422),
.B(n_1378),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1360),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_SL g1530 ( 
.A1(n_1375),
.A2(n_1470),
.B(n_1349),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1455),
.A2(n_1418),
.B1(n_1427),
.B2(n_1392),
.Y(n_1531)
);

AOI21x1_ASAP7_75t_SL g1532 ( 
.A1(n_1478),
.A2(n_1354),
.B(n_1436),
.Y(n_1532)
);

OA22x2_ASAP7_75t_L g1533 ( 
.A1(n_1400),
.A2(n_1390),
.B1(n_1382),
.B2(n_1349),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1397),
.B(n_1415),
.Y(n_1534)
);

BUFx12f_ASAP7_75t_L g1535 ( 
.A(n_1387),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1400),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1397),
.A2(n_1405),
.B1(n_1399),
.B2(n_1441),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1343),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1354),
.Y(n_1539)
);

O2A1O1Ixp33_ASAP7_75t_L g1540 ( 
.A1(n_1397),
.A2(n_1391),
.B(n_1359),
.C(n_1413),
.Y(n_1540)
);

NOR2xp67_ASAP7_75t_L g1541 ( 
.A(n_1434),
.B(n_1361),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1343),
.Y(n_1542)
);

O2A1O1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1390),
.A2(n_1422),
.B(n_1382),
.C(n_1393),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1436),
.Y(n_1544)
);

INVx8_ASAP7_75t_L g1545 ( 
.A(n_1343),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_SL g1546 ( 
.A1(n_1375),
.A2(n_1430),
.B(n_1382),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1447),
.A2(n_1476),
.B(n_1450),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1439),
.A2(n_1458),
.B(n_1457),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1401),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1387),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1389),
.B(n_1410),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1399),
.A2(n_1390),
.B1(n_1353),
.B2(n_1430),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1472),
.B(n_1430),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1361),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1363),
.B(n_1428),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1353),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1363),
.B(n_1347),
.Y(n_1557)
);

OA22x2_ASAP7_75t_L g1558 ( 
.A1(n_1420),
.A2(n_1472),
.B1(n_1411),
.B2(n_1414),
.Y(n_1558)
);

OAI31xp33_ASAP7_75t_L g1559 ( 
.A1(n_1402),
.A2(n_1348),
.A3(n_1350),
.B(n_1438),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1401),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1348),
.B(n_1350),
.Y(n_1561)
);

O2A1O1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1383),
.A2(n_1454),
.B(n_1423),
.C(n_1402),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_SL g1563 ( 
.A1(n_1365),
.A2(n_1383),
.B(n_1434),
.Y(n_1563)
);

O2A1O1Ixp5_ASAP7_75t_L g1564 ( 
.A1(n_1423),
.A2(n_1419),
.B(n_1352),
.C(n_1482),
.Y(n_1564)
);

O2A1O1Ixp33_ASAP7_75t_L g1565 ( 
.A1(n_1419),
.A2(n_1484),
.B(n_1352),
.C(n_1482),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1376),
.B(n_1417),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1439),
.A2(n_1432),
.B1(n_1481),
.B2(n_1366),
.Y(n_1567)
);

OA21x2_ASAP7_75t_L g1568 ( 
.A1(n_1467),
.A2(n_1355),
.B(n_1421),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1366),
.A2(n_1433),
.B1(n_1367),
.B2(n_1481),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1416),
.B(n_1377),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1403),
.B(n_1398),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1471),
.A2(n_1437),
.B1(n_1464),
.B2(n_1448),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1471),
.A2(n_1437),
.B1(n_1464),
.B2(n_1448),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1471),
.A2(n_1437),
.B1(n_1464),
.B2(n_1448),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1407),
.B(n_1380),
.Y(n_1575)
);

A2O1A1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1426),
.A2(n_1315),
.B(n_1448),
.C(n_1424),
.Y(n_1576)
);

O2A1O1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1471),
.A2(n_1315),
.B(n_1319),
.C(n_1437),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1429),
.B(n_1443),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1471),
.A2(n_1437),
.B1(n_1464),
.B2(n_1448),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1441),
.B(n_813),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1344),
.A2(n_1442),
.B(n_1425),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1429),
.B(n_1443),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1344),
.A2(n_1442),
.B(n_1425),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1429),
.B(n_1443),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1471),
.A2(n_1437),
.B1(n_1464),
.B2(n_1448),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1471),
.A2(n_1437),
.B1(n_1464),
.B2(n_1448),
.Y(n_1586)
);

AOI21xp5_ASAP7_75t_SL g1587 ( 
.A1(n_1426),
.A2(n_1315),
.B(n_1319),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1471),
.A2(n_1437),
.B1(n_1464),
.B2(n_1448),
.Y(n_1588)
);

INVxp67_ASAP7_75t_SL g1589 ( 
.A(n_1361),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1407),
.B(n_1380),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1394),
.B(n_1461),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1429),
.B(n_1443),
.Y(n_1592)
);

AOI31xp33_ASAP7_75t_L g1593 ( 
.A1(n_1455),
.A2(n_1460),
.A3(n_1448),
.B(n_1342),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1406),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1407),
.B(n_1380),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_SL g1596 ( 
.A1(n_1426),
.A2(n_1315),
.B(n_1319),
.Y(n_1596)
);

O2A1O1Ixp5_ASAP7_75t_L g1597 ( 
.A1(n_1460),
.A2(n_1342),
.B(n_1473),
.C(n_1459),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1429),
.B(n_1443),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1489),
.Y(n_1599)
);

CKINVDCx20_ASAP7_75t_R g1600 ( 
.A(n_1513),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1571),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1555),
.B(n_1557),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1507),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1554),
.Y(n_1604)
);

INVxp33_ASAP7_75t_L g1605 ( 
.A(n_1504),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1488),
.B(n_1575),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1526),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1570),
.B(n_1589),
.Y(n_1608)
);

OA21x2_ASAP7_75t_L g1609 ( 
.A1(n_1498),
.A2(n_1490),
.B(n_1548),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1564),
.Y(n_1610)
);

AO21x2_ASAP7_75t_L g1611 ( 
.A1(n_1528),
.A2(n_1523),
.B(n_1490),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1496),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1496),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1555),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1488),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1502),
.B(n_1514),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1575),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1590),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1522),
.B(n_1534),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1590),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1500),
.B(n_1566),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1595),
.Y(n_1622)
);

AO21x2_ASAP7_75t_L g1623 ( 
.A1(n_1567),
.A2(n_1500),
.B(n_1562),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1595),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1506),
.B(n_1497),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1511),
.Y(n_1626)
);

INVxp33_ASAP7_75t_L g1627 ( 
.A(n_1549),
.Y(n_1627)
);

AOI21x1_ASAP7_75t_L g1628 ( 
.A1(n_1487),
.A2(n_1566),
.B(n_1486),
.Y(n_1628)
);

AO21x2_ASAP7_75t_L g1629 ( 
.A1(n_1562),
.A2(n_1519),
.B(n_1593),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1499),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1557),
.Y(n_1631)
);

INVxp33_ASAP7_75t_L g1632 ( 
.A(n_1510),
.Y(n_1632)
);

AO31x2_ASAP7_75t_L g1633 ( 
.A1(n_1494),
.A2(n_1573),
.A3(n_1586),
.B(n_1585),
.Y(n_1633)
);

AO21x2_ASAP7_75t_L g1634 ( 
.A1(n_1506),
.A2(n_1561),
.B(n_1540),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1492),
.B(n_1503),
.Y(n_1635)
);

OR2x6_ASAP7_75t_L g1636 ( 
.A(n_1546),
.B(n_1530),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1521),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1568),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1594),
.B(n_1568),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1561),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1558),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1491),
.B(n_1493),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1578),
.B(n_1582),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1558),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1584),
.B(n_1592),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1515),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1485),
.A2(n_1597),
.B(n_1508),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1505),
.Y(n_1648)
);

AOI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1495),
.A2(n_1577),
.B(n_1587),
.Y(n_1649)
);

OA21x2_ASAP7_75t_L g1650 ( 
.A1(n_1576),
.A2(n_1518),
.B(n_1572),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1577),
.A2(n_1596),
.B(n_1574),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1591),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1547),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1581),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1581),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1598),
.B(n_1583),
.Y(n_1656)
);

OA21x2_ASAP7_75t_L g1657 ( 
.A1(n_1518),
.A2(n_1579),
.B(n_1588),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1509),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1569),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1541),
.Y(n_1660)
);

AO21x2_ASAP7_75t_L g1661 ( 
.A1(n_1540),
.A2(n_1524),
.B(n_1565),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1501),
.Y(n_1662)
);

INVxp67_ASAP7_75t_SL g1663 ( 
.A(n_1527),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1601),
.B(n_1553),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1646),
.Y(n_1665)
);

NOR2x1_ASAP7_75t_L g1666 ( 
.A(n_1636),
.B(n_1634),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1656),
.B(n_1501),
.Y(n_1667)
);

INVxp67_ASAP7_75t_SL g1668 ( 
.A(n_1614),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1599),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1646),
.Y(n_1670)
);

BUFx6f_ASAP7_75t_L g1671 ( 
.A(n_1609),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1599),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1602),
.B(n_1520),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1616),
.B(n_1563),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1603),
.Y(n_1675)
);

INVxp67_ASAP7_75t_SL g1676 ( 
.A(n_1614),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1653),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1653),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1621),
.B(n_1512),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1649),
.B(n_1517),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1609),
.Y(n_1681)
);

CKINVDCx14_ASAP7_75t_R g1682 ( 
.A(n_1600),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1612),
.B(n_1613),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1601),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1653),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1604),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1654),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1612),
.B(n_1559),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1609),
.B(n_1619),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1609),
.B(n_1533),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1611),
.B(n_1608),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1604),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1611),
.B(n_1533),
.Y(n_1693)
);

NOR2x1_ASAP7_75t_L g1694 ( 
.A(n_1636),
.B(n_1537),
.Y(n_1694)
);

INVxp67_ASAP7_75t_SL g1695 ( 
.A(n_1631),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_SL g1696 ( 
.A1(n_1629),
.A2(n_1650),
.B1(n_1657),
.B2(n_1663),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1611),
.B(n_1525),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1611),
.B(n_1551),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1654),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1602),
.B(n_1536),
.Y(n_1700)
);

INVx4_ASAP7_75t_L g1701 ( 
.A(n_1636),
.Y(n_1701)
);

INVxp67_ASAP7_75t_L g1702 ( 
.A(n_1613),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1604),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1631),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1652),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1639),
.B(n_1529),
.Y(n_1706)
);

OAI33xp33_ASAP7_75t_L g1707 ( 
.A1(n_1688),
.A2(n_1625),
.A3(n_1606),
.B1(n_1624),
.B2(n_1622),
.B3(n_1615),
.Y(n_1707)
);

INVxp67_ASAP7_75t_L g1708 ( 
.A(n_1706),
.Y(n_1708)
);

NOR2x1_ASAP7_75t_SL g1709 ( 
.A(n_1674),
.B(n_1636),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1704),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_1706),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1706),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1696),
.A2(n_1650),
.B1(n_1657),
.B2(n_1629),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1664),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1696),
.A2(n_1649),
.B1(n_1651),
.B2(n_1650),
.Y(n_1715)
);

INVx4_ASAP7_75t_L g1716 ( 
.A(n_1705),
.Y(n_1716)
);

OAI322xp33_ASAP7_75t_L g1717 ( 
.A1(n_1689),
.A2(n_1651),
.A3(n_1625),
.B1(n_1663),
.B2(n_1633),
.C1(n_1650),
.C2(n_1606),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1669),
.Y(n_1718)
);

AO21x2_ASAP7_75t_L g1719 ( 
.A1(n_1693),
.A2(n_1623),
.B(n_1638),
.Y(n_1719)
);

OAI31xp33_ASAP7_75t_L g1720 ( 
.A1(n_1680),
.A2(n_1531),
.A3(n_1650),
.B(n_1690),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1680),
.A2(n_1657),
.B1(n_1647),
.B2(n_1628),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1697),
.B(n_1615),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1694),
.A2(n_1647),
.B(n_1657),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1669),
.Y(n_1724)
);

BUFx3_ASAP7_75t_L g1725 ( 
.A(n_1673),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1667),
.B(n_1662),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1669),
.Y(n_1727)
);

NAND2xp33_ASAP7_75t_R g1728 ( 
.A(n_1674),
.B(n_1657),
.Y(n_1728)
);

NAND4xp25_ASAP7_75t_L g1729 ( 
.A(n_1689),
.B(n_1607),
.C(n_1635),
.D(n_1580),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1697),
.B(n_1617),
.Y(n_1730)
);

AOI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1693),
.A2(n_1629),
.B1(n_1661),
.B2(n_1633),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1694),
.A2(n_1629),
.B(n_1636),
.Y(n_1732)
);

OAI221xp5_ASAP7_75t_SL g1733 ( 
.A1(n_1689),
.A2(n_1633),
.B1(n_1641),
.B2(n_1644),
.C(n_1630),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1704),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1667),
.B(n_1662),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1697),
.B(n_1617),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1682),
.A2(n_1628),
.B1(n_1605),
.B2(n_1627),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1667),
.B(n_1679),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1679),
.B(n_1662),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1686),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1690),
.A2(n_1661),
.B1(n_1641),
.B2(n_1644),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1668),
.B(n_1648),
.Y(n_1742)
);

NOR4xp25_ASAP7_75t_SL g1743 ( 
.A(n_1684),
.B(n_1560),
.C(n_1550),
.D(n_1556),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1689),
.A2(n_1624),
.B1(n_1622),
.B2(n_1618),
.C(n_1620),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1672),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1686),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1668),
.B(n_1618),
.Y(n_1747)
);

OR2x6_ASAP7_75t_L g1748 ( 
.A(n_1701),
.B(n_1636),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1701),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1672),
.Y(n_1750)
);

AOI31xp67_ASAP7_75t_L g1751 ( 
.A1(n_1665),
.A2(n_1678),
.A3(n_1699),
.B(n_1677),
.Y(n_1751)
);

AOI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1688),
.A2(n_1620),
.B1(n_1634),
.B2(n_1637),
.C(n_1626),
.Y(n_1752)
);

AO21x2_ASAP7_75t_L g1753 ( 
.A1(n_1690),
.A2(n_1623),
.B(n_1638),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1676),
.B(n_1648),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1692),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1664),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1674),
.A2(n_1661),
.B1(n_1634),
.B2(n_1623),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1672),
.Y(n_1758)
);

CKINVDCx20_ASAP7_75t_R g1759 ( 
.A(n_1682),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1675),
.Y(n_1760)
);

NOR4xp25_ASAP7_75t_SL g1761 ( 
.A(n_1684),
.B(n_1607),
.C(n_1640),
.D(n_1626),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1666),
.A2(n_1661),
.B1(n_1634),
.B2(n_1659),
.Y(n_1762)
);

INVx1_ASAP7_75t_SL g1763 ( 
.A(n_1673),
.Y(n_1763)
);

AO21x2_ASAP7_75t_L g1764 ( 
.A1(n_1731),
.A2(n_1610),
.B(n_1655),
.Y(n_1764)
);

AO21x2_ASAP7_75t_L g1765 ( 
.A1(n_1731),
.A2(n_1610),
.B(n_1670),
.Y(n_1765)
);

OAI21x1_ASAP7_75t_L g1766 ( 
.A1(n_1732),
.A2(n_1666),
.B(n_1670),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1722),
.B(n_1683),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1723),
.B(n_1702),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1710),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1751),
.Y(n_1770)
);

AO21x2_ASAP7_75t_L g1771 ( 
.A1(n_1713),
.A2(n_1610),
.B(n_1670),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_SL g1772 ( 
.A1(n_1715),
.A2(n_1552),
.B(n_1671),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1711),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1720),
.B(n_1694),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1718),
.Y(n_1775)
);

NOR2x1p5_ASAP7_75t_L g1776 ( 
.A(n_1729),
.B(n_1539),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1738),
.B(n_1691),
.Y(n_1777)
);

BUFx2_ASAP7_75t_L g1778 ( 
.A(n_1759),
.Y(n_1778)
);

INVx3_ASAP7_75t_L g1779 ( 
.A(n_1714),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1718),
.Y(n_1780)
);

AO21x2_ASAP7_75t_L g1781 ( 
.A1(n_1713),
.A2(n_1678),
.B(n_1677),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1724),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1724),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1738),
.B(n_1691),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1727),
.Y(n_1785)
);

NOR2x1_ASAP7_75t_L g1786 ( 
.A(n_1716),
.B(n_1684),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1720),
.B(n_1691),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1759),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1727),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1745),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1745),
.Y(n_1791)
);

AO21x1_ASAP7_75t_SL g1792 ( 
.A1(n_1742),
.A2(n_1703),
.B(n_1692),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1739),
.B(n_1679),
.Y(n_1793)
);

INVx4_ASAP7_75t_SL g1794 ( 
.A(n_1748),
.Y(n_1794)
);

NAND3xp33_ASAP7_75t_L g1795 ( 
.A(n_1721),
.B(n_1681),
.C(n_1671),
.Y(n_1795)
);

BUFx2_ASAP7_75t_L g1796 ( 
.A(n_1734),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1750),
.Y(n_1797)
);

AND2x6_ASAP7_75t_SL g1798 ( 
.A(n_1748),
.B(n_1532),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1750),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1739),
.B(n_1679),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1742),
.Y(n_1801)
);

OAI21x1_ASAP7_75t_L g1802 ( 
.A1(n_1757),
.A2(n_1687),
.B(n_1685),
.Y(n_1802)
);

NOR3xp33_ASAP7_75t_L g1803 ( 
.A(n_1717),
.B(n_1702),
.C(n_1630),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1758),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1758),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1751),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1753),
.Y(n_1807)
);

AOI21x1_ASAP7_75t_L g1808 ( 
.A1(n_1737),
.A2(n_1687),
.B(n_1685),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1744),
.B(n_1676),
.Y(n_1809)
);

NAND3xp33_ASAP7_75t_SL g1810 ( 
.A(n_1761),
.B(n_1627),
.C(n_1698),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1760),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1753),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1749),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1754),
.Y(n_1814)
);

OR2x6_ASAP7_75t_L g1815 ( 
.A(n_1748),
.B(n_1543),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1768),
.B(n_1730),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1793),
.B(n_1714),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1775),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1793),
.B(n_1714),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1803),
.B(n_1752),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1800),
.B(n_1756),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1800),
.B(n_1756),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1775),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1777),
.B(n_1756),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1801),
.B(n_1736),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1809),
.B(n_1725),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1780),
.Y(n_1827)
);

INVxp67_ASAP7_75t_L g1828 ( 
.A(n_1778),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1814),
.B(n_1754),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1767),
.B(n_1747),
.Y(n_1830)
);

INVx3_ASAP7_75t_L g1831 ( 
.A(n_1813),
.Y(n_1831)
);

AOI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1787),
.A2(n_1717),
.B1(n_1707),
.B2(n_1733),
.C(n_1762),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1769),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1777),
.B(n_1726),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1781),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1784),
.B(n_1726),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1784),
.B(n_1735),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1767),
.B(n_1763),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1796),
.B(n_1725),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1780),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1792),
.B(n_1735),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1782),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1782),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1783),
.Y(n_1844)
);

INVxp67_ASAP7_75t_L g1845 ( 
.A(n_1778),
.Y(n_1845)
);

BUFx2_ASAP7_75t_L g1846 ( 
.A(n_1798),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1792),
.B(n_1711),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1773),
.B(n_1712),
.Y(n_1848)
);

NAND3xp33_ASAP7_75t_L g1849 ( 
.A(n_1795),
.B(n_1728),
.C(n_1681),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1796),
.B(n_1683),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1774),
.B(n_1695),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1776),
.B(n_1695),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1781),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1773),
.B(n_1712),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1783),
.B(n_1673),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1788),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1776),
.B(n_1658),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1785),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1785),
.B(n_1740),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1789),
.Y(n_1860)
);

BUFx2_ASAP7_75t_L g1861 ( 
.A(n_1798),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1789),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1813),
.B(n_1716),
.Y(n_1863)
);

AOI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1772),
.A2(n_1709),
.B(n_1743),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1790),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1795),
.B(n_1658),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1790),
.B(n_1746),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1791),
.B(n_1755),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1772),
.B(n_1642),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1791),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1797),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1813),
.B(n_1716),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1847),
.B(n_1813),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1828),
.B(n_1633),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1847),
.B(n_1813),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1860),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1831),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1841),
.B(n_1813),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1835),
.Y(n_1879)
);

NAND4xp25_ASAP7_75t_L g1880 ( 
.A(n_1846),
.B(n_1786),
.C(n_1770),
.D(n_1806),
.Y(n_1880)
);

AND3x2_ASAP7_75t_L g1881 ( 
.A(n_1846),
.B(n_1660),
.C(n_1600),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1838),
.B(n_1700),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1845),
.B(n_1786),
.Y(n_1883)
);

OAI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1820),
.A2(n_1810),
.B1(n_1815),
.B2(n_1808),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1832),
.A2(n_1771),
.B1(n_1765),
.B2(n_1781),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1838),
.B(n_1700),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1835),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1830),
.B(n_1700),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1830),
.B(n_1797),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1842),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1861),
.A2(n_1849),
.B1(n_1869),
.B2(n_1851),
.Y(n_1891)
);

HB1xp67_ASAP7_75t_L g1892 ( 
.A(n_1833),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1829),
.B(n_1799),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1861),
.B(n_1605),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1841),
.B(n_1779),
.Y(n_1895)
);

INVx1_ASAP7_75t_SL g1896 ( 
.A(n_1839),
.Y(n_1896)
);

INVx1_ASAP7_75t_SL g1897 ( 
.A(n_1848),
.Y(n_1897)
);

BUFx2_ASAP7_75t_SL g1898 ( 
.A(n_1863),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1848),
.B(n_1779),
.Y(n_1899)
);

AND2x2_ASAP7_75t_SL g1900 ( 
.A(n_1863),
.B(n_1701),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1854),
.B(n_1872),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1854),
.B(n_1779),
.Y(n_1902)
);

INVx2_ASAP7_75t_SL g1903 ( 
.A(n_1872),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1829),
.B(n_1799),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1856),
.B(n_1633),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1816),
.B(n_1804),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_SL g1907 ( 
.A1(n_1826),
.A2(n_1771),
.B1(n_1765),
.B2(n_1781),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1816),
.B(n_1804),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1853),
.Y(n_1909)
);

OAI21xp33_ASAP7_75t_L g1910 ( 
.A1(n_1866),
.A2(n_1852),
.B(n_1857),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1850),
.B(n_1633),
.Y(n_1911)
);

INVx1_ASAP7_75t_SL g1912 ( 
.A(n_1850),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1825),
.B(n_1633),
.Y(n_1913)
);

NOR4xp25_ASAP7_75t_L g1914 ( 
.A(n_1831),
.B(n_1770),
.C(n_1806),
.D(n_1853),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1825),
.B(n_1642),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1901),
.B(n_1834),
.Y(n_1916)
);

CKINVDCx16_ASAP7_75t_R g1917 ( 
.A(n_1894),
.Y(n_1917)
);

NOR2x1_ASAP7_75t_L g1918 ( 
.A(n_1894),
.B(n_1831),
.Y(n_1918)
);

INVxp67_ASAP7_75t_L g1919 ( 
.A(n_1892),
.Y(n_1919)
);

AO21x1_ASAP7_75t_SL g1920 ( 
.A1(n_1892),
.A2(n_1823),
.B(n_1818),
.Y(n_1920)
);

AOI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1885),
.A2(n_1771),
.B1(n_1765),
.B2(n_1764),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1912),
.B(n_1834),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1890),
.Y(n_1923)
);

NAND2xp33_ASAP7_75t_L g1924 ( 
.A(n_1897),
.B(n_1864),
.Y(n_1924)
);

CKINVDCx16_ASAP7_75t_R g1925 ( 
.A(n_1898),
.Y(n_1925)
);

INVx1_ASAP7_75t_SL g1926 ( 
.A(n_1881),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1876),
.Y(n_1927)
);

OAI221xp5_ASAP7_75t_L g1928 ( 
.A1(n_1907),
.A2(n_1808),
.B1(n_1770),
.B2(n_1806),
.C(n_1741),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1901),
.B(n_1878),
.Y(n_1929)
);

HB1xp67_ASAP7_75t_L g1930 ( 
.A(n_1896),
.Y(n_1930)
);

INVx1_ASAP7_75t_SL g1931 ( 
.A(n_1903),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1903),
.B(n_1836),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1906),
.Y(n_1933)
);

INVx4_ASAP7_75t_L g1934 ( 
.A(n_1877),
.Y(n_1934)
);

INVxp67_ASAP7_75t_SL g1935 ( 
.A(n_1884),
.Y(n_1935)
);

OR2x2_ASAP7_75t_L g1936 ( 
.A(n_1905),
.B(n_1855),
.Y(n_1936)
);

INVx1_ASAP7_75t_SL g1937 ( 
.A(n_1873),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1908),
.Y(n_1938)
);

OAI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1884),
.A2(n_1802),
.B(n_1766),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1874),
.B(n_1836),
.Y(n_1940)
);

INVx2_ASAP7_75t_SL g1941 ( 
.A(n_1900),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1893),
.Y(n_1942)
);

NAND2xp33_ASAP7_75t_L g1943 ( 
.A(n_1891),
.B(n_1855),
.Y(n_1943)
);

INVx1_ASAP7_75t_SL g1944 ( 
.A(n_1873),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1882),
.B(n_1859),
.Y(n_1945)
);

AOI22xp33_ASAP7_75t_SL g1946 ( 
.A1(n_1935),
.A2(n_1917),
.B1(n_1943),
.B2(n_1930),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1935),
.A2(n_1880),
.B(n_1911),
.Y(n_1947)
);

NAND3xp33_ASAP7_75t_L g1948 ( 
.A(n_1943),
.B(n_1913),
.C(n_1914),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1929),
.Y(n_1949)
);

O2A1O1Ixp33_ASAP7_75t_L g1950 ( 
.A1(n_1930),
.A2(n_1910),
.B(n_1883),
.C(n_1904),
.Y(n_1950)
);

INVx1_ASAP7_75t_SL g1951 ( 
.A(n_1926),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1923),
.Y(n_1952)
);

AOI222xp33_ASAP7_75t_L g1953 ( 
.A1(n_1928),
.A2(n_1812),
.B1(n_1807),
.B2(n_1909),
.C1(n_1887),
.C2(n_1879),
.Y(n_1953)
);

OA222x2_ASAP7_75t_L g1954 ( 
.A1(n_1919),
.A2(n_1886),
.B1(n_1877),
.B2(n_1815),
.C1(n_1748),
.C2(n_1889),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1925),
.A2(n_1900),
.B1(n_1888),
.B2(n_1915),
.Y(n_1955)
);

OAI211xp5_ASAP7_75t_L g1956 ( 
.A1(n_1918),
.A2(n_1875),
.B(n_1878),
.C(n_1895),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1931),
.B(n_1883),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1916),
.B(n_1883),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1932),
.B(n_1875),
.Y(n_1959)
);

INVxp67_ASAP7_75t_L g1960 ( 
.A(n_1920),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1932),
.Y(n_1961)
);

OR2x2_ASAP7_75t_L g1962 ( 
.A(n_1922),
.B(n_1859),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1919),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1932),
.Y(n_1964)
);

AOI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1921),
.A2(n_1771),
.B1(n_1765),
.B2(n_1764),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1924),
.A2(n_1939),
.B1(n_1933),
.B2(n_1938),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1934),
.B(n_1877),
.Y(n_1967)
);

OAI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1924),
.A2(n_1895),
.B(n_1802),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1961),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1961),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1959),
.B(n_1937),
.Y(n_1971)
);

INVx4_ASAP7_75t_L g1972 ( 
.A(n_1964),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1949),
.Y(n_1973)
);

INVx1_ASAP7_75t_SL g1974 ( 
.A(n_1951),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1946),
.B(n_1944),
.Y(n_1975)
);

INVx2_ASAP7_75t_SL g1976 ( 
.A(n_1967),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1946),
.B(n_1942),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1960),
.B(n_1941),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1966),
.B(n_1934),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1947),
.B(n_1927),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1963),
.B(n_1945),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1962),
.B(n_1940),
.Y(n_1982)
);

NOR2x1_ASAP7_75t_L g1983 ( 
.A(n_1948),
.B(n_1544),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1952),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1957),
.Y(n_1985)
);

O2A1O1Ixp33_ASAP7_75t_L g1986 ( 
.A1(n_1979),
.A2(n_1950),
.B(n_1966),
.C(n_1960),
.Y(n_1986)
);

OAI211xp5_ASAP7_75t_SL g1987 ( 
.A1(n_1975),
.A2(n_1968),
.B(n_1967),
.C(n_1958),
.Y(n_1987)
);

OAI221xp5_ASAP7_75t_L g1988 ( 
.A1(n_1977),
.A2(n_1965),
.B1(n_1953),
.B2(n_1955),
.C(n_1956),
.Y(n_1988)
);

AOI211xp5_ASAP7_75t_L g1989 ( 
.A1(n_1979),
.A2(n_1936),
.B(n_1954),
.C(n_1899),
.Y(n_1989)
);

AOI21xp33_ASAP7_75t_SL g1990 ( 
.A1(n_1976),
.A2(n_1902),
.B(n_1899),
.Y(n_1990)
);

AOI221xp5_ASAP7_75t_L g1991 ( 
.A1(n_1980),
.A2(n_1812),
.B1(n_1807),
.B2(n_1887),
.C(n_1879),
.Y(n_1991)
);

AOI22xp33_ASAP7_75t_SL g1992 ( 
.A1(n_1974),
.A2(n_1807),
.B1(n_1812),
.B2(n_1764),
.Y(n_1992)
);

AOI221xp5_ASAP7_75t_L g1993 ( 
.A1(n_1985),
.A2(n_1909),
.B1(n_1764),
.B2(n_1671),
.C(n_1681),
.Y(n_1993)
);

NAND2xp33_ASAP7_75t_R g1994 ( 
.A(n_1971),
.B(n_1743),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1976),
.B(n_1902),
.Y(n_1995)
);

AOI211xp5_ASAP7_75t_L g1996 ( 
.A1(n_1978),
.A2(n_1681),
.B(n_1671),
.C(n_1842),
.Y(n_1996)
);

NAND4xp25_ASAP7_75t_SL g1997 ( 
.A(n_1981),
.B(n_1824),
.C(n_1819),
.D(n_1821),
.Y(n_1997)
);

AOI221xp5_ASAP7_75t_L g1998 ( 
.A1(n_1984),
.A2(n_1681),
.B1(n_1671),
.B2(n_1844),
.C(n_1719),
.Y(n_1998)
);

OAI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1973),
.A2(n_1982),
.B1(n_1983),
.B2(n_1969),
.Y(n_1999)
);

OAI211xp5_ASAP7_75t_SL g2000 ( 
.A1(n_1970),
.A2(n_1844),
.B(n_1870),
.C(n_1871),
.Y(n_2000)
);

OAI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1989),
.A2(n_1973),
.B1(n_1972),
.B2(n_1978),
.Y(n_2001)
);

INVx2_ASAP7_75t_SL g2002 ( 
.A(n_1995),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1999),
.Y(n_2003)
);

AOI221xp5_ASAP7_75t_L g2004 ( 
.A1(n_1988),
.A2(n_1972),
.B1(n_1671),
.B2(n_1681),
.C(n_1865),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1994),
.Y(n_2005)
);

AOI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1987),
.A2(n_1972),
.B1(n_1535),
.B2(n_1753),
.Y(n_2006)
);

OAI221xp5_ASAP7_75t_L g2007 ( 
.A1(n_1986),
.A2(n_1516),
.B1(n_1862),
.B2(n_1858),
.C(n_1843),
.Y(n_2007)
);

AOI211xp5_ASAP7_75t_L g2008 ( 
.A1(n_1990),
.A2(n_1671),
.B(n_1681),
.C(n_1840),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_2002),
.B(n_1837),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_2003),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_2007),
.Y(n_2011)
);

AOI32xp33_ASAP7_75t_L g2012 ( 
.A1(n_2001),
.A2(n_2000),
.A3(n_1992),
.B1(n_1996),
.B2(n_1998),
.Y(n_2012)
);

NOR2x1_ASAP7_75t_L g2013 ( 
.A(n_2005),
.B(n_1997),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_2006),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_2004),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_2008),
.B(n_1867),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_2009),
.B(n_1993),
.Y(n_2017)
);

OAI21xp33_ASAP7_75t_SL g2018 ( 
.A1(n_2012),
.A2(n_1991),
.B(n_1827),
.Y(n_2018)
);

NOR2x1_ASAP7_75t_L g2019 ( 
.A(n_2013),
.B(n_1867),
.Y(n_2019)
);

HB1xp67_ASAP7_75t_L g2020 ( 
.A(n_2010),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_2015),
.B(n_1868),
.Y(n_2021)
);

AOI322xp5_ASAP7_75t_L g2022 ( 
.A1(n_2014),
.A2(n_2011),
.A3(n_2016),
.B1(n_1698),
.B2(n_1837),
.C1(n_1671),
.C2(n_1681),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_R g2023 ( 
.A(n_2010),
.B(n_1779),
.Y(n_2023)
);

INVxp67_ASAP7_75t_L g2024 ( 
.A(n_2020),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_L g2025 ( 
.A(n_2018),
.B(n_1868),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_2019),
.B(n_2021),
.Y(n_2026)
);

AND2x4_ASAP7_75t_L g2027 ( 
.A(n_2017),
.B(n_1817),
.Y(n_2027)
);

OAI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_2024),
.A2(n_2022),
.B1(n_2023),
.B2(n_1824),
.Y(n_2028)
);

OAI221xp5_ASAP7_75t_SL g2029 ( 
.A1(n_2028),
.A2(n_2026),
.B1(n_2025),
.B2(n_2027),
.C(n_1815),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_2029),
.B(n_1822),
.Y(n_2030)
);

CKINVDCx16_ASAP7_75t_R g2031 ( 
.A(n_2029),
.Y(n_2031)
);

OAI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_2031),
.A2(n_1822),
.B1(n_1821),
.B2(n_1819),
.Y(n_2032)
);

NAND2x1p5_ASAP7_75t_L g2033 ( 
.A(n_2030),
.B(n_1538),
.Y(n_2033)
);

HB1xp67_ASAP7_75t_L g2034 ( 
.A(n_2033),
.Y(n_2034)
);

OAI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_2032),
.A2(n_1817),
.B1(n_1811),
.B2(n_1805),
.Y(n_2035)
);

AOI22xp5_ASAP7_75t_SL g2036 ( 
.A1(n_2034),
.A2(n_1708),
.B1(n_1645),
.B2(n_1643),
.Y(n_2036)
);

OAI321xp33_ASAP7_75t_L g2037 ( 
.A1(n_2036),
.A2(n_2035),
.A3(n_1815),
.B1(n_1805),
.B2(n_1811),
.C(n_1749),
.Y(n_2037)
);

NOR2x1_ASAP7_75t_SL g2038 ( 
.A(n_2037),
.B(n_1538),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2038),
.Y(n_2039)
);

AOI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_2039),
.A2(n_1794),
.B1(n_1545),
.B2(n_1538),
.Y(n_2040)
);

AOI211xp5_ASAP7_75t_L g2041 ( 
.A1(n_2040),
.A2(n_1542),
.B(n_1632),
.C(n_1749),
.Y(n_2041)
);


endmodule