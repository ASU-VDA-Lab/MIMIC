module fake_jpeg_22289_n_246 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_246);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_246;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_19),
.Y(n_65)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_24),
.B1(n_33),
.B2(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_29),
.B1(n_33),
.B2(n_22),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_56),
.B1(n_69),
.B2(n_39),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_47),
.A2(n_52),
.B(n_61),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_59),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_33),
.B1(n_29),
.B2(n_30),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_43),
.B1(n_37),
.B2(n_38),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_57),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_30),
.B1(n_31),
.B2(n_17),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_31),
.B1(n_19),
.B2(n_28),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_39),
.B1(n_43),
.B2(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_35),
.B(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_67),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_65),
.B(n_36),
.Y(n_92)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_32),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_32),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_36),
.A2(n_19),
.B1(n_17),
.B2(n_34),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_79),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_37),
.B1(n_43),
.B2(n_45),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_80),
.B1(n_81),
.B2(n_89),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_34),
.B1(n_17),
.B2(n_28),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_37),
.B1(n_43),
.B2(n_45),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_47),
.B1(n_52),
.B2(n_60),
.Y(n_105)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_85),
.Y(n_101)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_94),
.Y(n_112)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_36),
.B1(n_41),
.B2(n_28),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_34),
.B1(n_31),
.B2(n_26),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_48),
.B(n_79),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_25),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_50),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_55),
.B(n_60),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_27),
.B1(n_25),
.B2(n_23),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_89),
.B1(n_81),
.B2(n_74),
.Y(n_110)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_51),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_111),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_68),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_104),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_93),
.B1(n_62),
.B2(n_84),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_65),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_86),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_55),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_78),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_110),
.A2(n_113),
.B1(n_97),
.B2(n_61),
.Y(n_129)
);

CKINVDCx12_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

AO21x2_ASAP7_75t_SL g113 ( 
.A1(n_80),
.A2(n_69),
.B(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_59),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_117),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g116 ( 
.A(n_92),
.B(n_69),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_118),
.B(n_123),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_65),
.B(n_50),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_122),
.A2(n_84),
.B1(n_97),
.B2(n_51),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_50),
.Y(n_123)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_94),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_72),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_139),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_136),
.B1(n_154),
.B2(n_100),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_113),
.B(n_122),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_110),
.B1(n_113),
.B2(n_103),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_51),
.B1(n_82),
.B2(n_62),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_73),
.C(n_48),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_102),
.C(n_40),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_64),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_113),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_20),
.B(n_18),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_71),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_112),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_125),
.B(n_126),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_71),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_149),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_77),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_104),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_99),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_115),
.B(n_83),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_113),
.A2(n_106),
.B1(n_110),
.B2(n_116),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_155),
.A2(n_99),
.B(n_113),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_131),
.B(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_156),
.B(n_164),
.Y(n_191)
);

AO21x1_ASAP7_75t_L g194 ( 
.A1(n_157),
.A2(n_151),
.B(n_107),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_158),
.A2(n_168),
.B(n_134),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_165),
.Y(n_187)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_180),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_162),
.A2(n_173),
.B1(n_135),
.B2(n_130),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_136),
.B(n_141),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_122),
.B(n_111),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_120),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_169),
.B(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_172),
.C(n_176),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_102),
.C(n_121),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_133),
.B1(n_137),
.B2(n_155),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_40),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_179),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_40),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_130),
.B(n_166),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_121),
.B(n_107),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_121),
.C(n_40),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_199),
.B1(n_179),
.B2(n_175),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_189),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_161),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_188),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_134),
.B(n_149),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_163),
.B(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_88),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_124),
.C(n_18),
.Y(n_208)
);

AOI21x1_ASAP7_75t_L g197 ( 
.A1(n_158),
.A2(n_18),
.B(n_104),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_162),
.A2(n_144),
.B1(n_58),
.B2(n_88),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_185),
.B(n_160),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_205),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_165),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_207),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_206),
.A2(n_23),
.B(n_16),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_18),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_209),
.C(n_183),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_119),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_213),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_183),
.C(n_195),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_210),
.A2(n_197),
.B1(n_193),
.B2(n_194),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_204),
.A2(n_191),
.B1(n_186),
.B2(n_195),
.Y(n_217)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_23),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_222),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_220),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_201),
.A2(n_9),
.B(n_15),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_27),
.C(n_16),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_205),
.Y(n_223)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_207),
.B(n_1),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_8),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_221),
.C(n_214),
.Y(n_232)
);

AND2x6_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_216),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_231),
.A2(n_7),
.B(n_8),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_233),
.C(n_234),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_225),
.C(n_223),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_3),
.C(n_4),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_228),
.B(n_226),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_233),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_239),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_234),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_235),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_237),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_242),
.A2(n_13),
.B(n_241),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_243),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_244),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);


endmodule