module fake_jpeg_1799_n_378 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_378);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_378;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx9p33_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_11),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_58),
.B(n_62),
.C(n_78),
.Y(n_141)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_32),
.A2(n_9),
.B(n_14),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_73),
.Y(n_116)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_9),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_18),
.Y(n_63)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_63),
.Y(n_150)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_67),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_6),
.B1(n_12),
.B2(n_13),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_68),
.A2(n_29),
.B1(n_37),
.B2(n_50),
.Y(n_115)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_19),
.B(n_12),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_79),
.Y(n_167)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_19),
.B(n_13),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_86),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_83),
.Y(n_142)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_84),
.B(n_85),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_91),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_88),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_89),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

BUFx24_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

BUFx4f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_101),
.B1(n_107),
.B2(n_34),
.Y(n_118)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

NAND2x1_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_100),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_96),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g95 ( 
.A(n_33),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_95),
.B(n_99),
.Y(n_170)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_98),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_21),
.B(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_103),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_53),
.Y(n_117)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_109),
.Y(n_139)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_21),
.B(n_16),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_94),
.A2(n_53),
.B1(n_54),
.B2(n_52),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_114),
.A2(n_142),
.B1(n_152),
.B2(n_155),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_115),
.B(n_117),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_118),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_78),
.A2(n_53),
.B1(n_52),
.B2(n_51),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_121),
.A2(n_138),
.B1(n_144),
.B2(n_149),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_62),
.B(n_50),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_123),
.B(n_136),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_46),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_65),
.A2(n_39),
.B1(n_34),
.B2(n_51),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_70),
.A2(n_39),
.B1(n_47),
.B2(n_38),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_28),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_146),
.B(n_162),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_81),
.B(n_46),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_148),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_37),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_92),
.A2(n_29),
.B1(n_38),
.B2(n_31),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_82),
.A2(n_26),
.B1(n_31),
.B2(n_28),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_152),
.A2(n_159),
.B1(n_161),
.B2(n_165),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_74),
.B(n_25),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_160),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_88),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_76),
.B(n_27),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_95),
.A2(n_47),
.B1(n_1),
.B2(n_3),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_67),
.B(n_0),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_63),
.B(n_0),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_164),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_61),
.B(n_1),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_77),
.A2(n_3),
.B1(n_64),
.B2(n_103),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_89),
.A2(n_104),
.B1(n_90),
.B2(n_100),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_57),
.B1(n_71),
.B2(n_117),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_116),
.A2(n_91),
.B1(n_80),
.B2(n_102),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_171),
.A2(n_189),
.B1(n_174),
.B2(n_187),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_172),
.A2(n_179),
.B1(n_181),
.B2(n_211),
.Y(n_235)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVxp67_ASAP7_75t_SL g240 ( 
.A(n_173),
.Y(n_240)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_112),
.Y(n_175)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_175),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_123),
.B(n_147),
.C(n_136),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g223 ( 
.A1(n_176),
.A2(n_151),
.B(n_132),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_177),
.B(n_178),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_131),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_160),
.B1(n_166),
.B2(n_159),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_129),
.A2(n_168),
.B1(n_154),
.B2(n_167),
.Y(n_181)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_170),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_185),
.B(n_190),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_203),
.Y(n_232)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_140),
.A2(n_139),
.B1(n_130),
.B2(n_127),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_115),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_192),
.Y(n_238)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_195),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_157),
.Y(n_196)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_198),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_119),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_210),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_200),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_115),
.B(n_133),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_201),
.B(n_208),
.Y(n_244)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_137),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_202),
.Y(n_249)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_142),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_206),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_155),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_126),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_209),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_115),
.B(n_157),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_142),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_119),
.B(n_155),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_134),
.A2(n_145),
.B1(n_113),
.B2(n_120),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_134),
.B(n_122),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_209),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_156),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_216),
.Y(n_226)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_151),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_113),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_218),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_112),
.B(n_120),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_L g219 ( 
.A1(n_125),
.A2(n_143),
.B1(n_156),
.B2(n_132),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_219),
.A2(n_172),
.B1(n_211),
.B2(n_179),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_231),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_137),
.C(n_125),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_236),
.C(n_239),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_143),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_193),
.C(n_182),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_215),
.B(n_199),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_L g271 ( 
.A1(n_237),
.A2(n_175),
.B(n_221),
.C(n_248),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_182),
.C(n_180),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_248),
.B1(n_250),
.B2(n_183),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_254),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_180),
.A2(n_186),
.B1(n_215),
.B2(n_184),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_180),
.A2(n_213),
.B1(n_197),
.B2(n_212),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_196),
.B(n_194),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_253),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_176),
.B(n_196),
.Y(n_254)
);

AND2x2_ASAP7_75t_SL g255 ( 
.A(n_188),
.B(n_217),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_251),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_252),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_278),
.Y(n_292)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_234),
.Y(n_259)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

A2O1A1O1Ixp25_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_207),
.B(n_203),
.C(n_219),
.D(n_195),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_260),
.A2(n_261),
.B(n_263),
.Y(n_287)
);

NAND2xp67_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_237),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_230),
.A2(n_200),
.B1(n_198),
.B2(n_202),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_264),
.A2(n_269),
.B1(n_270),
.B2(n_273),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_175),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_274),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_250),
.A2(n_221),
.B1(n_232),
.B2(n_254),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_230),
.A2(n_244),
.B1(n_232),
.B2(n_253),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_249),
.B(n_220),
.Y(n_291)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_232),
.A2(n_228),
.B1(n_247),
.B2(n_222),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_227),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_245),
.A2(n_235),
.B1(n_251),
.B2(n_226),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_275),
.A2(n_281),
.B1(n_241),
.B2(n_256),
.Y(n_297)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_277),
.B(n_285),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_225),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_251),
.Y(n_279)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_242),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_280),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_235),
.A2(n_256),
.B1(n_249),
.B2(n_234),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_242),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_282),
.B(n_284),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_238),
.B(n_255),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_224),
.C(n_246),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_255),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_220),
.B(n_238),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_291),
.A2(n_284),
.B(n_268),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_264),
.B1(n_269),
.B2(n_271),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_295),
.A2(n_268),
.B1(n_281),
.B2(n_265),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_258),
.B(n_241),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_300),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_258),
.B(n_246),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_306),
.C(n_274),
.Y(n_315)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_304),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_280),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_233),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_267),
.B(n_224),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_272),
.Y(n_307)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_307),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_292),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_313),
.Y(n_327)
);

NAND2x1_ASAP7_75t_SL g328 ( 
.A(n_309),
.B(n_290),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_311),
.A2(n_319),
.B1(n_321),
.B2(n_301),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_300),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_291),
.A2(n_287),
.B(n_295),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_318),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_315),
.B(n_322),
.C(n_302),
.Y(n_335)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_316),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_288),
.A2(n_267),
.B1(n_268),
.B2(n_263),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_303),
.B(n_257),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_324),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_297),
.A2(n_266),
.B1(n_261),
.B2(n_283),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_277),
.C(n_279),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_293),
.Y(n_323)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_323),
.Y(n_337)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_296),
.Y(n_325)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_325),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_313),
.A2(n_288),
.B1(n_299),
.B2(n_287),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_326),
.A2(n_316),
.B1(n_323),
.B2(n_317),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_328),
.A2(n_309),
.B(n_314),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_299),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_334),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_330),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_298),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_331),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_290),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_335),
.B(n_298),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_276),
.C(n_294),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_321),
.C(n_319),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_329),
.B(n_322),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_328),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_345),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_335),
.B(n_320),
.C(n_318),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_348),
.C(n_333),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_347),
.B(n_349),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_311),
.C(n_310),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_327),
.B(n_305),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_333),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_340),
.A2(n_326),
.B1(n_332),
.B2(n_336),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_357),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_339),
.B(n_334),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_354),
.B(n_356),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_355),
.A2(n_358),
.B(n_350),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_348),
.B(n_325),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_286),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_359),
.B(n_342),
.C(n_343),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_362),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_351),
.A2(n_359),
.B(n_353),
.Y(n_364)
);

A2O1A1Ixp33_ASAP7_75t_L g369 ( 
.A1(n_364),
.A2(n_355),
.B(n_286),
.C(n_312),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_346),
.C(n_333),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_358),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_366),
.B(n_368),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_363),
.A2(n_341),
.B1(n_337),
.B2(n_324),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_369),
.B(n_312),
.C(n_317),
.Y(n_372)
);

AO21x1_ASAP7_75t_L g370 ( 
.A1(n_367),
.A2(n_360),
.B(n_294),
.Y(n_370)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_370),
.Y(n_373)
);

A2O1A1Ixp33_ASAP7_75t_L g374 ( 
.A1(n_372),
.A2(n_366),
.B(n_307),
.C(n_260),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_374),
.B(n_373),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_375),
.A2(n_376),
.B(n_289),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_373),
.B(n_371),
.C(n_289),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_259),
.Y(n_378)
);


endmodule