module fake_jpeg_19742_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_46),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_29),
.B1(n_35),
.B2(n_23),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_50),
.B1(n_23),
.B2(n_16),
.Y(n_78)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_29),
.B1(n_35),
.B2(n_23),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_53),
.Y(n_70)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_57),
.Y(n_71)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_22),
.Y(n_75)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_67),
.Y(n_128)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_46),
.B1(n_29),
.B2(n_35),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_69),
.A2(n_89),
.B1(n_95),
.B2(n_30),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_45),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_83),
.Y(n_114)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_75),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_79),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_78),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_13),
.B(n_14),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_80),
.A2(n_94),
.B(n_106),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_17),
.B(n_20),
.C(n_34),
.Y(n_81)
);

OAI32xp33_ASAP7_75t_L g129 ( 
.A1(n_81),
.A2(n_98),
.A3(n_99),
.B1(n_101),
.B2(n_20),
.Y(n_129)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_26),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_53),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_33),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_86),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_40),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_19),
.B1(n_16),
.B2(n_26),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_32),
.B(n_34),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_88),
.A2(n_20),
.B(n_18),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_19),
.B1(n_16),
.B2(n_38),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_91),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_19),
.B1(n_16),
.B2(n_32),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_57),
.B(n_17),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_51),
.A2(n_27),
.B1(n_34),
.B2(n_31),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_52),
.A2(n_40),
.B1(n_27),
.B2(n_31),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_44),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_31),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_30),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_60),
.A2(n_30),
.B1(n_27),
.B2(n_18),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_64),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_107),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_109),
.A2(n_24),
.B1(n_25),
.B2(n_105),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_24),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_93),
.C(n_71),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_24),
.B1(n_105),
.B2(n_25),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_25),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_132),
.B(n_133),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_72),
.B(n_18),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_75),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_R g163 ( 
.A(n_129),
.B(n_77),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_88),
.A2(n_0),
.B(n_1),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_85),
.A2(n_24),
.B1(n_25),
.B2(n_15),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_134),
.A2(n_99),
.B1(n_101),
.B2(n_84),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_25),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_70),
.B(n_74),
.Y(n_147)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_139),
.A2(n_148),
.B1(n_162),
.B2(n_117),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_154),
.Y(n_170)
);

BUFx4f_ASAP7_75t_SL g142 ( 
.A(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_81),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_152),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_144),
.A2(n_149),
.B(n_151),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_145),
.A2(n_166),
.B1(n_168),
.B2(n_109),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_150),
.Y(n_179)
);

NAND2xp33_ASAP7_75t_SL g183 ( 
.A(n_147),
.B(n_163),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_96),
.B1(n_90),
.B2(n_76),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_70),
.B(n_79),
.Y(n_149)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_77),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_129),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_158),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_131),
.A2(n_95),
.B(n_107),
.C(n_67),
.Y(n_157)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_21),
.B1(n_3),
.B2(n_4),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_122),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_104),
.B(n_68),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_159),
.A2(n_133),
.B(n_114),
.Y(n_173)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_111),
.B(n_73),
.C(n_102),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_105),
.C(n_25),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_90),
.B1(n_97),
.B2(n_100),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_82),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_164),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_109),
.B(n_136),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_116),
.A2(n_67),
.B1(n_105),
.B2(n_24),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_122),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_1),
.Y(n_199)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_173),
.A2(n_202),
.B(n_151),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_152),
.A2(n_114),
.B1(n_134),
.B2(n_135),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_174),
.A2(n_188),
.B1(n_191),
.B2(n_198),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_155),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_2),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_157),
.A2(n_128),
.B1(n_115),
.B2(n_126),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_182),
.B1(n_187),
.B2(n_194),
.Y(n_214)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_125),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_200),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_157),
.A2(n_126),
.B1(n_113),
.B2(n_119),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_189),
.A2(n_150),
.B1(n_156),
.B2(n_169),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_157),
.A2(n_120),
.B1(n_119),
.B2(n_118),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_120),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_197),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_166),
.A2(n_136),
.B1(n_118),
.B2(n_117),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_121),
.B1(n_105),
.B2(n_14),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_139),
.B1(n_14),
.B2(n_13),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_165),
.C(n_147),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_1),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_163),
.A2(n_24),
.B1(n_21),
.B2(n_3),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_144),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_140),
.B(n_21),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_153),
.A2(n_159),
.B1(n_149),
.B2(n_141),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_12),
.B1(n_7),
.B2(n_8),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_181),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_205),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_176),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_208),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_207),
.B(n_212),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_176),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_210),
.C(n_220),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_154),
.C(n_141),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_151),
.Y(n_211)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_167),
.B(n_158),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_213),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_184),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_216),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_196),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_192),
.A2(n_201),
.B(n_188),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_145),
.C(n_142),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_224),
.B1(n_174),
.B2(n_198),
.Y(n_237)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_223),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_13),
.B1(n_4),
.B2(n_5),
.Y(n_224)
);

NOR2x1_ASAP7_75t_R g226 ( 
.A(n_183),
.B(n_2),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_202),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_2),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_227),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_178),
.B(n_4),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_229),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_5),
.C(n_6),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_230),
.B(n_197),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_231),
.A2(n_187),
.B1(n_173),
.B2(n_194),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_243),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_237),
.A2(n_250),
.B1(n_231),
.B2(n_228),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_240),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_186),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_210),
.B(n_200),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_249),
.C(n_251),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_215),
.B(n_189),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_190),
.C(n_171),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_179),
.C(n_185),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_217),
.C(n_206),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_256),
.A2(n_269),
.B1(n_245),
.B2(n_254),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_214),
.B1(n_227),
.B2(n_211),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_262),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_241),
.B(n_207),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_258),
.B(n_268),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_203),
.Y(n_260)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_242),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_267),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_205),
.Y(n_265)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_270),
.C(n_273),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_216),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_225),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_219),
.C(n_204),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_274),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_204),
.C(n_218),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_208),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_243),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_283),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_232),
.C(n_246),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_285),
.C(n_288),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_249),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_232),
.C(n_234),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_260),
.A2(n_245),
.B(n_247),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_263),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_287),
.A2(n_257),
.B1(n_250),
.B2(n_226),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_225),
.C(n_218),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_265),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_175),
.C(n_239),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_175),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_269),
.B(n_272),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_291),
.A2(n_297),
.B(n_303),
.Y(n_312)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_292),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_255),
.B1(n_281),
.B2(n_282),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_301),
.B1(n_302),
.B2(n_289),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_296),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_277),
.A2(n_259),
.B(n_267),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_276),
.A2(n_259),
.B(n_266),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_288),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_300),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_276),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_290),
.C(n_280),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_309),
.C(n_311),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

XOR2x2_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_285),
.Y(n_308)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_278),
.C(n_283),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_222),
.C(n_212),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_291),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_313),
.B(n_314),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_299),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_235),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_304),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_308),
.B(n_312),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_322),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_315),
.B(n_305),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_318),
.B(n_317),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_321),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_325),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_323),
.B(n_316),
.Y(n_327)
);

AOI21xp33_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_309),
.B(n_202),
.Y(n_328)
);

AOI21x1_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_12),
.B(n_7),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_330)
);


endmodule