module fake_jpeg_18812_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_40),
.Y(n_69)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_20),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_18),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_25),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_45),
.A2(n_19),
.B1(n_16),
.B2(n_22),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_22),
.B1(n_25),
.B2(n_32),
.Y(n_90)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_22),
.B1(n_20),
.B2(n_27),
.Y(n_54)
);

AO22x2_ASAP7_75t_L g100 ( 
.A1(n_54),
.A2(n_20),
.B1(n_27),
.B2(n_21),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_35),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_56),
.A2(n_27),
.B1(n_20),
.B2(n_21),
.Y(n_98)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_29),
.Y(n_84)
);

NAND2x1_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_27),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_21),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_30),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_61),
.B(n_65),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_20),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_30),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g85 ( 
.A(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_18),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_72),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_44),
.B1(n_38),
.B2(n_45),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_73),
.A2(n_75),
.B1(n_90),
.B2(n_100),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_76),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_69),
.B1(n_38),
.B2(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_91),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_79),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_39),
.B1(n_54),
.B2(n_70),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_82),
.A2(n_64),
.B1(n_66),
.B2(n_70),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_88),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_29),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_89),
.B(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_63),
.B(n_32),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_98),
.B(n_10),
.Y(n_132)
);

INVxp67_ASAP7_75t_SL g94 ( 
.A(n_67),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_35),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_66),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_63),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_56),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_26),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_51),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_50),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_23),
.B1(n_24),
.B2(n_57),
.Y(n_124)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_124),
.B1(n_130),
.B2(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_123),
.B(n_109),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_27),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_86),
.C(n_81),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_79),
.A2(n_51),
.B1(n_55),
.B2(n_34),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_82),
.A2(n_55),
.B1(n_31),
.B2(n_33),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_82),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_80),
.A2(n_34),
.B1(n_33),
.B2(n_28),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_78),
.A2(n_0),
.B(n_1),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_142),
.A2(n_126),
.B1(n_127),
.B2(n_124),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_78),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_75),
.C(n_96),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_145),
.B(n_163),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_82),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_100),
.B1(n_110),
.B2(n_73),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_147),
.A2(n_162),
.B1(n_168),
.B2(n_135),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_100),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_148),
.B(n_149),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_113),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_100),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_130),
.B(n_139),
.C(n_140),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_157),
.B(n_165),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_98),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_120),
.B(n_7),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_160),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_95),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_139),
.A2(n_111),
.B1(n_109),
.B2(n_103),
.Y(n_162)
);

MAJx3_ASAP7_75t_L g164 ( 
.A(n_112),
.B(n_102),
.C(n_81),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_116),
.B(n_126),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_139),
.A2(n_104),
.B(n_87),
.C(n_107),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_112),
.B(n_87),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_129),
.B(n_134),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_77),
.B1(n_34),
.B2(n_33),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_77),
.B1(n_86),
.B2(n_13),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_170),
.A2(n_136),
.B1(n_116),
.B2(n_115),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_28),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_115),
.B(n_136),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_113),
.Y(n_173)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_174),
.A2(n_164),
.B(n_148),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_134),
.B(n_129),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_175),
.A2(n_1),
.B(n_2),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_127),
.C(n_118),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_200),
.C(n_143),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_177),
.A2(n_183),
.B(n_196),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_199),
.B1(n_155),
.B2(n_156),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_150),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_189),
.B(n_192),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_85),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_171),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_194),
.A2(n_201),
.B1(n_170),
.B2(n_205),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_135),
.B1(n_12),
.B2(n_14),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_195),
.A2(n_204),
.B1(n_164),
.B2(n_166),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_146),
.A2(n_135),
.B(n_85),
.C(n_83),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_167),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_203),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_161),
.A2(n_153),
.B1(n_156),
.B2(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_167),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_157),
.A2(n_10),
.B1(n_12),
.B2(n_11),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_217),
.B1(n_224),
.B2(n_231),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_178),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_SL g251 ( 
.A(n_208),
.B(n_178),
.C(n_190),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_202),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_210),
.B(n_213),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_184),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_161),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_214),
.B(n_191),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_222),
.C(n_174),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_223),
.B1(n_232),
.B2(n_234),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_227),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_228),
.B(n_230),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_145),
.C(n_142),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_194),
.A2(n_142),
.B1(n_169),
.B2(n_28),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_199),
.A2(n_10),
.B1(n_12),
.B2(n_11),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_31),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_175),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_179),
.A2(n_85),
.B(n_71),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_31),
.B1(n_5),
.B2(n_4),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_182),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_181),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_233),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_196),
.A2(n_6),
.B1(n_11),
.B2(n_3),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_176),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_252),
.Y(n_259)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_221),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_244),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_212),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_254),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_215),
.B(n_186),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_249),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_251),
.A2(n_228),
.B(n_234),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_256),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_209),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_209),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_257),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_185),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_223),
.A2(n_187),
.B1(n_185),
.B2(n_179),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_225),
.C(n_229),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_264),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_225),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_246),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_219),
.B(n_230),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_224),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_218),
.B1(n_217),
.B2(n_207),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_263),
.A2(n_245),
.B1(n_232),
.B2(n_195),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_208),
.C(n_198),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_275),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_288),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_218),
.B1(n_237),
.B2(n_256),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_285),
.Y(n_295)
);

OAI21x1_ASAP7_75t_L g282 ( 
.A1(n_262),
.A2(n_238),
.B(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_270),
.B(n_263),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_284),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_271),
.B(n_241),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_266),
.A2(n_243),
.B1(n_245),
.B2(n_257),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_287),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_198),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_265),
.B(n_180),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_260),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_184),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_291),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_188),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_188),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_269),
.Y(n_294)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_293),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_297),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_264),
.C(n_261),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_276),
.C(n_280),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_274),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_291),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_258),
.C(n_268),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_305),
.C(n_298),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_268),
.C(n_273),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_306),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_304),
.A2(n_272),
.B(n_273),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_236),
.B(n_286),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_310),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_299),
.A2(n_240),
.B1(n_236),
.B2(n_278),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_287),
.B1(n_206),
.B2(n_301),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_295),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_303),
.C(n_305),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_317),
.A2(n_318),
.B(n_319),
.Y(n_322)
);

AOI211xp5_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_313),
.B(n_314),
.C(n_309),
.Y(n_321)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_315),
.A2(n_308),
.B(n_298),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_323),
.A2(n_324),
.B(n_317),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_SL g324 ( 
.A(n_320),
.B(n_302),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_325),
.A2(n_322),
.B(n_320),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_326),
.B(n_301),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_6),
.B(n_2),
.Y(n_329)
);

AO21x1_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_3),
.B(n_1),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_3),
.C(n_1),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_2),
.Y(n_332)
);


endmodule