module fake_aes_1417_n_47 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_47);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_47;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_46;
wire n_30;
wire n_16;
wire n_26;
wire n_33;
wire n_25;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_8), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_7), .B(n_11), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_6), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_13), .Y(n_20) );
BUFx6f_ASAP7_75t_L g21 ( .A(n_4), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_4), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_3), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_21), .Y(n_25) );
OR2x6_ASAP7_75t_L g26 ( .A(n_22), .B(n_0), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
NOR3xp33_ASAP7_75t_L g28 ( .A(n_27), .B(n_16), .C(n_17), .Y(n_28) );
AO21x2_ASAP7_75t_L g29 ( .A1(n_24), .A2(n_18), .B(n_19), .Y(n_29) );
AOI22xp33_ASAP7_75t_L g30 ( .A1(n_26), .A2(n_21), .B1(n_19), .B2(n_18), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
OR2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_26), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
AND2x2_ASAP7_75t_L g34 ( .A(n_32), .B(n_28), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
OR2x2_ASAP7_75t_L g36 ( .A(n_34), .B(n_0), .Y(n_36) );
INVx1_ASAP7_75t_SL g37 ( .A(n_33), .Y(n_37) );
OAI211xp5_ASAP7_75t_SL g38 ( .A1(n_36), .A2(n_25), .B(n_34), .C(n_21), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_35), .Y(n_39) );
OAI22xp33_ASAP7_75t_L g40 ( .A1(n_37), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_40) );
NOR3xp33_ASAP7_75t_L g41 ( .A(n_38), .B(n_1), .C(n_2), .Y(n_41) );
NOR2x1_ASAP7_75t_L g42 ( .A(n_40), .B(n_5), .Y(n_42) );
NAND3xp33_ASAP7_75t_L g43 ( .A(n_39), .B(n_9), .C(n_10), .Y(n_43) );
INVx1_ASAP7_75t_L g44 ( .A(n_42), .Y(n_44) );
NAND2xp5_ASAP7_75t_L g45 ( .A(n_41), .B(n_12), .Y(n_45) );
OAI22xp5_ASAP7_75t_L g46 ( .A1(n_44), .A2(n_45), .B1(n_43), .B2(n_14), .Y(n_46) );
INVx1_ASAP7_75t_L g47 ( .A(n_46), .Y(n_47) );
endmodule