module fake_jpeg_4637_n_109 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_19),
.B(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_23),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_0),
.C(n_1),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_0),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx6p67_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_18),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_18),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_14),
.C(n_1),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_29),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_23),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_37),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_24),
.B1(n_22),
.B2(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_29),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_32),
.B1(n_40),
.B2(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_52),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_49),
.B(n_45),
.Y(n_62)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_57),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_33),
.Y(n_55)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_38),
.B(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_53),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_58),
.B(n_61),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_14),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_27),
.B(n_20),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_50),
.B1(n_43),
.B2(n_27),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_21),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_59),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_11),
.B(n_16),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_72),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_56),
.A3(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_77),
.Y(n_84)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_56),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_81),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_66),
.B(n_54),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_85),
.B(n_21),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_66),
.C(n_51),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_76),
.B1(n_82),
.B2(n_73),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_91),
.B(n_2),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_89),
.B1(n_15),
.B2(n_12),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_75),
.B1(n_69),
.B2(n_70),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_75),
.B1(n_51),
.B2(n_46),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_90),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_78),
.C(n_16),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_95),
.C(n_96),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_3),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_2),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_97),
.B(n_100),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_87),
.C(n_3),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_99),
.B(n_98),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_101),
.B(n_102),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_92),
.Y(n_102)
);

NOR2x1_ASAP7_75t_SL g105 ( 
.A(n_102),
.B(n_93),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_103),
.C(n_4),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_5),
.B(n_7),
.Y(n_107)
);

BUFx24_ASAP7_75t_SL g108 ( 
.A(n_107),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_104),
.Y(n_109)
);


endmodule