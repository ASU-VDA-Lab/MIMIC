module fake_jpeg_9655_n_132 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_4),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_31),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_21),
.A2(n_1),
.B(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx2_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_27),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_20),
.B1(n_19),
.B2(n_14),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_14),
.B1(n_29),
.B2(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_25),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_28),
.C(n_33),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_56),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_32),
.C(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_25),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_64),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_16),
.C(n_29),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_3),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_61),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_37),
.B1(n_34),
.B2(n_20),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_23),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_66),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_19),
.B1(n_18),
.B2(n_23),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_71),
.B1(n_15),
.B2(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_18),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_24),
.B(n_2),
.C(n_3),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_22),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_27),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_10),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_22),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_1),
.Y(n_70)
);

AOI32xp33_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_26),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_15),
.B1(n_27),
.B2(n_26),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_75),
.B1(n_86),
.B2(n_82),
.Y(n_93)
);

NOR3xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_76),
.C(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_85),
.Y(n_91)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_8),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_10),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_11),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_55),
.B(n_59),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_78),
.B(n_76),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_69),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_98),
.C(n_76),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_94),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_63),
.B(n_7),
.C(n_5),
.Y(n_109)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_78),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_53),
.C(n_70),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_65),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_81),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_98),
.A2(n_75),
.B1(n_77),
.B2(n_81),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_102),
.A2(n_104),
.B(n_105),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

FAx1_ASAP7_75t_SL g112 ( 
.A(n_106),
.B(n_89),
.CI(n_96),
.CON(n_112),
.SN(n_112)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_91),
.C(n_99),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_109),
.A2(n_99),
.B1(n_95),
.B2(n_100),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_90),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_115),
.C(n_109),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_103),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_114),
.B1(n_109),
.B2(n_110),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_112),
.B(n_60),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_113),
.C(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_119),
.B(n_120),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_110),
.B(n_84),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_122),
.B(n_60),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_123),
.A2(n_117),
.B(n_118),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_68),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_126),
.C(n_60),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_127),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_128),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_129),
.Y(n_132)
);


endmodule