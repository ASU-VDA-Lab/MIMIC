module fake_jpeg_31461_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_6),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_18),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_7),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_17),
.A2(n_20),
.B1(n_23),
.B2(n_8),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_22),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_10),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_3),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_14),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_12),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_12),
.B(n_8),
.Y(n_24)
);

BUFx24_ASAP7_75t_SL g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_30),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_23),
.A2(n_20),
.B1(n_16),
.B2(n_15),
.Y(n_26)
);

AO21x1_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_31),
.B(n_8),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_17),
.A2(n_8),
.B1(n_15),
.B2(n_19),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_29),
.B1(n_32),
.B2(n_27),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_36),
.B1(n_35),
.B2(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_43),
.B(n_44),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_36),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_45),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_46),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_47)
);


endmodule