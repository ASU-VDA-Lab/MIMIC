module real_aes_6176_n_10 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
output n_10;
wire n_28;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_41;
wire n_34;
wire n_12;
wire n_19;
wire n_40;
wire n_25;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
INVx1_ASAP7_75t_L g21 ( .A(n_0), .Y(n_21) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_1), .Y(n_25) );
AND2x6_ASAP7_75t_L g35 ( .A(n_1), .B(n_27), .Y(n_35) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_2), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_3), .Y(n_18) );
AOI221xp5_ASAP7_75t_L g10 ( .A1(n_4), .A2(n_11), .B1(n_15), .B2(n_28), .C(n_40), .Y(n_10) );
NOR2xp33_ASAP7_75t_L g42 ( .A(n_4), .B(n_30), .Y(n_42) );
INVx2_ASAP7_75t_L g39 ( .A(n_5), .Y(n_39) );
INVx1_ASAP7_75t_L g32 ( .A(n_6), .Y(n_32) );
INVx1_ASAP7_75t_L g38 ( .A(n_7), .Y(n_38) );
INVx1_ASAP7_75t_L g31 ( .A(n_8), .Y(n_31) );
INVx1_ASAP7_75t_L g27 ( .A(n_9), .Y(n_27) );
CKINVDCx20_ASAP7_75t_R g11 ( .A(n_12), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_14), .Y(n_13) );
INVx1_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_16), .B(n_34), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_17), .B(n_22), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_18), .B(n_19), .Y(n_17) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_21), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_23), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_24), .B(n_26), .Y(n_23) );
OAI21xp33_ASAP7_75t_SL g28 ( .A1(n_24), .A2(n_29), .B(n_33), .Y(n_28) );
CKINVDCx16_ASAP7_75t_R g24 ( .A(n_25), .Y(n_24) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_27), .Y(n_26) );
CKINVDCx20_ASAP7_75t_R g29 ( .A(n_30), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_31), .B(n_32), .Y(n_30) );
NOR2xp33_ASAP7_75t_L g40 ( .A(n_34), .B(n_41), .Y(n_40) );
NAND2xp5_ASAP7_75t_SL g34 ( .A(n_35), .B(n_36), .Y(n_34) );
NOR2xp33_ASAP7_75t_L g36 ( .A(n_37), .B(n_39), .Y(n_36) );
HB1xp67_ASAP7_75t_L g37 ( .A(n_38), .Y(n_37) );
INVxp33_ASAP7_75t_L g41 ( .A(n_42), .Y(n_41) );
endmodule