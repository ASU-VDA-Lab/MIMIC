module fake_jpeg_15316_n_212 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_212);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_2),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_26),
.Y(n_56)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_58),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_49),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_29),
.B1(n_20),
.B2(n_21),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_21),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_20),
.B1(n_29),
.B2(n_21),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_29),
.B1(n_20),
.B2(n_27),
.Y(n_51)
);

CKINVDCx9p33_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_59),
.B(n_30),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_65),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_81),
.B1(n_72),
.B2(n_67),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_17),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_41),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_74),
.Y(n_90)
);

AO22x1_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_36),
.B1(n_27),
.B2(n_37),
.Y(n_71)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_72),
.B(n_75),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_41),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_30),
.C(n_19),
.Y(n_102)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_60),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_76),
.B(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_40),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_39),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_39),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_93),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_48),
.B1(n_57),
.B2(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_83),
.B(n_100),
.Y(n_115)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_84),
.B(n_99),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_51),
.B1(n_46),
.B2(n_57),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_87),
.A2(n_92),
.B(n_95),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_27),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_97),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_55),
.B1(n_42),
.B2(n_37),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_69),
.A2(n_27),
.B(n_15),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_19),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_67),
.A2(n_36),
.B1(n_39),
.B2(n_37),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_32),
.B1(n_31),
.B2(n_17),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_103),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_54),
.C(n_32),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_106),
.B(n_101),
.Y(n_130)
);

AND2x6_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_87),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_112),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_80),
.B1(n_31),
.B2(n_71),
.Y(n_111)
);

OA21x2_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_61),
.B(n_79),
.Y(n_133)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_16),
.B(n_25),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_118),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_78),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_119),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_16),
.B(n_25),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_78),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_71),
.B(n_66),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_109),
.B1(n_123),
.B2(n_111),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_96),
.A2(n_61),
.B(n_32),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_15),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_94),
.B1(n_100),
.B2(n_92),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_115),
.B1(n_111),
.B2(n_122),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_88),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_132),
.Y(n_146)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_94),
.A3(n_89),
.B1(n_102),
.B2(n_15),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_86),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_135),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_86),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_122),
.B(n_26),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_15),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_105),
.B(n_109),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_144),
.A2(n_142),
.B(n_138),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_104),
.C(n_116),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_148),
.C(n_153),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_150),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_116),
.C(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_125),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_120),
.C(n_121),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_115),
.B1(n_111),
.B2(n_105),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_156),
.B1(n_4),
.B2(n_5),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_119),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_108),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_146),
.B(n_154),
.Y(n_174)
);

NOR4xp25_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_126),
.C(n_131),
.D(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_127),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_163),
.C(n_164),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_136),
.C(n_126),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_118),
.Y(n_164)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_166),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_133),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_169),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_133),
.C(n_111),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_154),
.B1(n_150),
.B2(n_143),
.Y(n_177)
);

NOR2xp67_ASAP7_75t_SL g172 ( 
.A(n_147),
.B(n_61),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_172),
.A2(n_149),
.B(n_155),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_23),
.B(n_22),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_171),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_176),
.A2(n_180),
.B1(n_166),
.B2(n_183),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_177),
.A2(n_168),
.B1(n_161),
.B2(n_7),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_152),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_183),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_164),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_175),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_188),
.B(n_190),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_161),
.C(n_162),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_191),
.C(n_192),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_189),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_23),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_23),
.C(n_11),
.Y(n_192)
);

AOI322xp5_ASAP7_75t_L g194 ( 
.A1(n_184),
.A2(n_185),
.A3(n_182),
.B1(n_174),
.B2(n_191),
.C1(n_186),
.C2(n_178),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_195),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_184),
.A2(n_178),
.A3(n_23),
.B1(n_12),
.B2(n_14),
.C1(n_13),
.C2(n_7),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_28),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_197),
.B(n_198),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_12),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_5),
.C(n_6),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_200),
.B(n_204),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_193),
.A2(n_5),
.B(n_6),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_202),
.A2(n_203),
.B(n_197),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_28),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_203),
.B(n_6),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_207),
.B(n_208),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_8),
.B1(n_9),
.B2(n_28),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_205),
.B(n_8),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_209),
.Y(n_212)
);


endmodule