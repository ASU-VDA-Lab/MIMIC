module fake_jpeg_22176_n_105 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_10),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_22),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_11),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

NAND3xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_13),
.C(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_41),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_48),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_51),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_18),
.C(n_23),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_29),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_26),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

AO21x1_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_35),
.B(n_33),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_57),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_24),
.B1(n_17),
.B2(n_26),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_56),
.B1(n_13),
.B2(n_23),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_33),
.B(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_24),
.B1(n_14),
.B2(n_21),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_46),
.B(n_45),
.Y(n_77)
);

AND2x6_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_5),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_50),
.C(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_14),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_69),
.B(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_59),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_63),
.B(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_47),
.B1(n_57),
.B2(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_44),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_63),
.C(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_61),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_72),
.B(n_68),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_70),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_25),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_88),
.B(n_92),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_84),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_91),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_68),
.B1(n_62),
.B2(n_20),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_95),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_96),
.B(n_12),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g97 ( 
.A1(n_94),
.A2(n_86),
.A3(n_19),
.B1(n_21),
.B2(n_12),
.C1(n_25),
.C2(n_62),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_99),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

AOI322xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_25),
.A3(n_42),
.B1(n_10),
.B2(n_8),
.C1(n_27),
.C2(n_2),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_100),
.B1(n_2),
.B2(n_3),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_102),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_1),
.Y(n_105)
);


endmodule