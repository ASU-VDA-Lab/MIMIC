module real_aes_6746_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g552 ( .A1(n_0), .A2(n_159), .B(n_553), .C(n_556), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_1), .B(n_497), .Y(n_557) );
INVx1_ASAP7_75t_L g107 ( .A(n_2), .Y(n_107) );
INVx1_ASAP7_75t_L g193 ( .A(n_3), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_4), .B(n_151), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_5), .A2(n_466), .B(n_491), .Y(n_490) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_6), .A2(n_136), .B(n_482), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_7), .A2(n_36), .B1(n_145), .B2(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_8), .B(n_136), .Y(n_162) );
AND2x6_ASAP7_75t_L g160 ( .A(n_9), .B(n_161), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_10), .A2(n_160), .B(n_456), .C(n_458), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_11), .B(n_37), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_11), .B(n_37), .Y(n_122) );
INVx1_ASAP7_75t_L g141 ( .A(n_12), .Y(n_141) );
INVx1_ASAP7_75t_L g186 ( .A(n_13), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_14), .B(n_149), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_15), .B(n_151), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_16), .B(n_137), .Y(n_198) );
AO32x2_ASAP7_75t_L g220 ( .A1(n_17), .A2(n_136), .A3(n_166), .B1(n_177), .B2(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_18), .B(n_145), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_19), .B(n_137), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_20), .A2(n_53), .B1(n_145), .B2(n_223), .Y(n_224) );
AOI22xp33_ASAP7_75t_SL g245 ( .A1(n_21), .A2(n_80), .B1(n_145), .B2(n_149), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_22), .B(n_145), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_23), .A2(n_177), .B(n_456), .C(n_517), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_24), .A2(n_177), .B(n_456), .C(n_485), .Y(n_484) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_25), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_26), .B(n_179), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_27), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_28), .A2(n_466), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_29), .B(n_179), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_30), .A2(n_101), .B1(n_111), .B2(n_750), .Y(n_100) );
INVx2_ASAP7_75t_L g147 ( .A(n_31), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_32), .A2(n_468), .B(n_476), .C(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_33), .B(n_145), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_34), .B(n_179), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_35), .B(n_231), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_38), .B(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_39), .Y(n_462) );
AOI222xp33_ASAP7_75t_SL g124 ( .A1(n_40), .A2(n_78), .B1(n_125), .B2(n_731), .C1(n_732), .C2(n_736), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g731 ( .A(n_40), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_41), .B(n_151), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_42), .B(n_466), .Y(n_483) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_43), .A2(n_77), .B1(n_439), .B2(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_43), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_44), .A2(n_468), .B(n_470), .C(n_476), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_45), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g554 ( .A(n_46), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_47), .A2(n_89), .B1(n_223), .B2(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g471 ( .A(n_48), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_49), .B(n_145), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_50), .B(n_145), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_51), .B(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_52), .B(n_157), .Y(n_156) );
AOI22xp33_ASAP7_75t_SL g202 ( .A1(n_54), .A2(n_58), .B1(n_145), .B2(n_149), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_55), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_56), .B(n_145), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_57), .B(n_145), .Y(n_228) );
INVx1_ASAP7_75t_L g161 ( .A(n_59), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_60), .B(n_466), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_61), .B(n_497), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_62), .A2(n_157), .B(n_189), .C(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_63), .B(n_145), .Y(n_194) );
INVx1_ASAP7_75t_L g140 ( .A(n_64), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_65), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_66), .B(n_151), .Y(n_507) );
AO32x2_ASAP7_75t_L g241 ( .A1(n_67), .A2(n_136), .A3(n_177), .B1(n_242), .B2(n_246), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_68), .B(n_152), .Y(n_459) );
INVx1_ASAP7_75t_L g172 ( .A(n_69), .Y(n_172) );
INVx1_ASAP7_75t_L g212 ( .A(n_70), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g551 ( .A(n_71), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_72), .B(n_473), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_73), .A2(n_456), .B(n_476), .C(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_74), .B(n_149), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_75), .Y(n_492) );
INVx1_ASAP7_75t_L g110 ( .A(n_76), .Y(n_110) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_77), .A2(n_128), .B1(n_438), .B2(n_439), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_77), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_79), .B(n_472), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_81), .B(n_223), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_82), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_83), .B(n_149), .Y(n_216) );
INVx2_ASAP7_75t_L g138 ( .A(n_84), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_85), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_86), .B(n_176), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_87), .B(n_149), .Y(n_148) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_88), .B(n_107), .C(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g119 ( .A(n_88), .B(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g442 ( .A(n_88), .B(n_121), .Y(n_442) );
INVx2_ASAP7_75t_L g730 ( .A(n_88), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_90), .A2(n_99), .B1(n_149), .B2(n_150), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_91), .B(n_466), .Y(n_503) );
INVx1_ASAP7_75t_L g506 ( .A(n_92), .Y(n_506) );
INVxp67_ASAP7_75t_L g495 ( .A(n_93), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_94), .B(n_149), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_95), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g452 ( .A(n_96), .Y(n_452) );
INVx1_ASAP7_75t_L g530 ( .A(n_97), .Y(n_530) );
AND2x2_ASAP7_75t_L g478 ( .A(n_98), .B(n_179), .Y(n_478) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g750 ( .A(n_103), .Y(n_750) );
CKINVDCx12_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
OR2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AND2x2_ASAP7_75t_L g121 ( .A(n_107), .B(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AOI22x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_124), .B1(n_739), .B2(n_740), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_117), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_SL g739 ( .A(n_115), .Y(n_739) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_117), .A2(n_741), .B(n_748), .Y(n_740) );
NOR2xp33_ASAP7_75t_SL g117 ( .A(n_118), .B(n_123), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g749 ( .A(n_119), .Y(n_749) );
NOR2x2_ASAP7_75t_L g738 ( .A(n_120), .B(n_730), .Y(n_738) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g729 ( .A(n_121), .B(n_730), .Y(n_729) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_440), .B1(n_443), .B2(n_727), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_127), .A2(n_733), .B1(n_734), .B2(n_735), .Y(n_732) );
INVx2_ASAP7_75t_L g438 ( .A(n_128), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_128), .A2(n_438), .B1(n_745), .B2(n_746), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g128 ( .A(n_129), .B(n_362), .Y(n_128) );
AND2x2_ASAP7_75t_SL g129 ( .A(n_130), .B(n_320), .Y(n_129) );
NOR4xp25_ASAP7_75t_L g130 ( .A(n_131), .B(n_260), .C(n_296), .D(n_310), .Y(n_130) );
OAI221xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_204), .B1(n_236), .B2(n_247), .C(n_251), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_132), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_180), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_163), .Y(n_134) );
AND2x2_ASAP7_75t_L g257 ( .A(n_135), .B(n_164), .Y(n_257) );
INVx3_ASAP7_75t_L g265 ( .A(n_135), .Y(n_265) );
AND2x2_ASAP7_75t_L g319 ( .A(n_135), .B(n_183), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_135), .B(n_182), .Y(n_355) );
AND2x2_ASAP7_75t_L g413 ( .A(n_135), .B(n_275), .Y(n_413) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_142), .B(n_162), .Y(n_135) );
INVx4_ASAP7_75t_L g203 ( .A(n_136), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_136), .A2(n_483), .B(n_484), .Y(n_482) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_136), .Y(n_489) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g166 ( .A(n_137), .Y(n_166) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g179 ( .A(n_138), .B(n_139), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
OAI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_154), .B(n_160), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_148), .B(n_151), .Y(n_143) );
INVx3_ASAP7_75t_L g211 ( .A(n_145), .Y(n_211) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_145), .Y(n_532) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g223 ( .A(n_146), .Y(n_223) );
BUFx3_ASAP7_75t_L g244 ( .A(n_146), .Y(n_244) );
AND2x6_ASAP7_75t_L g456 ( .A(n_146), .B(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g150 ( .A(n_147), .Y(n_150) );
INVx1_ASAP7_75t_L g158 ( .A(n_147), .Y(n_158) );
INVx2_ASAP7_75t_L g187 ( .A(n_149), .Y(n_187) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_151), .A2(n_169), .B(n_170), .Y(n_168) );
O2A1O1Ixp5_ASAP7_75t_SL g210 ( .A1(n_151), .A2(n_211), .B(n_212), .C(n_213), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_151), .B(n_495), .Y(n_494) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OAI22xp5_ASAP7_75t_SL g242 ( .A1(n_152), .A2(n_176), .B1(n_243), .B2(n_245), .Y(n_242) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_153), .Y(n_176) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_153), .Y(n_191) );
INVx1_ASAP7_75t_L g231 ( .A(n_153), .Y(n_231) );
AND2x2_ASAP7_75t_L g454 ( .A(n_153), .B(n_158), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_153), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_159), .Y(n_154) );
INVx2_ASAP7_75t_L g173 ( .A(n_157), .Y(n_173) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_159), .A2(n_173), .B(n_193), .C(n_194), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_159), .A2(n_176), .B1(n_201), .B2(n_202), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_159), .A2(n_176), .B1(n_222), .B2(n_224), .Y(n_221) );
BUFx3_ASAP7_75t_L g177 ( .A(n_160), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g184 ( .A1(n_160), .A2(n_185), .B(n_192), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_160), .A2(n_210), .B(n_214), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g226 ( .A1(n_160), .A2(n_227), .B(n_232), .Y(n_226) );
NAND2x1p5_ASAP7_75t_L g453 ( .A(n_160), .B(n_454), .Y(n_453) );
AND2x4_ASAP7_75t_L g466 ( .A(n_160), .B(n_454), .Y(n_466) );
INVx4_ASAP7_75t_SL g477 ( .A(n_160), .Y(n_477) );
AND2x2_ASAP7_75t_L g248 ( .A(n_163), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g262 ( .A(n_163), .B(n_183), .Y(n_262) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_164), .B(n_183), .Y(n_277) );
AND2x2_ASAP7_75t_L g289 ( .A(n_164), .B(n_265), .Y(n_289) );
OR2x2_ASAP7_75t_L g291 ( .A(n_164), .B(n_249), .Y(n_291) );
AND2x2_ASAP7_75t_L g326 ( .A(n_164), .B(n_249), .Y(n_326) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_164), .Y(n_371) );
INVx1_ASAP7_75t_L g379 ( .A(n_164), .Y(n_379) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_167), .B(n_178), .Y(n_164) );
OA21x2_ASAP7_75t_L g183 ( .A1(n_165), .A2(n_184), .B(n_195), .Y(n_183) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_166), .B(n_462), .Y(n_461) );
OAI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_171), .B(n_177), .Y(n_167) );
O2A1O1Ixp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_174), .C(n_175), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_173), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_175), .A2(n_233), .B(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx4_ASAP7_75t_L g555 ( .A(n_176), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g199 ( .A(n_177), .B(n_200), .C(n_203), .Y(n_199) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_179), .A2(n_209), .B(n_217), .Y(n_208) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_179), .A2(n_226), .B(n_235), .Y(n_225) );
INVx2_ASAP7_75t_L g246 ( .A(n_179), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_179), .A2(n_465), .B(n_467), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_179), .A2(n_503), .B(n_504), .Y(n_502) );
INVx1_ASAP7_75t_L g523 ( .A(n_179), .Y(n_523) );
OAI221xp5_ASAP7_75t_L g296 ( .A1(n_180), .A2(n_297), .B1(n_301), .B2(n_305), .C(n_306), .Y(n_296) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g256 ( .A(n_181), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_196), .Y(n_181) );
INVx2_ASAP7_75t_L g255 ( .A(n_182), .Y(n_255) );
AND2x2_ASAP7_75t_L g308 ( .A(n_182), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g327 ( .A(n_182), .B(n_265), .Y(n_327) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g390 ( .A(n_183), .B(n_265), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_188), .C(n_189), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_187), .A2(n_459), .B(n_460), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_187), .A2(n_486), .B(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_189), .A2(n_530), .B(n_531), .C(n_532), .Y(n_529) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_190), .A2(n_215), .B(n_216), .Y(n_214) );
INVx4_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g473 ( .A(n_191), .Y(n_473) );
AND2x2_ASAP7_75t_L g312 ( .A(n_196), .B(n_257), .Y(n_312) );
OAI322xp33_ASAP7_75t_L g380 ( .A1(n_196), .A2(n_336), .A3(n_381), .B1(n_383), .B2(n_386), .C1(n_388), .C2(n_392), .Y(n_380) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2x1_ASAP7_75t_L g263 ( .A(n_197), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g276 ( .A(n_197), .Y(n_276) );
AND2x2_ASAP7_75t_L g385 ( .A(n_197), .B(n_265), .Y(n_385) );
AND2x2_ASAP7_75t_L g417 ( .A(n_197), .B(n_289), .Y(n_417) );
OR2x2_ASAP7_75t_L g420 ( .A(n_197), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
INVx1_ASAP7_75t_L g250 ( .A(n_198), .Y(n_250) );
AO21x1_ASAP7_75t_L g249 ( .A1(n_200), .A2(n_203), .B(n_250), .Y(n_249) );
AO21x2_ASAP7_75t_L g450 ( .A1(n_203), .A2(n_451), .B(n_461), .Y(n_450) );
INVx3_ASAP7_75t_L g497 ( .A(n_203), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_203), .B(n_509), .Y(n_508) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_203), .A2(n_527), .B(n_534), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_203), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_218), .Y(n_205) );
INVx1_ASAP7_75t_L g433 ( .A(n_206), .Y(n_433) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_L g238 ( .A(n_207), .B(n_225), .Y(n_238) );
INVx2_ASAP7_75t_L g273 ( .A(n_207), .Y(n_273) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g295 ( .A(n_208), .Y(n_295) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_208), .Y(n_303) );
OR2x2_ASAP7_75t_L g427 ( .A(n_208), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g252 ( .A(n_218), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g292 ( .A(n_218), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g344 ( .A(n_218), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_225), .Y(n_218) );
AND2x2_ASAP7_75t_L g239 ( .A(n_219), .B(n_240), .Y(n_239) );
NOR2xp67_ASAP7_75t_L g299 ( .A(n_219), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g353 ( .A(n_219), .B(n_241), .Y(n_353) );
OR2x2_ASAP7_75t_L g361 ( .A(n_219), .B(n_295), .Y(n_361) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
BUFx2_ASAP7_75t_L g270 ( .A(n_220), .Y(n_270) );
AND2x2_ASAP7_75t_L g280 ( .A(n_220), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g304 ( .A(n_220), .B(n_225), .Y(n_304) );
AND2x2_ASAP7_75t_L g368 ( .A(n_220), .B(n_241), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_225), .B(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_225), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g281 ( .A(n_225), .Y(n_281) );
INVx1_ASAP7_75t_L g286 ( .A(n_225), .Y(n_286) );
AND2x2_ASAP7_75t_L g298 ( .A(n_225), .B(n_299), .Y(n_298) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_225), .Y(n_376) );
INVx1_ASAP7_75t_L g428 ( .A(n_225), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_230), .Y(n_227) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_239), .Y(n_236) );
AND2x2_ASAP7_75t_L g405 ( .A(n_237), .B(n_314), .Y(n_405) );
INVx2_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g332 ( .A(n_239), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g431 ( .A(n_239), .B(n_366), .Y(n_431) );
INVx1_ASAP7_75t_L g253 ( .A(n_240), .Y(n_253) );
AND2x2_ASAP7_75t_L g279 ( .A(n_240), .B(n_273), .Y(n_279) );
BUFx2_ASAP7_75t_L g338 ( .A(n_240), .Y(n_338) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_241), .Y(n_259) );
INVx1_ASAP7_75t_L g269 ( .A(n_241), .Y(n_269) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_244), .Y(n_475) );
INVx2_ASAP7_75t_L g556 ( .A(n_244), .Y(n_556) );
INVx1_ASAP7_75t_L g520 ( .A(n_246), .Y(n_520) );
NOR2xp67_ASAP7_75t_L g407 ( .A(n_247), .B(n_254), .Y(n_407) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AOI32xp33_ASAP7_75t_L g251 ( .A1(n_248), .A2(n_252), .A3(n_254), .B1(n_256), .B2(n_258), .Y(n_251) );
AND2x2_ASAP7_75t_L g391 ( .A(n_248), .B(n_264), .Y(n_391) );
AND2x2_ASAP7_75t_L g429 ( .A(n_248), .B(n_327), .Y(n_429) );
INVx1_ASAP7_75t_L g309 ( .A(n_249), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_253), .B(n_315), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_254), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_254), .B(n_257), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_254), .B(n_326), .Y(n_408) );
OR2x2_ASAP7_75t_L g422 ( .A(n_254), .B(n_291), .Y(n_422) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g349 ( .A(n_255), .B(n_257), .Y(n_349) );
OR2x2_ASAP7_75t_L g358 ( .A(n_255), .B(n_345), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_257), .B(n_308), .Y(n_330) );
INVx2_ASAP7_75t_L g345 ( .A(n_259), .Y(n_345) );
OR2x2_ASAP7_75t_L g360 ( .A(n_259), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g375 ( .A(n_259), .B(n_376), .Y(n_375) );
A2O1A1Ixp33_ASAP7_75t_L g432 ( .A1(n_259), .A2(n_352), .B(n_433), .C(n_434), .Y(n_432) );
OAI321xp33_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_266), .A3(n_271), .B1(n_274), .B2(n_278), .C(n_282), .Y(n_260) );
INVx1_ASAP7_75t_L g373 ( .A(n_261), .Y(n_373) );
NAND2x1p5_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
AND2x2_ASAP7_75t_L g384 ( .A(n_262), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g336 ( .A(n_264), .Y(n_336) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_265), .B(n_379), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g403 ( .A1(n_266), .A2(n_404), .B1(n_406), .B2(n_408), .C(n_409), .Y(n_403) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
AND2x2_ASAP7_75t_L g341 ( .A(n_268), .B(n_315), .Y(n_341) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_269), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g314 ( .A(n_270), .Y(n_314) );
A2O1A1Ixp33_ASAP7_75t_L g356 ( .A1(n_271), .A2(n_312), .B(n_357), .C(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g323 ( .A(n_273), .B(n_280), .Y(n_323) );
BUFx2_ASAP7_75t_L g333 ( .A(n_273), .Y(n_333) );
INVx1_ASAP7_75t_L g348 ( .A(n_273), .Y(n_348) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
OR2x2_ASAP7_75t_L g354 ( .A(n_276), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g437 ( .A(n_276), .Y(n_437) );
INVx1_ASAP7_75t_L g430 ( .A(n_277), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g283 ( .A(n_279), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g387 ( .A(n_279), .B(n_304), .Y(n_387) );
INVx1_ASAP7_75t_L g316 ( .A(n_280), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_287), .B1(n_290), .B2(n_292), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_284), .B(n_400), .Y(n_399) );
INVxp67_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g352 ( .A(n_285), .B(n_353), .Y(n_352) );
BUFx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_SL g315 ( .A(n_286), .B(n_295), .Y(n_315) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g307 ( .A(n_289), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g317 ( .A(n_291), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_294), .A2(n_412), .B1(n_414), .B2(n_415), .C(n_416), .Y(n_411) );
INVx1_ASAP7_75t_L g300 ( .A(n_295), .Y(n_300) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_295), .Y(n_366) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_298), .B(n_417), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g306 ( .A1(n_299), .A2(n_304), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_302), .B(n_312), .Y(n_409) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_L g378 ( .A(n_303), .Y(n_378) );
AND2x2_ASAP7_75t_L g337 ( .A(n_304), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g426 ( .A(n_304), .Y(n_426) );
INVx1_ASAP7_75t_L g342 ( .A(n_307), .Y(n_342) );
INVx1_ASAP7_75t_L g397 ( .A(n_308), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_313), .B1(n_316), .B2(n_317), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_314), .B(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g382 ( .A(n_315), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_315), .B(n_353), .Y(n_419) );
OR2x2_ASAP7_75t_L g392 ( .A(n_316), .B(n_345), .Y(n_392) );
INVx1_ASAP7_75t_L g331 ( .A(n_317), .Y(n_331) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_319), .B(n_370), .Y(n_369) );
NOR3xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_339), .C(n_350), .Y(n_320) );
OAI211xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_324), .B(n_328), .C(n_334), .Y(n_321) );
INVxp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_323), .A2(n_394), .B1(n_398), .B2(n_401), .C(n_403), .Y(n_393) );
INVx1_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
AND2x2_ASAP7_75t_L g335 ( .A(n_326), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g389 ( .A(n_326), .B(n_390), .Y(n_389) );
OAI211xp5_ASAP7_75t_L g374 ( .A1(n_327), .A2(n_375), .B(n_377), .C(n_379), .Y(n_374) );
INVx2_ASAP7_75t_L g421 ( .A(n_327), .Y(n_421) );
OAI21xp5_ASAP7_75t_SL g328 ( .A1(n_329), .A2(n_331), .B(n_332), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g400 ( .A(n_333), .B(n_353), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
OAI21xp5_ASAP7_75t_SL g339 ( .A1(n_340), .A2(n_342), .B(n_343), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI21xp5_ASAP7_75t_SL g343 ( .A1(n_344), .A2(n_346), .B(n_349), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_344), .B(n_373), .Y(n_372) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_349), .B(n_436), .Y(n_435) );
OAI21xp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_354), .B(n_356), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g377 ( .A(n_353), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND4x1_ASAP7_75t_L g362 ( .A(n_363), .B(n_393), .C(n_410), .D(n_432), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_380), .Y(n_363) );
OAI211xp5_ASAP7_75t_SL g364 ( .A1(n_365), .A2(n_369), .B(n_372), .C(n_374), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_368), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_379), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
INVx1_ASAP7_75t_L g414 ( .A(n_389), .Y(n_414) );
INVx2_ASAP7_75t_SL g402 ( .A(n_390), .Y(n_402) );
OR2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g415 ( .A(n_400), .Y(n_415) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_SL g410 ( .A(n_411), .B(n_418), .Y(n_410) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
OAI221xp5_ASAP7_75t_SL g418 ( .A1(n_419), .A2(n_420), .B1(n_422), .B2(n_423), .C(n_424), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_424) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g733 ( .A(n_441), .Y(n_733) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g734 ( .A(n_443), .Y(n_734) );
OR3x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_625), .C(n_690), .Y(n_443) );
NAND4xp25_ASAP7_75t_SL g444 ( .A(n_445), .B(n_566), .C(n_592), .D(n_615), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_498), .B1(n_536), .B2(n_543), .C(n_558), .Y(n_445) );
CKINVDCx14_ASAP7_75t_R g446 ( .A(n_447), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_447), .A2(n_559), .B1(n_583), .B2(n_714), .Y(n_713) );
OR2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_479), .Y(n_447) );
INVx1_ASAP7_75t_SL g619 ( .A(n_448), .Y(n_619) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_463), .Y(n_448) );
OR2x2_ASAP7_75t_L g541 ( .A(n_449), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g561 ( .A(n_449), .B(n_480), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_449), .B(n_488), .Y(n_574) );
AND2x2_ASAP7_75t_L g591 ( .A(n_449), .B(n_463), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_449), .B(n_539), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_449), .B(n_590), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_449), .B(n_479), .Y(n_712) );
AOI211xp5_ASAP7_75t_SL g723 ( .A1(n_449), .A2(n_629), .B(n_724), .C(n_725), .Y(n_723) );
INVx5_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_450), .B(n_480), .Y(n_595) );
AND2x2_ASAP7_75t_L g598 ( .A(n_450), .B(n_481), .Y(n_598) );
OR2x2_ASAP7_75t_L g643 ( .A(n_450), .B(n_480), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_450), .B(n_488), .Y(n_652) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B(n_455), .Y(n_451) );
INVx5_ASAP7_75t_L g469 ( .A(n_456), .Y(n_469) );
INVx5_ASAP7_75t_SL g542 ( .A(n_463), .Y(n_542) );
AND2x2_ASAP7_75t_L g560 ( .A(n_463), .B(n_561), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_463), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g646 ( .A(n_463), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g678 ( .A(n_463), .B(n_488), .Y(n_678) );
OR2x2_ASAP7_75t_L g684 ( .A(n_463), .B(n_574), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_463), .B(n_634), .Y(n_693) );
OR2x6_ASAP7_75t_L g463 ( .A(n_464), .B(n_478), .Y(n_463) );
BUFx2_ASAP7_75t_L g515 ( .A(n_466), .Y(n_515) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_469), .A2(n_477), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g550 ( .A1(n_469), .A2(n_477), .B(n_551), .C(n_552), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_474), .C(n_475), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_472), .A2(n_475), .B(n_506), .C(n_507), .Y(n_505) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_488), .Y(n_479) );
AND2x2_ASAP7_75t_L g575 ( .A(n_480), .B(n_542), .Y(n_575) );
INVx1_ASAP7_75t_SL g588 ( .A(n_480), .Y(n_588) );
OR2x2_ASAP7_75t_L g623 ( .A(n_480), .B(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g629 ( .A(n_480), .B(n_488), .Y(n_629) );
AND2x2_ASAP7_75t_L g687 ( .A(n_480), .B(n_539), .Y(n_687) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_481), .B(n_542), .Y(n_614) );
INVx3_ASAP7_75t_L g539 ( .A(n_488), .Y(n_539) );
OR2x2_ASAP7_75t_L g580 ( .A(n_488), .B(n_542), .Y(n_580) );
AND2x2_ASAP7_75t_L g590 ( .A(n_488), .B(n_588), .Y(n_590) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_488), .Y(n_638) );
AND2x2_ASAP7_75t_L g647 ( .A(n_488), .B(n_561), .Y(n_647) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_496), .Y(n_488) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_497), .A2(n_549), .B(n_557), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_498), .A2(n_664), .B1(n_666), .B2(n_668), .C(n_671), .Y(n_663) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_510), .Y(n_499) );
AND2x2_ASAP7_75t_L g637 ( .A(n_500), .B(n_618), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_500), .B(n_696), .Y(n_700) );
OR2x2_ASAP7_75t_L g721 ( .A(n_500), .B(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_500), .B(n_726), .Y(n_725) );
BUFx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx5_ASAP7_75t_L g568 ( .A(n_501), .Y(n_568) );
AND2x2_ASAP7_75t_L g645 ( .A(n_501), .B(n_512), .Y(n_645) );
AND2x2_ASAP7_75t_L g706 ( .A(n_501), .B(n_585), .Y(n_706) );
AND2x2_ASAP7_75t_L g719 ( .A(n_501), .B(n_539), .Y(n_719) );
OR2x6_ASAP7_75t_L g501 ( .A(n_502), .B(n_508), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_524), .Y(n_510) );
AND2x4_ASAP7_75t_L g546 ( .A(n_511), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g564 ( .A(n_511), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g571 ( .A(n_511), .Y(n_571) );
AND2x2_ASAP7_75t_L g640 ( .A(n_511), .B(n_618), .Y(n_640) );
AND2x2_ASAP7_75t_L g650 ( .A(n_511), .B(n_568), .Y(n_650) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_511), .Y(n_658) );
AND2x2_ASAP7_75t_L g670 ( .A(n_511), .B(n_548), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_511), .B(n_602), .Y(n_674) );
AND2x2_ASAP7_75t_L g711 ( .A(n_511), .B(n_706), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_511), .B(n_585), .Y(n_722) );
OR2x2_ASAP7_75t_L g724 ( .A(n_511), .B(n_660), .Y(n_724) );
INVx5_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g610 ( .A(n_512), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g620 ( .A(n_512), .B(n_565), .Y(n_620) );
AND2x2_ASAP7_75t_L g632 ( .A(n_512), .B(n_548), .Y(n_632) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_512), .Y(n_662) );
AND2x4_ASAP7_75t_L g696 ( .A(n_512), .B(n_547), .Y(n_696) );
OR2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_521), .Y(n_512) );
AOI21xp5_ASAP7_75t_SL g513 ( .A1(n_514), .A2(n_516), .B(n_520), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
BUFx2_ASAP7_75t_L g545 ( .A(n_524), .Y(n_545) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g585 ( .A(n_525), .Y(n_585) );
AND2x2_ASAP7_75t_L g618 ( .A(n_525), .B(n_548), .Y(n_618) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g565 ( .A(n_526), .B(n_548), .Y(n_565) );
BUFx2_ASAP7_75t_L g611 ( .A(n_526), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_533), .Y(n_527) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_538), .B(n_619), .Y(n_698) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_539), .B(n_561), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_539), .B(n_542), .Y(n_600) );
AND2x2_ASAP7_75t_L g655 ( .A(n_539), .B(n_591), .Y(n_655) );
AOI221xp5_ASAP7_75t_SL g592 ( .A1(n_540), .A2(n_593), .B1(n_601), .B2(n_603), .C(n_607), .Y(n_592) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OR2x2_ASAP7_75t_L g587 ( .A(n_541), .B(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g628 ( .A(n_541), .B(n_629), .Y(n_628) );
OAI321xp33_ASAP7_75t_L g635 ( .A1(n_541), .A2(n_594), .A3(n_636), .B1(n_638), .B2(n_639), .C(n_641), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_542), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_545), .B(n_696), .Y(n_714) );
AND2x2_ASAP7_75t_L g601 ( .A(n_546), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_546), .B(n_605), .Y(n_604) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_547), .Y(n_577) );
AND2x2_ASAP7_75t_L g584 ( .A(n_547), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_547), .B(n_659), .Y(n_689) );
INVx1_ASAP7_75t_L g726 ( .A(n_547), .Y(n_726) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_562), .B(n_563), .Y(n_558) );
INVx1_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_560), .A2(n_670), .B(n_719), .C(n_720), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_561), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_561), .B(n_599), .Y(n_665) );
INVx1_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g608 ( .A(n_565), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_565), .B(n_568), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_565), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_565), .B(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_569), .B1(n_581), .B2(n_586), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g582 ( .A(n_568), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g605 ( .A(n_568), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g617 ( .A(n_568), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_568), .B(n_611), .Y(n_653) );
OR2x2_ASAP7_75t_L g660 ( .A(n_568), .B(n_585), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_568), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g710 ( .A(n_568), .B(n_696), .Y(n_710) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_572), .B1(n_576), .B2(n_578), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g616 ( .A(n_571), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g656 ( .A1(n_574), .A2(n_589), .B1(n_657), .B2(n_661), .Y(n_656) );
INVx1_ASAP7_75t_L g704 ( .A(n_575), .Y(n_704) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_579), .A2(n_616), .B1(n_619), .B2(n_620), .C(n_621), .Y(n_615) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g594 ( .A(n_580), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_584), .B(n_650), .Y(n_682) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_585), .Y(n_602) );
INVx1_ASAP7_75t_L g606 ( .A(n_585), .Y(n_606) );
NAND2xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g624 ( .A(n_591), .Y(n_624) );
AND2x2_ASAP7_75t_L g633 ( .A(n_591), .B(n_634), .Y(n_633) );
NAND2xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
INVx2_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g677 ( .A(n_598), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_601), .A2(n_627), .B1(n_630), .B2(n_633), .C(n_635), .Y(n_626) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_605), .B(n_662), .Y(n_661) );
AOI21xp33_ASAP7_75t_SL g607 ( .A1(n_608), .A2(n_609), .B(n_612), .Y(n_607) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
CKINVDCx16_ASAP7_75t_R g709 ( .A(n_612), .Y(n_709) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
OR2x2_ASAP7_75t_L g651 ( .A(n_614), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_SL g672 ( .A(n_617), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_617), .B(n_677), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_620), .B(n_642), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND4xp25_ASAP7_75t_L g625 ( .A(n_626), .B(n_644), .C(n_663), .D(n_676), .Y(n_625) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g634 ( .A(n_629), .Y(n_634) );
INVxp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g667 ( .A(n_638), .B(n_643), .Y(n_667) );
INVxp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AOI211xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B(n_648), .C(n_656), .Y(n_644) );
AOI211xp5_ASAP7_75t_L g715 ( .A1(n_646), .A2(n_688), .B(n_716), .C(n_723), .Y(n_715) );
INVx1_ASAP7_75t_SL g675 ( .A(n_647), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_651), .B1(n_653), .B2(n_654), .Y(n_648) );
INVx1_ASAP7_75t_L g679 ( .A(n_653), .Y(n_679) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_659), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_659), .B(n_670), .Y(n_703) );
INVx2_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g680 ( .A(n_670), .Y(n_680) );
AOI21xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B(n_675), .Y(n_671) );
INVxp33_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AOI322xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .A3(n_680), .B1(n_681), .B2(n_683), .C1(n_685), .C2(n_688), .Y(n_676) );
INVxp67_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND3xp33_ASAP7_75t_SL g690 ( .A(n_691), .B(n_708), .C(n_715), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_694), .B1(n_697), .B2(n_699), .C(n_701), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_SL g707 ( .A(n_696), .Y(n_707) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVxp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_710), .B1(n_711), .B2(n_712), .C(n_713), .Y(n_708) );
NAND2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g735 ( .A(n_728), .Y(n_735) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx3_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVxp67_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
endmodule