module fake_jpeg_16108_n_247 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_38),
.Y(n_55)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_20),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_22),
.B1(n_27),
.B2(n_29),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_35),
.B1(n_39),
.B2(n_36),
.Y(n_60)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_31),
.Y(n_68)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_25),
.C(n_23),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_54),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_22),
.B1(n_32),
.B2(n_20),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_53),
.A2(n_56),
.B1(n_57),
.B2(n_31),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_17),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_35),
.A2(n_22),
.B1(n_32),
.B2(n_18),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_18),
.B1(n_19),
.B2(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_65),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_63),
.B(n_67),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_42),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_66),
.A2(n_69),
.B(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_78),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_0),
.B(n_1),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_34),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_45),
.Y(n_74)
);

OA22x2_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_42),
.B1(n_40),
.B2(n_34),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_39),
.B(n_38),
.C(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_46),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_79),
.B(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_21),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_40),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_43),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_83),
.C(n_89),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_43),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_48),
.B(n_38),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_36),
.B1(n_39),
.B2(n_38),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_87),
.B1(n_36),
.B2(n_40),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_38),
.B(n_33),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_25),
.B(n_42),
.C(n_40),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_47),
.B(n_33),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_58),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_94),
.Y(n_140)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_113),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_98),
.A2(n_101),
.B1(n_71),
.B2(n_75),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_108),
.B1(n_114),
.B2(n_118),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_59),
.A2(n_63),
.B1(n_70),
.B2(n_67),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_66),
.A2(n_30),
.B1(n_28),
.B2(n_21),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_66),
.A2(n_28),
.B1(n_19),
.B2(n_24),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_61),
.A2(n_24),
.B1(n_25),
.B2(n_23),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_61),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_87),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_121),
.B(n_127),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_69),
.B1(n_61),
.B2(n_72),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_128),
.B1(n_143),
.B2(n_100),
.Y(n_156)
);

AO22x1_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_76),
.B1(n_77),
.B2(n_85),
.Y(n_124)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_88),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_126),
.B(n_131),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_111),
.B(n_108),
.Y(n_127)
);

AO21x2_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_94),
.B(n_76),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_81),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_138),
.C(n_143),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_85),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_142),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_64),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_102),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_64),
.Y(n_137)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_73),
.C(n_91),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_111),
.B(n_84),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_141),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_105),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_65),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_135),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_160),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_96),
.B(n_100),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_122),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_128),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_23),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_156),
.A2(n_167),
.B1(n_128),
.B2(n_132),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_99),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_159),
.C(n_162),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_97),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_161),
.B(n_124),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_25),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_140),
.A2(n_113),
.B(n_117),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_138),
.C(n_128),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_117),
.B1(n_3),
.B2(n_5),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_170),
.A2(n_184),
.B1(n_187),
.B2(n_150),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_164),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_180),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_166),
.C(n_158),
.Y(n_190)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_124),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_183),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_185),
.Y(n_191)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_10),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_16),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_167),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_194),
.C(n_197),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_152),
.B(n_149),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_187),
.B(n_173),
.Y(n_214)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_159),
.C(n_146),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_146),
.C(n_156),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_162),
.C(n_147),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_190),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_201),
.B(n_191),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_200),
.B(n_178),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_203),
.B(n_206),
.Y(n_218)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_169),
.B1(n_155),
.B2(n_180),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_8),
.B(n_11),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_182),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_209),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_188),
.A2(n_169),
.B1(n_198),
.B2(n_189),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_210),
.B(n_211),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_174),
.B1(n_170),
.B2(n_172),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_202),
.B(n_151),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_214),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_165),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_6),
.Y(n_225)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_222),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_221),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_2),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_217),
.C(n_218),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_215),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_213),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_227),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_215),
.C(n_209),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_220),
.C(n_225),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_232),
.Y(n_236)
);

NOR2xp67_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_11),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_229),
.C(n_231),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_235),
.Y(n_240)
);

XNOR2x1_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_223),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_12),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_241),
.C(n_236),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_235),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_233),
.B(n_7),
.C(n_14),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_238),
.C(n_12),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_240),
.C(n_7),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_245),
.C(n_7),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_14),
.Y(n_247)
);


endmodule