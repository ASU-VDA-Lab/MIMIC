module real_aes_6428_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1177;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_1066;
wire n_684;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_1175;
wire n_1170;
wire n_778;
wire n_800;
wire n_522;
wire n_1106;
wire n_838;
wire n_933;
wire n_1092;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_673;
wire n_1067;
wire n_518;
wire n_792;
wire n_905;
wire n_878;
wire n_1192;
wire n_665;
wire n_991;
wire n_667;
wire n_1114;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_1123;
wire n_571;
wire n_491;
wire n_694;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_1137;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_551;
wire n_537;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_1160;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_1078;
wire n_495;
wire n_1072;
wire n_892;
wire n_994;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_1098;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_976;
wire n_466;
wire n_636;
wire n_1182;
wire n_559;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_1189;
wire n_726;
wire n_1070;
wire n_1180;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_962;
wire n_693;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_1168;
wire n_755;
wire n_1025;
wire n_1148;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_874;
wire n_796;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_725;
wire n_973;
wire n_455;
wire n_960;
wire n_504;
wire n_671;
wire n_1081;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_1121;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_1135;
wire n_828;
wire n_940;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_1167;
wire n_1100;
wire n_1193;
wire n_1174;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_449;
wire n_417;
wire n_607;
wire n_1006;
wire n_754;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_505;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1103;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_1145;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_1179;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_1171;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_1157;
wire n_471;
wire n_902;
wire n_1105;
wire n_1158;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_1136;
wire n_579;
wire n_699;
wire n_533;
wire n_1187;
wire n_1000;
wire n_1003;
wire n_1014;
wire n_1028;
wire n_1083;
wire n_727;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_1002;
wire n_1155;
wire n_934;
wire n_1165;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1127;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_637;
wire n_526;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_1194;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1071;
wire n_1052;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_1090;
wire n_456;
wire n_717;
wire n_982;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_1162;
wire n_705;
wire n_1191;
wire n_1195;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1186;
wire n_1010;
wire n_811;
wire n_1185;
wire n_1015;
wire n_459;
wire n_558;
wire n_1172;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1184;
wire n_1166;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_1143;
wire n_929;
wire n_686;
wire n_776;
wire n_1190;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_1045;
wire n_871;
wire n_1159;
wire n_474;
wire n_1156;
wire n_829;
wire n_1030;
wire n_988;
wire n_1088;
wire n_1055;
wire n_921;
wire n_597;
wire n_1176;
wire n_483;
wire n_611;
wire n_640;
wire n_1151;
wire n_1036;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_652;
wire n_703;
wire n_1040;
wire n_601;
wire n_500;
wire n_1097;
wire n_661;
wire n_463;
wire n_1076;
wire n_804;
wire n_1101;
wire n_447;
wire n_1033;
wire n_1102;
wire n_1173;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1119;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_SL g938 ( .A1(n_0), .A2(n_177), .B1(n_939), .B2(n_940), .Y(n_938) );
XOR2x2_ASAP7_75t_L g907 ( .A(n_1), .B(n_908), .Y(n_907) );
CKINVDCx20_ASAP7_75t_R g1085 ( .A(n_2), .Y(n_1085) );
OA22x2_ASAP7_75t_L g854 ( .A1(n_3), .A2(n_855), .B1(n_856), .B2(n_882), .Y(n_854) );
CKINVDCx20_ASAP7_75t_R g855 ( .A(n_3), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_4), .A2(n_308), .B1(n_492), .B2(n_1154), .Y(n_1153) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_5), .A2(n_165), .B1(n_575), .B2(n_576), .C(n_577), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_6), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_7), .A2(n_84), .B1(n_763), .B2(n_1157), .Y(n_1156) );
CKINVDCx20_ASAP7_75t_R g1169 ( .A(n_8), .Y(n_1169) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_9), .A2(n_297), .B1(n_544), .B2(n_602), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_10), .A2(n_355), .B1(n_523), .B2(n_524), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_11), .Y(n_708) );
AO22x2_ASAP7_75t_L g424 ( .A1(n_12), .A2(n_222), .B1(n_425), .B2(n_426), .Y(n_424) );
INVx1_ASAP7_75t_L g1134 ( .A(n_12), .Y(n_1134) );
AOI22xp33_ASAP7_75t_SL g656 ( .A1(n_13), .A2(n_207), .B1(n_657), .B2(n_658), .Y(n_656) );
AOI22xp5_ASAP7_75t_SL g997 ( .A1(n_14), .A2(n_393), .B1(n_718), .B2(n_940), .Y(n_997) );
AOI222xp33_ASAP7_75t_L g1070 ( .A1(n_15), .A2(n_59), .B1(n_334), .B2(n_549), .C1(n_583), .C2(n_797), .Y(n_1070) );
AOI22xp5_ASAP7_75t_SL g993 ( .A1(n_16), .A2(n_255), .B1(n_712), .B2(n_808), .Y(n_993) );
AO22x1_ASAP7_75t_L g951 ( .A1(n_17), .A2(n_952), .B1(n_973), .B2(n_974), .Y(n_951) );
INVx1_ASAP7_75t_L g973 ( .A(n_17), .Y(n_973) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_18), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_19), .A2(n_26), .B1(n_540), .B2(n_544), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_20), .A2(n_397), .B1(n_502), .B2(n_565), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_21), .A2(n_326), .B1(n_572), .B2(n_766), .Y(n_1170) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_22), .A2(n_385), .B1(n_866), .B2(n_967), .Y(n_966) );
CKINVDCx20_ASAP7_75t_R g899 ( .A(n_23), .Y(n_899) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_24), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g913 ( .A1(n_25), .A2(n_380), .B1(n_554), .B2(n_720), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_27), .A2(n_272), .B1(n_479), .B2(n_622), .Y(n_898) );
INVx1_ASAP7_75t_L g920 ( .A(n_28), .Y(n_920) );
AOI221xp5_ASAP7_75t_L g1065 ( .A1(n_29), .A2(n_256), .B1(n_576), .B2(n_1066), .C(n_1067), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_30), .A2(n_373), .B1(n_554), .B2(n_1159), .Y(n_1158) );
AOI22xp33_ASAP7_75t_SL g990 ( .A1(n_31), .A2(n_178), .B1(n_918), .B2(n_991), .Y(n_990) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_32), .A2(n_93), .B1(n_451), .B2(n_798), .Y(n_921) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_33), .A2(n_822), .B1(n_850), .B2(n_851), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g850 ( .A(n_33), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g1049 ( .A1(n_34), .A2(n_1050), .B1(n_1071), .B2(n_1072), .Y(n_1049) );
INVx1_ASAP7_75t_L g1071 ( .A(n_34), .Y(n_1071) );
CKINVDCx20_ASAP7_75t_R g1150 ( .A(n_35), .Y(n_1150) );
AO22x2_ASAP7_75t_L g428 ( .A1(n_36), .A2(n_106), .B1(n_425), .B2(n_429), .Y(n_428) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_37), .A2(n_265), .B1(n_477), .B2(n_482), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_38), .A2(n_200), .B1(n_515), .B2(n_866), .Y(n_865) );
AOI22xp33_ASAP7_75t_SL g796 ( .A1(n_39), .A2(n_98), .B1(n_450), .B2(n_797), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g1069 ( .A(n_40), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_41), .A2(n_287), .B1(n_527), .B2(n_614), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g958 ( .A(n_42), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_43), .A2(n_261), .B1(n_533), .B2(n_609), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g1016 ( .A(n_44), .Y(n_1016) );
AOI22xp33_ASAP7_75t_SL g605 ( .A1(n_45), .A2(n_344), .B1(n_606), .B2(n_607), .Y(n_605) );
AOI22xp33_ASAP7_75t_SL g941 ( .A1(n_46), .A2(n_337), .B1(n_767), .B2(n_942), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g1103 ( .A1(n_47), .A2(n_231), .B1(n_518), .B2(n_746), .Y(n_1103) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_48), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g886 ( .A1(n_49), .A2(n_282), .B1(n_488), .B2(n_506), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_50), .A2(n_236), .B1(n_518), .B2(n_524), .Y(n_972) );
AOI222xp33_ASAP7_75t_L g848 ( .A1(n_51), .A2(n_145), .B1(n_303), .B2(n_549), .C1(n_677), .C2(n_849), .Y(n_848) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_52), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g963 ( .A(n_53), .Y(n_963) );
AOI22xp33_ASAP7_75t_SL g929 ( .A1(n_54), .A2(n_195), .B1(n_585), .B2(n_601), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_55), .B(n_547), .Y(n_706) );
AOI222xp33_ASAP7_75t_L g582 ( .A1(n_56), .A2(n_215), .B1(n_327), .B2(n_449), .C1(n_583), .C2(n_585), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_57), .Y(n_435) );
AOI22xp33_ASAP7_75t_SL g1093 ( .A1(n_58), .A2(n_341), .B1(n_507), .B2(n_763), .Y(n_1093) );
CKINVDCx20_ASAP7_75t_R g1061 ( .A(n_60), .Y(n_1061) );
CKINVDCx20_ASAP7_75t_R g1031 ( .A(n_61), .Y(n_1031) );
CKINVDCx20_ASAP7_75t_R g1010 ( .A(n_62), .Y(n_1010) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_63), .Y(n_831) );
AOI22xp5_ASAP7_75t_SL g1077 ( .A1(n_64), .A2(n_1078), .B1(n_1098), .B2(n_1099), .Y(n_1077) );
CKINVDCx16_ASAP7_75t_R g1099 ( .A(n_64), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_65), .A2(n_208), .B1(n_497), .B2(n_501), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_66), .A2(n_102), .B1(n_487), .B2(n_572), .Y(n_969) );
INVx1_ASAP7_75t_L g999 ( .A(n_67), .Y(n_999) );
CKINVDCx20_ASAP7_75t_R g1012 ( .A(n_68), .Y(n_1012) );
CKINVDCx20_ASAP7_75t_R g1090 ( .A(n_69), .Y(n_1090) );
AOI222xp33_ASAP7_75t_L g1113 ( .A1(n_70), .A2(n_204), .B1(n_248), .B2(n_737), .C1(n_738), .C2(n_780), .Y(n_1113) );
AOI22xp33_ASAP7_75t_SL g1034 ( .A1(n_71), .A2(n_209), .B1(n_540), .B2(n_545), .Y(n_1034) );
AOI22xp33_ASAP7_75t_SL g615 ( .A1(n_72), .A2(n_75), .B1(n_616), .B2(n_618), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g947 ( .A1(n_73), .A2(n_277), .B1(n_529), .B2(n_720), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_74), .A2(n_97), .B1(n_529), .B2(n_861), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_76), .A2(n_144), .B1(n_558), .B2(n_665), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_77), .A2(n_262), .B1(n_458), .B2(n_542), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_78), .A2(n_240), .B1(n_624), .B2(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_79), .A2(n_249), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp5_ASAP7_75t_SL g994 ( .A1(n_80), .A2(n_259), .B1(n_715), .B2(n_995), .Y(n_994) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_81), .Y(n_418) );
OA22x2_ASAP7_75t_L g590 ( .A1(n_82), .A2(n_591), .B1(n_592), .B2(n_628), .Y(n_590) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_82), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_83), .Y(n_764) );
AOI22xp33_ASAP7_75t_SL g1097 ( .A1(n_85), .A2(n_127), .B1(n_520), .B2(n_715), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_86), .A2(n_314), .B1(n_565), .B2(n_654), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_87), .A2(n_113), .B1(n_712), .B2(n_1111), .Y(n_1110) );
CKINVDCx20_ASAP7_75t_R g890 ( .A(n_88), .Y(n_890) );
AO22x2_ASAP7_75t_L g432 ( .A1(n_89), .A2(n_264), .B1(n_425), .B2(n_426), .Y(n_432) );
INVx1_ASAP7_75t_L g1131 ( .A(n_89), .Y(n_1131) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_90), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_91), .A2(n_186), .B1(n_544), .B2(n_776), .Y(n_775) );
AOI22xp33_ASAP7_75t_SL g805 ( .A1(n_92), .A2(n_328), .B1(n_626), .B2(n_806), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_94), .Y(n_836) );
AOI22xp5_ASAP7_75t_SL g998 ( .A1(n_95), .A2(n_213), .B1(n_497), .B2(n_529), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_96), .A2(n_307), .B1(n_520), .B2(n_660), .Y(n_1112) );
AOI211xp5_ASAP7_75t_L g807 ( .A1(n_99), .A2(n_808), .B(n_809), .C(n_812), .Y(n_807) );
AOI22xp33_ASAP7_75t_SL g800 ( .A1(n_100), .A2(n_293), .B1(n_606), .B2(n_607), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_101), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_103), .A2(n_201), .B1(n_536), .B2(n_881), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_104), .A2(n_111), .B1(n_737), .B2(n_738), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_105), .A2(n_180), .B1(n_542), .B2(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g1135 ( .A(n_106), .Y(n_1135) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_107), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g1007 ( .A(n_108), .Y(n_1007) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_109), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g1068 ( .A(n_110), .Y(n_1068) );
CKINVDCx20_ASAP7_75t_R g1183 ( .A(n_112), .Y(n_1183) );
AOI22xp33_ASAP7_75t_SL g1108 ( .A1(n_114), .A2(n_345), .B1(n_542), .B2(n_544), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_115), .A2(n_363), .B1(n_523), .B2(n_612), .Y(n_770) );
AOI22xp33_ASAP7_75t_SL g945 ( .A1(n_116), .A2(n_199), .B1(n_507), .B2(n_946), .Y(n_945) );
CKINVDCx20_ASAP7_75t_R g1142 ( .A(n_117), .Y(n_1142) );
CKINVDCx20_ASAP7_75t_R g1167 ( .A(n_118), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_119), .B(n_533), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_120), .A2(n_342), .B1(n_482), .B2(n_665), .Y(n_1038) );
AOI22xp33_ASAP7_75t_SL g933 ( .A1(n_121), .A2(n_211), .B1(n_934), .B2(n_935), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_122), .A2(n_370), .B1(n_477), .B2(n_501), .Y(n_1041) );
CKINVDCx20_ASAP7_75t_R g1179 ( .A(n_123), .Y(n_1179) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_124), .A2(n_280), .B1(n_621), .B2(n_622), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_125), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_126), .A2(n_139), .B1(n_457), .B2(n_550), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_128), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_129), .A2(n_347), .B1(n_492), .B2(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g1180 ( .A(n_130), .Y(n_1180) );
AOI22xp33_ASAP7_75t_SL g879 ( .A1(n_131), .A2(n_257), .B1(n_606), .B2(n_607), .Y(n_879) );
AOI22xp33_ASAP7_75t_SL g985 ( .A1(n_132), .A2(n_354), .B1(n_550), .B2(n_585), .Y(n_985) );
AOI22xp33_ASAP7_75t_SL g867 ( .A1(n_133), .A2(n_206), .B1(n_868), .B2(n_870), .Y(n_867) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_134), .A2(n_153), .B1(n_624), .B2(n_626), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_135), .A2(n_190), .B1(n_533), .B2(n_536), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_136), .A2(n_371), .B1(n_501), .B2(n_524), .Y(n_1024) );
XNOR2x2_ASAP7_75t_L g511 ( .A(n_137), .B(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_138), .A2(n_151), .B1(n_626), .B2(n_746), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g1051 ( .A1(n_140), .A2(n_217), .B1(n_477), .B2(n_1052), .C(n_1054), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_141), .B(n_538), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g1172 ( .A(n_142), .Y(n_1172) );
AND2x6_ASAP7_75t_L g401 ( .A(n_143), .B(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g1128 ( .A(n_143), .Y(n_1128) );
AOI22xp33_ASAP7_75t_SL g717 ( .A1(n_146), .A2(n_379), .B1(n_565), .B2(n_718), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_147), .A2(n_188), .B1(n_505), .B2(n_507), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g1081 ( .A(n_148), .Y(n_1081) );
NAND2xp5_ASAP7_75t_SL g932 ( .A(n_149), .B(n_575), .Y(n_932) );
CKINVDCx20_ASAP7_75t_R g959 ( .A(n_150), .Y(n_959) );
AOI22xp33_ASAP7_75t_SL g719 ( .A1(n_152), .A2(n_358), .B1(n_612), .B2(n_720), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g910 ( .A1(n_154), .A2(n_191), .B1(n_558), .B2(n_614), .Y(n_910) );
NAND2xp5_ASAP7_75t_SL g931 ( .A(n_155), .B(n_609), .Y(n_931) );
AOI22xp33_ASAP7_75t_SL g1032 ( .A1(n_156), .A2(n_276), .B1(n_449), .B2(n_548), .Y(n_1032) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_157), .Y(n_825) );
CKINVDCx20_ASAP7_75t_R g1106 ( .A(n_158), .Y(n_1106) );
AO22x1_ASAP7_75t_L g551 ( .A1(n_159), .A2(n_552), .B1(n_587), .B2(n_588), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_159), .Y(n_587) );
AOI22xp33_ASAP7_75t_SL g679 ( .A1(n_160), .A2(n_181), .B1(n_505), .B2(n_680), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_161), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g838 ( .A(n_162), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g1175 ( .A(n_163), .Y(n_1175) );
AOI222xp33_ASAP7_75t_L g546 ( .A1(n_164), .A2(n_210), .B1(n_351), .B2(n_547), .C1(n_548), .C2(n_549), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_166), .A2(n_312), .B1(n_657), .B2(n_746), .Y(n_971) );
AOI22xp33_ASAP7_75t_SL g801 ( .A1(n_167), .A2(n_241), .B1(n_533), .B2(n_609), .Y(n_801) );
AO22x2_ASAP7_75t_L g434 ( .A1(n_168), .A2(n_258), .B1(n_425), .B2(n_429), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g1132 ( .A(n_168), .B(n_1133), .Y(n_1132) );
CKINVDCx20_ASAP7_75t_R g1002 ( .A(n_169), .Y(n_1002) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_170), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_171), .Y(n_813) );
AOI22xp33_ASAP7_75t_SL g897 ( .A1(n_172), .A2(n_300), .B1(n_499), .B2(n_508), .Y(n_897) );
AOI221xp5_ASAP7_75t_L g1059 ( .A1(n_173), .A2(n_198), .B1(n_515), .B2(n_558), .C(n_1060), .Y(n_1059) );
AOI22xp33_ASAP7_75t_SL g1019 ( .A1(n_174), .A2(n_184), .B1(n_523), .B2(n_1020), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g803 ( .A1(n_175), .A2(n_275), .B1(n_612), .B2(n_804), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_176), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_179), .A2(n_203), .B1(n_505), .B2(n_720), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_182), .A2(n_266), .B1(n_479), .B2(n_520), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_183), .A2(n_189), .B1(n_536), .B2(n_881), .Y(n_1035) );
AOI22xp33_ASAP7_75t_SL g1021 ( .A1(n_185), .A2(n_335), .B1(n_767), .B2(n_868), .Y(n_1021) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_187), .A2(n_202), .B1(n_515), .B2(n_554), .C(n_555), .Y(n_553) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_192), .A2(n_399), .B(n_407), .C(n_1136), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_193), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g1145 ( .A(n_194), .Y(n_1145) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_196), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_197), .A2(n_310), .B1(n_627), .B2(n_660), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g1163 ( .A1(n_205), .A2(n_1164), .B1(n_1188), .B2(n_1189), .Y(n_1163) );
INVx1_ASAP7_75t_L g1188 ( .A(n_205), .Y(n_1188) );
XNOR2xp5_ASAP7_75t_L g790 ( .A(n_212), .B(n_791), .Y(n_790) );
AOI22xp33_ASAP7_75t_SL g711 ( .A1(n_214), .A2(n_250), .B1(n_624), .B2(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g713 ( .A1(n_216), .A2(n_239), .B1(n_714), .B2(n_715), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g563 ( .A1(n_218), .A2(n_244), .B1(n_564), .B2(n_565), .C(n_566), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_219), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_220), .A2(n_348), .B1(n_766), .B2(n_767), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_221), .A2(n_246), .B1(n_565), .B2(n_627), .Y(n_914) );
NAND2xp5_ASAP7_75t_SL g989 ( .A(n_223), .B(n_575), .Y(n_989) );
CKINVDCx20_ASAP7_75t_R g1182 ( .A(n_224), .Y(n_1182) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_225), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_226), .A2(n_362), .B1(n_550), .B2(n_598), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g1176 ( .A1(n_227), .A2(n_247), .B1(n_804), .B2(n_1111), .Y(n_1176) );
CKINVDCx20_ASAP7_75t_R g1062 ( .A(n_228), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_229), .A2(n_271), .B1(n_517), .B2(n_666), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_230), .A2(n_283), .B1(n_598), .B2(n_1147), .Y(n_1146) );
AOI22xp33_ASAP7_75t_SL g486 ( .A1(n_232), .A2(n_315), .B1(n_487), .B2(n_492), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_233), .B(n_767), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_234), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_235), .A2(n_369), .B1(n_558), .B2(n_564), .Y(n_1094) );
OA22x2_ASAP7_75t_L g695 ( .A1(n_237), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_237), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g559 ( .A(n_238), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_242), .A2(n_260), .B1(n_654), .B2(n_665), .Y(n_1104) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_243), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_245), .A2(n_339), .B1(n_515), .B2(n_518), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g1015 ( .A(n_251), .Y(n_1015) );
CKINVDCx20_ASAP7_75t_R g984 ( .A(n_252), .Y(n_984) );
AOI22xp33_ASAP7_75t_SL g664 ( .A1(n_253), .A2(n_304), .B1(n_665), .B2(n_666), .Y(n_664) );
AND2x2_ASAP7_75t_L g405 ( .A(n_254), .B(n_406), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_263), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_267), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_268), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_269), .A2(n_758), .B1(n_785), .B2(n_786), .Y(n_757) );
INVx1_ASAP7_75t_L g785 ( .A(n_269), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g956 ( .A(n_270), .Y(n_956) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_273), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_274), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g1143 ( .A(n_278), .Y(n_1143) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_279), .Y(n_774) );
OA22x2_ASAP7_75t_L g1025 ( .A1(n_281), .A2(n_1026), .B1(n_1027), .B2(n_1043), .Y(n_1025) );
CKINVDCx20_ASAP7_75t_R g1026 ( .A(n_281), .Y(n_1026) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_284), .Y(n_755) );
AOI22xp33_ASAP7_75t_SL g1023 ( .A1(n_285), .A2(n_305), .B1(n_763), .B2(n_863), .Y(n_1023) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_286), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_288), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_289), .Y(n_462) );
OA22x2_ASAP7_75t_L g722 ( .A1(n_290), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_722) );
CKINVDCx16_ASAP7_75t_R g723 ( .A(n_290), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_291), .B(n_575), .Y(n_1107) );
AOI22xp5_ASAP7_75t_L g911 ( .A1(n_292), .A2(n_360), .B1(n_658), .B2(n_715), .Y(n_911) );
INVx1_ASAP7_75t_L g425 ( .A(n_294), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_294), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_295), .Y(n_1013) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_296), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_298), .A2(n_350), .B1(n_487), .B2(n_660), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_299), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g843 ( .A1(n_301), .A2(n_395), .B1(n_536), .B2(n_575), .C(n_844), .Y(n_843) );
AOI22xp33_ASAP7_75t_SL g859 ( .A1(n_302), .A2(n_377), .B1(n_507), .B2(n_806), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_306), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_309), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g1057 ( .A(n_311), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g955 ( .A(n_313), .Y(n_955) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_316), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_317), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_318), .A2(n_924), .B1(n_925), .B2(n_948), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_318), .Y(n_924) );
XNOR2x1_ASAP7_75t_L g632 ( .A(n_319), .B(n_633), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g1088 ( .A(n_320), .Y(n_1088) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_321), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_322), .Y(n_875) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_323), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_324), .A2(n_367), .B1(n_545), .B2(n_918), .Y(n_917) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_325), .Y(n_682) );
INVx1_ASAP7_75t_L g406 ( .A(n_329), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g1151 ( .A(n_330), .Y(n_1151) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_331), .Y(n_447) );
INVx1_ASAP7_75t_L g402 ( .A(n_332), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_333), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g1187 ( .A(n_336), .Y(n_1187) );
AOI22xp33_ASAP7_75t_SL g1096 ( .A1(n_338), .A2(n_376), .B1(n_517), .B2(n_554), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_340), .A2(n_386), .B1(n_451), .B2(n_607), .Y(n_643) );
XOR2x2_ASAP7_75t_L g414 ( .A(n_343), .B(n_415), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_346), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_349), .B(n_674), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_352), .A2(n_384), .B1(n_544), .B2(n_602), .Y(n_671) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_353), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_356), .A2(n_396), .B1(n_576), .B2(n_674), .Y(n_916) );
CKINVDCx20_ASAP7_75t_R g1055 ( .A(n_357), .Y(n_1055) );
CKINVDCx20_ASAP7_75t_R g1082 ( .A(n_359), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_361), .A2(n_372), .B1(n_527), .B2(n_529), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_364), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_365), .A2(n_388), .B1(n_520), .B2(n_767), .Y(n_1042) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_366), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_368), .B(n_538), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_374), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_375), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g960 ( .A(n_378), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_381), .B(n_457), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_382), .Y(n_928) );
CKINVDCx20_ASAP7_75t_R g1006 ( .A(n_383), .Y(n_1006) );
CKINVDCx20_ASAP7_75t_R g1114 ( .A(n_387), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_389), .B(n_988), .Y(n_987) );
CKINVDCx20_ASAP7_75t_R g1184 ( .A(n_390), .Y(n_1184) );
CKINVDCx20_ASAP7_75t_R g962 ( .A(n_391), .Y(n_962) );
CKINVDCx20_ASAP7_75t_R g1186 ( .A(n_392), .Y(n_1186) );
XOR2xp5_ASAP7_75t_L g1137 ( .A(n_394), .B(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_402), .Y(n_1127) );
OAI21xp5_ASAP7_75t_L g1194 ( .A1(n_403), .A2(n_1126), .B(n_1195), .Y(n_1194) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_976), .B1(n_1121), .B2(n_1122), .C(n_1123), .Y(n_407) );
INVx1_ASAP7_75t_L g1122 ( .A(n_408), .Y(n_1122) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_688), .B2(n_689), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_589), .B1(n_686), .B2(n_687), .Y(n_410) );
INVx1_ASAP7_75t_L g686 ( .A(n_411), .Y(n_686) );
XOR2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_551), .Y(n_411) );
OAI22xp5_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_414), .B1(n_510), .B2(n_511), .Y(n_412) );
OA22x2_ASAP7_75t_L g630 ( .A1(n_413), .A2(n_414), .B1(n_631), .B2(n_683), .Y(n_630) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_474), .Y(n_415) );
NOR3xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_441), .C(n_461), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_435), .B2(n_436), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g954 ( .A1(n_419), .A2(n_638), .B1(n_955), .B2(n_956), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g1178 ( .A1(n_419), .A2(n_1083), .B1(n_1179), .B2(n_1180), .Y(n_1178) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_421), .A2(n_636), .B1(n_637), .B2(n_638), .Y(n_635) );
BUFx3_ASAP7_75t_L g702 ( .A(n_421), .Y(n_702) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_421), .Y(n_730) );
OR2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_430), .Y(n_421) );
INVx2_ASAP7_75t_L g500 ( .A(n_422), .Y(n_500) );
OR2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_428), .Y(n_422) );
AND2x2_ASAP7_75t_L g440 ( .A(n_423), .B(n_428), .Y(n_440) );
AND2x2_ASAP7_75t_L g481 ( .A(n_423), .B(n_460), .Y(n_481) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g444 ( .A(n_424), .B(n_428), .Y(n_444) );
AND2x2_ASAP7_75t_L g454 ( .A(n_424), .B(n_434), .Y(n_454) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_427), .Y(n_429) );
INVx2_ASAP7_75t_L g460 ( .A(n_428), .Y(n_460) );
INVx1_ASAP7_75t_L g494 ( .A(n_428), .Y(n_494) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_431), .B(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g503 ( .A(n_431), .B(n_481), .Y(n_503) );
AND2x4_ASAP7_75t_L g535 ( .A(n_431), .B(n_500), .Y(n_535) );
AND2x6_ASAP7_75t_L g538 ( .A(n_431), .B(n_440), .Y(n_538) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g446 ( .A(n_432), .Y(n_446) );
INVx1_ASAP7_75t_L g453 ( .A(n_432), .Y(n_453) );
INVx1_ASAP7_75t_L g473 ( .A(n_432), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_432), .B(n_434), .Y(n_485) );
AND2x2_ASAP7_75t_L g445 ( .A(n_433), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g491 ( .A(n_434), .B(n_473), .Y(n_491) );
OAI221xp5_ASAP7_75t_SL g772 ( .A1(n_436), .A2(n_730), .B1(n_773), .B2(n_774), .C(n_775), .Y(n_772) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_438), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_700) );
BUFx3_ASAP7_75t_L g732 ( .A(n_438), .Y(n_732) );
OAI22xp5_ASAP7_75t_SL g1005 ( .A1(n_438), .A2(n_730), .B1(n_1006), .B2(n_1007), .Y(n_1005) );
BUFx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g639 ( .A(n_439), .Y(n_639) );
AND2x2_ASAP7_75t_L g490 ( .A(n_440), .B(n_491), .Y(n_490) );
AND2x4_ASAP7_75t_L g506 ( .A(n_440), .B(n_445), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_440), .B(n_491), .Y(n_569) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_447), .B1(n_448), .B2(n_455), .C(n_456), .Y(n_441) );
OAI21xp33_ASAP7_75t_L g1144 ( .A1(n_442), .A2(n_1145), .B(n_1146), .Y(n_1144) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx3_ASAP7_75t_L g547 ( .A(n_443), .Y(n_547) );
INVx4_ASAP7_75t_L g584 ( .A(n_443), .Y(n_584) );
BUFx6f_ASAP7_75t_L g780 ( .A(n_443), .Y(n_780) );
INVx2_ASAP7_75t_SL g1011 ( .A(n_443), .Y(n_1011) );
INVx2_ASAP7_75t_L g1030 ( .A(n_443), .Y(n_1030) );
AND2x6_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx1_ASAP7_75t_L g470 ( .A(n_444), .Y(n_470) );
AND2x4_ASAP7_75t_L g545 ( .A(n_444), .B(n_472), .Y(n_545) );
AND2x2_ASAP7_75t_L g480 ( .A(n_445), .B(n_481), .Y(n_480) );
AND2x6_ASAP7_75t_L g499 ( .A(n_445), .B(n_500), .Y(n_499) );
OAI222xp33_ASAP7_75t_L g957 ( .A1(n_448), .A2(n_646), .B1(n_779), .B2(n_958), .C1(n_959), .C2(n_960), .Y(n_957) );
OAI222xp33_ASAP7_75t_L g1181 ( .A1(n_448), .A2(n_597), .B1(n_794), .B2(n_1182), .C1(n_1183), .C2(n_1184), .Y(n_1181) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx2_ASAP7_75t_L g783 ( .A(n_450), .Y(n_783) );
INVx2_ASAP7_75t_L g1148 ( .A(n_450), .Y(n_1148) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx12f_ASAP7_75t_L g550 ( .A(n_451), .Y(n_550) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_451), .Y(n_602) );
INVx1_ASAP7_75t_L g876 ( .A(n_451), .Y(n_876) );
AND2x4_ASAP7_75t_L g451 ( .A(n_452), .B(n_454), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g459 ( .A(n_453), .B(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g458 ( .A(n_454), .B(n_459), .Y(n_458) );
NAND2x1p5_ASAP7_75t_L g464 ( .A(n_454), .B(n_465), .Y(n_464) );
AND2x4_ASAP7_75t_L g542 ( .A(n_454), .B(n_543), .Y(n_542) );
INVx4_ASAP7_75t_L g586 ( .A(n_457), .Y(n_586) );
BUFx2_ASAP7_75t_L g737 ( .A(n_457), .Y(n_737) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g548 ( .A(n_458), .Y(n_548) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_458), .Y(n_598) );
BUFx4f_ASAP7_75t_SL g677 ( .A(n_458), .Y(n_677) );
BUFx6f_ASAP7_75t_L g798 ( .A(n_458), .Y(n_798) );
INVx1_ASAP7_75t_L g465 ( .A(n_460), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B1(n_466), .B2(n_467), .Y(n_461) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g579 ( .A(n_464), .Y(n_579) );
INVx4_ASAP7_75t_L g649 ( .A(n_464), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_464), .A2(n_469), .B1(n_708), .B2(n_709), .Y(n_707) );
OAI22xp33_ASAP7_75t_SL g740 ( .A1(n_464), .A2(n_467), .B1(n_741), .B2(n_742), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g1141 ( .A1(n_464), .A2(n_581), .B1(n_1142), .B2(n_1143), .Y(n_1141) );
AND2x2_ASAP7_75t_L g666 ( .A(n_465), .B(n_484), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_467), .A2(n_579), .B1(n_962), .B2(n_963), .Y(n_961) );
OAI22xp5_ASAP7_75t_SL g1014 ( .A1(n_467), .A2(n_579), .B1(n_1015), .B2(n_1016), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g1185 ( .A1(n_467), .A2(n_579), .B1(n_1186), .B2(n_1187), .Y(n_1185) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g581 ( .A(n_468), .Y(n_581) );
CKINVDCx16_ASAP7_75t_R g468 ( .A(n_469), .Y(n_468) );
BUFx2_ASAP7_75t_L g847 ( .A(n_469), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_469), .A2(n_1088), .B1(n_1089), .B2(n_1090), .Y(n_1087) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_495), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_486), .Y(n_475) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OAI221xp5_ASAP7_75t_SL g1171 ( .A1(n_478), .A2(n_1172), .B1(n_1173), .B2(n_1175), .C(n_1176), .Y(n_1171) );
INVx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx3_ASAP7_75t_L g523 ( .A(n_479), .Y(n_523) );
BUFx3_ASAP7_75t_L g866 ( .A(n_479), .Y(n_866) );
BUFx6f_ASAP7_75t_L g946 ( .A(n_479), .Y(n_946) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx2_ASAP7_75t_SL g554 ( .A(n_480), .Y(n_554) );
INVx2_ASAP7_75t_L g625 ( .A(n_480), .Y(n_625) );
BUFx2_ASAP7_75t_SL g808 ( .A(n_480), .Y(n_808) );
AND2x4_ASAP7_75t_L g483 ( .A(n_481), .B(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g509 ( .A(n_481), .B(n_491), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_481), .B(n_491), .Y(n_562) );
BUFx2_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
BUFx3_ASAP7_75t_L g518 ( .A(n_483), .Y(n_518) );
BUFx3_ASAP7_75t_L g565 ( .A(n_483), .Y(n_565) );
BUFx3_ASAP7_75t_L g622 ( .A(n_483), .Y(n_622) );
INVx1_ASAP7_75t_L g756 ( .A(n_483), .Y(n_756) );
BUFx2_ASAP7_75t_SL g763 ( .A(n_483), .Y(n_763) );
BUFx3_ASAP7_75t_L g829 ( .A(n_483), .Y(n_829) );
BUFx2_ASAP7_75t_L g940 ( .A(n_483), .Y(n_940) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OR2x6_ASAP7_75t_L g493 ( .A(n_485), .B(n_494), .Y(n_493) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g869 ( .A(n_488), .Y(n_869) );
BUFx2_ASAP7_75t_L g995 ( .A(n_488), .Y(n_995) );
INVx4_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx3_ASAP7_75t_L g520 ( .A(n_489), .Y(n_520) );
INVx1_ASAP7_75t_L g617 ( .A(n_489), .Y(n_617) );
INVx2_ASAP7_75t_L g658 ( .A(n_489), .Y(n_658) );
INVx5_ASAP7_75t_L g714 ( .A(n_489), .Y(n_714) );
BUFx3_ASAP7_75t_L g943 ( .A(n_489), .Y(n_943) );
INVx8_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx6_ASAP7_75t_SL g573 ( .A(n_493), .Y(n_573) );
INVx1_ASAP7_75t_SL g767 ( .A(n_493), .Y(n_767) );
INVx1_ASAP7_75t_SL g870 ( .A(n_493), .Y(n_870) );
INVx1_ASAP7_75t_L g543 ( .A(n_494), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_504), .Y(n_495) );
INVx1_ASAP7_75t_L g837 ( .A(n_497), .Y(n_837) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g564 ( .A(n_498), .Y(n_564) );
INVx4_ASAP7_75t_L g720 ( .A(n_498), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_498), .B(n_813), .Y(n_812) );
INVx4_ASAP7_75t_L g1157 ( .A(n_498), .Y(n_1157) );
OAI221xp5_ASAP7_75t_SL g1166 ( .A1(n_498), .A2(n_1167), .B1(n_1168), .B2(n_1169), .C(n_1170), .Y(n_1166) );
INVx11_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx11_ASAP7_75t_L g528 ( .A(n_499), .Y(n_528) );
BUFx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_503), .Y(n_517) );
BUFx3_ASAP7_75t_L g627 ( .A(n_503), .Y(n_627) );
BUFx3_ASAP7_75t_L g712 ( .A(n_503), .Y(n_712) );
INVx2_ASAP7_75t_L g968 ( .A(n_503), .Y(n_968) );
BUFx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx6_ASAP7_75t_L g530 ( .A(n_506), .Y(n_530) );
BUFx3_ASAP7_75t_L g612 ( .A(n_506), .Y(n_612) );
BUFx3_ASAP7_75t_L g1020 ( .A(n_506), .Y(n_1020) );
BUFx4f_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g525 ( .A(n_508), .Y(n_525) );
BUFx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx3_ASAP7_75t_L g614 ( .A(n_509), .Y(n_614) );
BUFx3_ASAP7_75t_L g665 ( .A(n_509), .Y(n_665) );
BUFx3_ASAP7_75t_L g718 ( .A(n_509), .Y(n_718) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND4xp75_ASAP7_75t_L g512 ( .A(n_513), .B(n_521), .C(n_531), .D(n_546), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_519), .Y(n_513) );
INVx4_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx3_ASAP7_75t_L g939 ( .A(n_516), .Y(n_939) );
INVx4_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_526), .Y(n_521) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_SL g1056 ( .A(n_527), .Y(n_1056) );
INVx4_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g621 ( .A(n_528), .Y(n_621) );
INVx2_ASAP7_75t_SL g680 ( .A(n_528), .Y(n_680) );
INVx2_ASAP7_75t_L g746 ( .A(n_528), .Y(n_746) );
INVx5_ASAP7_75t_SL g863 ( .A(n_528), .Y(n_863) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g558 ( .A(n_530), .Y(n_558) );
INVx2_ASAP7_75t_L g657 ( .A(n_530), .Y(n_657) );
INVx3_ASAP7_75t_L g1111 ( .A(n_530), .Y(n_1111) );
AND2x2_ASAP7_75t_SL g531 ( .A(n_532), .B(n_539), .Y(n_531) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_533), .Y(n_575) );
INVx5_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g674 ( .A(n_534), .Y(n_674) );
INVx2_ASAP7_75t_L g881 ( .A(n_534), .Y(n_881) );
INVx4_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_SL g988 ( .A(n_537), .Y(n_988) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
BUFx4f_ASAP7_75t_L g576 ( .A(n_538), .Y(n_576) );
BUFx2_ASAP7_75t_L g609 ( .A(n_538), .Y(n_609) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g934 ( .A(n_541), .Y(n_934) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx2_ASAP7_75t_L g606 ( .A(n_542), .Y(n_606) );
BUFx2_ASAP7_75t_L g776 ( .A(n_542), .Y(n_776) );
BUFx3_ASAP7_75t_L g918 ( .A(n_542), .Y(n_918) );
INVx1_ASAP7_75t_SL g936 ( .A(n_544), .Y(n_936) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx3_ASAP7_75t_L g607 ( .A(n_545), .Y(n_607) );
BUFx2_ASAP7_75t_SL g991 ( .A(n_545), .Y(n_991) );
INVx3_ASAP7_75t_L g642 ( .A(n_547), .Y(n_642) );
INVx1_ASAP7_75t_L g646 ( .A(n_548), .Y(n_646) );
BUFx4f_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g739 ( .A(n_550), .Y(n_739) );
INVx1_ASAP7_75t_L g588 ( .A(n_552), .Y(n_588) );
AND4x1_ASAP7_75t_L g552 ( .A(n_553), .B(n_563), .C(n_574), .D(n_582), .Y(n_552) );
INVx1_ASAP7_75t_L g841 ( .A(n_554), .Y(n_841) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_559), .B2(n_560), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_557), .A2(n_749), .B1(n_750), .B2(n_751), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_557), .A2(n_836), .B1(n_837), .B2(n_838), .Y(n_835) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OAI221xp5_ASAP7_75t_SL g760 ( .A1(n_560), .A2(n_761), .B1(n_762), .B2(n_764), .C(n_765), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_560), .A2(n_840), .B1(n_841), .B2(n_842), .Y(n_839) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g751 ( .A(n_561), .Y(n_751) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g1058 ( .A(n_565), .Y(n_1058) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_570), .B2(n_571), .Y(n_566) );
OAI21xp33_ASAP7_75t_L g809 ( .A1(n_568), .A2(n_810), .B(n_811), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_568), .A2(n_831), .B1(n_832), .B2(n_833), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g1060 ( .A1(n_568), .A2(n_1061), .B1(n_1062), .B2(n_1063), .Y(n_1060) );
BUFx2_ASAP7_75t_R g568 ( .A(n_569), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_572), .Y(n_571) );
BUFx4f_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_L g618 ( .A(n_573), .Y(n_618) );
BUFx2_ASAP7_75t_L g660 ( .A(n_573), .Y(n_660) );
BUFx2_ASAP7_75t_L g715 ( .A(n_573), .Y(n_715) );
BUFx2_ASAP7_75t_L g1064 ( .A(n_573), .Y(n_1064) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_579), .B1(n_580), .B2(n_581), .Y(n_577) );
INVx4_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx2_ASAP7_75t_L g595 ( .A(n_584), .Y(n_595) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_584), .A2(n_670), .B(n_671), .Y(n_669) );
OAI21xp5_ASAP7_75t_L g889 ( .A1(n_584), .A2(n_890), .B(n_891), .Y(n_889) );
OAI21xp5_ASAP7_75t_SL g983 ( .A1(n_584), .A2(n_984), .B(n_985), .Y(n_983) );
INVx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g687 ( .A(n_589), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_629), .B1(n_684), .B2(n_685), .Y(n_589) );
INVx1_ASAP7_75t_L g684 ( .A(n_590), .Y(n_684) );
INVx1_ASAP7_75t_L g628 ( .A(n_592), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_610), .C(n_619), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_604), .Y(n_593) );
OAI222xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_597), .B2(n_599), .C1(n_600), .C2(n_603), .Y(n_594) );
INVx1_ASAP7_75t_L g849 ( .A(n_595), .Y(n_849) );
OAI222xp33_ASAP7_75t_L g777 ( .A1(n_597), .A2(n_778), .B1(n_779), .B2(n_781), .C1(n_782), .C2(n_784), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_598), .Y(n_597) );
OAI222xp33_ASAP7_75t_L g1008 ( .A1(n_600), .A2(n_1009), .B1(n_1010), .B2(n_1011), .C1(n_1012), .C2(n_1013), .Y(n_1008) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
BUFx4f_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .Y(n_604) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_615), .Y(n_610) );
BUFx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVxp67_ASAP7_75t_L g833 ( .A(n_618), .Y(n_833) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_623), .Y(n_619) );
INVx2_ASAP7_75t_L g1168 ( .A(n_622), .Y(n_1168) );
INVx3_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx3_ASAP7_75t_L g654 ( .A(n_625), .Y(n_654) );
INVx1_ASAP7_75t_L g826 ( .A(n_626), .Y(n_826) );
BUFx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g685 ( .A(n_630), .Y(n_685) );
INVx2_ASAP7_75t_L g683 ( .A(n_631), .Y(n_683) );
XOR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_661), .Y(n_631) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_650), .Y(n_633) );
NOR3xp33_ASAP7_75t_L g634 ( .A(n_635), .B(n_640), .C(n_644), .Y(n_634) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g1083 ( .A(n_639), .Y(n_1083) );
OAI21xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B(n_643), .Y(n_640) );
OAI21xp33_ASAP7_75t_SL g734 ( .A1(n_642), .A2(n_735), .B(n_736), .Y(n_734) );
OAI21xp5_ASAP7_75t_SL g919 ( .A1(n_642), .A2(n_920), .B(n_921), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B1(n_647), .B2(n_648), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_648), .A2(n_845), .B1(n_846), .B2(n_847), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_648), .A2(n_847), .B1(n_1068), .B2(n_1069), .Y(n_1067) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx3_ASAP7_75t_SL g1089 ( .A(n_649), .Y(n_1089) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_655), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_659), .Y(n_655) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_658), .Y(n_766) );
INVx2_ASAP7_75t_L g814 ( .A(n_661), .Y(n_814) );
XOR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_682), .Y(n_661) );
NAND3x1_ASAP7_75t_L g662 ( .A(n_663), .B(n_668), .C(n_678), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_667), .Y(n_663) );
NOR2x1_ASAP7_75t_L g668 ( .A(n_669), .B(n_672), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .C(n_676), .Y(n_672) );
BUFx2_ASAP7_75t_L g1066 ( .A(n_674), .Y(n_1066) );
INVx1_ASAP7_75t_L g874 ( .A(n_677), .Y(n_874) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
XNOR2xp5_ASAP7_75t_SL g689 ( .A(n_690), .B(n_818), .Y(n_689) );
OAI22xp5_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_788), .B1(n_789), .B2(n_817), .Y(n_690) );
INVx2_ASAP7_75t_L g817 ( .A(n_691), .Y(n_817) );
AO22x2_ASAP7_75t_SL g691 ( .A1(n_692), .A2(n_693), .B1(n_757), .B2(n_787), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_721), .B2(n_722), .Y(n_693) );
INVx2_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND3x1_ASAP7_75t_L g698 ( .A(n_699), .B(n_710), .C(n_716), .Y(n_698) );
NOR3xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_704), .C(n_707), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_713), .Y(n_710) );
INVx1_ASAP7_75t_L g754 ( .A(n_712), .Y(n_754) );
HB1xp67_ASAP7_75t_L g1174 ( .A(n_712), .Y(n_1174) );
BUFx2_ASAP7_75t_L g1154 ( .A(n_714), .Y(n_1154) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
BUFx2_ASAP7_75t_L g804 ( .A(n_718), .Y(n_804) );
INVx1_ASAP7_75t_L g1053 ( .A(n_718), .Y(n_1053) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_726), .B(n_743), .Y(n_725) );
NOR3xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_734), .C(n_740), .Y(n_726) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_728), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g1080 ( .A1(n_730), .A2(n_1081), .B1(n_1082), .B2(n_1083), .Y(n_1080) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_730), .A2(n_1083), .B1(n_1150), .B2(n_1151), .Y(n_1149) );
INVx3_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NOR3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_748), .C(n_752), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B1(n_755), .B2(n_756), .Y(n_752) );
INVx1_ASAP7_75t_L g806 ( .A(n_756), .Y(n_806) );
INVx2_ASAP7_75t_L g787 ( .A(n_757), .Y(n_787) );
INVx1_ASAP7_75t_L g786 ( .A(n_758), .Y(n_786) );
AND2x2_ASAP7_75t_SL g758 ( .A(n_759), .B(n_771), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_768), .Y(n_759) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
NOR2xp33_ASAP7_75t_SL g771 ( .A(n_772), .B(n_777), .Y(n_771) );
OAI222xp33_ASAP7_75t_L g872 ( .A1(n_779), .A2(n_873), .B1(n_874), .B2(n_875), .C1(n_876), .C2(n_877), .Y(n_872) );
INVx2_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
INVx2_ASAP7_75t_L g794 ( .A(n_780), .Y(n_794) );
INVxp67_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
OAI22x1_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_814), .B1(n_815), .B2(n_816), .Y(n_789) );
INVx1_ASAP7_75t_L g815 ( .A(n_790), .Y(n_815) );
NAND3x1_ASAP7_75t_L g791 ( .A(n_792), .B(n_802), .C(n_807), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_799), .Y(n_792) );
OAI21xp5_ASAP7_75t_SL g793 ( .A1(n_794), .A2(n_795), .B(n_796), .Y(n_793) );
OAI21xp5_ASAP7_75t_SL g927 ( .A1(n_794), .A2(n_928), .B(n_929), .Y(n_927) );
INVx2_ASAP7_75t_SL g1009 ( .A(n_797), .Y(n_1009) );
BUFx6f_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
AND2x2_ASAP7_75t_L g802 ( .A(n_803), .B(n_805), .Y(n_802) );
INVx1_ASAP7_75t_L g816 ( .A(n_814), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_820), .B1(n_903), .B2(n_975), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_852), .B1(n_901), .B2(n_902), .Y(n_820) );
INVx1_ASAP7_75t_L g902 ( .A(n_821), .Y(n_902) );
INVx1_ASAP7_75t_L g851 ( .A(n_822), .Y(n_851) );
AND4x1_ASAP7_75t_L g822 ( .A(n_823), .B(n_834), .C(n_843), .D(n_848), .Y(n_822) );
NOR2xp33_ASAP7_75t_SL g823 ( .A(n_824), .B(n_830), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_826), .B1(n_827), .B2(n_828), .Y(n_824) );
INVxp67_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_835), .B(n_839), .Y(n_834) );
INVx2_ASAP7_75t_L g901 ( .A(n_852), .Y(n_901) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_853), .A2(n_854), .B1(n_883), .B2(n_900), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g882 ( .A(n_856), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_857), .B(n_871), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_858), .B(n_864), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
INVx2_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_867), .Y(n_864) );
INVx3_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_872), .B(n_878), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
INVx3_ASAP7_75t_L g900 ( .A(n_883), .Y(n_900) );
XOR2x2_ASAP7_75t_L g883 ( .A(n_884), .B(n_899), .Y(n_883) );
NAND3x1_ASAP7_75t_SL g884 ( .A(n_885), .B(n_888), .C(n_896), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
NOR2x1_ASAP7_75t_L g888 ( .A(n_889), .B(n_892), .Y(n_888) );
NAND3xp33_ASAP7_75t_L g892 ( .A(n_893), .B(n_894), .C(n_895), .Y(n_892) );
AND2x2_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
INVx2_ASAP7_75t_L g975 ( .A(n_903), .Y(n_975) );
BUFx3_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_906), .B1(n_950), .B2(n_951), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
AO22x1_ASAP7_75t_L g906 ( .A1(n_907), .A2(n_922), .B1(n_923), .B2(n_949), .Y(n_906) );
INVx1_ASAP7_75t_SL g949 ( .A(n_907), .Y(n_949) );
NOR4xp75_ASAP7_75t_L g908 ( .A(n_909), .B(n_912), .C(n_915), .D(n_919), .Y(n_908) );
NAND2xp5_ASAP7_75t_SL g909 ( .A(n_910), .B(n_911), .Y(n_909) );
NAND2xp5_ASAP7_75t_SL g912 ( .A(n_913), .B(n_914), .Y(n_912) );
NAND2xp5_ASAP7_75t_SL g915 ( .A(n_916), .B(n_917), .Y(n_915) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g948 ( .A(n_925), .Y(n_948) );
NAND3x1_ASAP7_75t_L g925 ( .A(n_926), .B(n_937), .C(n_944), .Y(n_925) );
NOR2x1_ASAP7_75t_L g926 ( .A(n_927), .B(n_930), .Y(n_926) );
NAND3xp33_ASAP7_75t_L g930 ( .A(n_931), .B(n_932), .C(n_933), .Y(n_930) );
INVx2_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
AND2x2_ASAP7_75t_L g937 ( .A(n_938), .B(n_941), .Y(n_937) );
INVx3_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
AND2x2_ASAP7_75t_L g944 ( .A(n_945), .B(n_947), .Y(n_944) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx1_ASAP7_75t_SL g974 ( .A(n_952), .Y(n_974) );
AND2x2_ASAP7_75t_L g952 ( .A(n_953), .B(n_964), .Y(n_952) );
NOR3xp33_ASAP7_75t_L g953 ( .A(n_954), .B(n_957), .C(n_961), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g964 ( .A(n_965), .B(n_970), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_966), .B(n_969), .Y(n_965) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx2_ASAP7_75t_L g1159 ( .A(n_968), .Y(n_1159) );
NAND2xp5_ASAP7_75t_SL g970 ( .A(n_971), .B(n_972), .Y(n_970) );
INVx1_ASAP7_75t_L g1121 ( .A(n_976), .Y(n_1121) );
AOI22xp5_ASAP7_75t_L g976 ( .A1(n_977), .A2(n_1048), .B1(n_1119), .B2(n_1120), .Y(n_976) );
INVx1_ASAP7_75t_L g1119 ( .A(n_977), .Y(n_1119) );
HB1xp67_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
AOI22xp5_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_1000), .B1(n_1046), .B2(n_1047), .Y(n_978) );
INVx2_ASAP7_75t_L g1047 ( .A(n_979), .Y(n_1047) );
HB1xp67_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
XOR2x2_ASAP7_75t_L g980 ( .A(n_981), .B(n_999), .Y(n_980) );
NAND3x1_ASAP7_75t_L g981 ( .A(n_982), .B(n_992), .C(n_996), .Y(n_981) );
NOR2x1_ASAP7_75t_L g982 ( .A(n_983), .B(n_986), .Y(n_982) );
NAND3xp33_ASAP7_75t_L g986 ( .A(n_987), .B(n_989), .C(n_990), .Y(n_986) );
AND2x2_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
AND2x2_ASAP7_75t_L g996 ( .A(n_997), .B(n_998), .Y(n_996) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1000), .Y(n_1046) );
AOI22xp5_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1025), .B1(n_1044), .B2(n_1045), .Y(n_1000) );
INVx2_ASAP7_75t_L g1044 ( .A(n_1001), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g1074 ( .A1(n_1001), .A2(n_1044), .B1(n_1075), .B2(n_1076), .Y(n_1074) );
XNOR2x2_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1003), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1017), .Y(n_1003) );
NOR3xp33_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1008), .C(n_1014), .Y(n_1004) );
OAI21xp5_ASAP7_75t_SL g1084 ( .A1(n_1011), .A2(n_1085), .B(n_1086), .Y(n_1084) );
NOR2xp33_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1022), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1021), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1024), .Y(n_1022) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1025), .Y(n_1045) );
INVx2_ASAP7_75t_L g1043 ( .A(n_1027), .Y(n_1043) );
NAND2x1_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1036), .Y(n_1027) );
NOR2xp33_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1033), .Y(n_1028) );
OAI21xp5_ASAP7_75t_SL g1029 ( .A1(n_1030), .A2(n_1031), .B(n_1032), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1035), .Y(n_1033) );
NOR2x1_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1040), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1039), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1042), .Y(n_1040) );
INVx2_ASAP7_75t_L g1120 ( .A(n_1048), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g1048 ( .A1(n_1049), .A2(n_1073), .B1(n_1117), .B2(n_1118), .Y(n_1048) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1049), .Y(n_1117) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1050), .Y(n_1072) );
AND4x2_ASAP7_75t_L g1050 ( .A(n_1051), .B(n_1059), .C(n_1065), .D(n_1070), .Y(n_1050) );
INVx2_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
OAI22xp5_ASAP7_75t_L g1054 ( .A1(n_1055), .A2(n_1056), .B1(n_1057), .B2(n_1058), .Y(n_1054) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx2_ASAP7_75t_L g1118 ( .A(n_1073), .Y(n_1118) );
BUFx2_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
AO22x1_ASAP7_75t_L g1076 ( .A1(n_1077), .A2(n_1100), .B1(n_1115), .B2(n_1116), .Y(n_1076) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1077), .Y(n_1115) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1078), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1091), .Y(n_1078) );
NOR3xp33_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1084), .C(n_1087), .Y(n_1079) );
OA211x2_ASAP7_75t_L g1105 ( .A1(n_1083), .A2(n_1106), .B(n_1107), .C(n_1108), .Y(n_1105) );
NOR2xp33_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1095), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1094), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1097), .Y(n_1095) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1100), .Y(n_1116) );
XOR2x2_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1114), .Y(n_1100) );
NAND4xp75_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1105), .C(n_1109), .D(n_1113), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1104), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1112), .Y(n_1109) );
INVx1_ASAP7_75t_SL g1123 ( .A(n_1124), .Y(n_1123) );
NOR2x1_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1129), .Y(n_1124) );
OR2x2_ASAP7_75t_SL g1192 ( .A(n_1125), .B(n_1130), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1128), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_1126), .B(n_1161), .Y(n_1160) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1127), .B(n_1161), .Y(n_1195) );
CKINVDCx16_ASAP7_75t_R g1161 ( .A(n_1128), .Y(n_1161) );
CKINVDCx20_ASAP7_75t_R g1129 ( .A(n_1130), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1132), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1135), .Y(n_1133) );
OAI222xp33_ASAP7_75t_L g1136 ( .A1(n_1137), .A2(n_1160), .B1(n_1162), .B2(n_1188), .C1(n_1190), .C2(n_1193), .Y(n_1136) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
NAND2x1_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1152), .Y(n_1139) );
NOR3xp33_ASAP7_75t_SL g1140 ( .A(n_1141), .B(n_1144), .C(n_1149), .Y(n_1140) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
AND4x1_ASAP7_75t_L g1152 ( .A(n_1153), .B(n_1155), .C(n_1156), .D(n_1158), .Y(n_1152) );
BUFx3_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1164), .Y(n_1189) );
AND2x2_ASAP7_75t_SL g1164 ( .A(n_1165), .B(n_1177), .Y(n_1164) );
NOR2xp33_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1171), .Y(n_1165) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
NOR3xp33_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1181), .C(n_1185), .Y(n_1177) );
CKINVDCx20_ASAP7_75t_R g1190 ( .A(n_1191), .Y(n_1190) );
CKINVDCx20_ASAP7_75t_R g1191 ( .A(n_1192), .Y(n_1191) );
CKINVDCx20_ASAP7_75t_R g1193 ( .A(n_1194), .Y(n_1193) );
endmodule