module fake_jpeg_12939_n_526 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_49),
.Y(n_149)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_15),
.B(n_13),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_59),
.B(n_85),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_66),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_18),
.B(n_12),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_93),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_81),
.Y(n_150)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_84),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_18),
.B(n_0),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_86),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_15),
.B(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_87),
.B(n_38),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_33),
.B(n_0),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_34),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_98),
.B(n_46),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_27),
.B1(n_37),
.B2(n_48),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_102),
.A2(n_110),
.B1(n_120),
.B2(n_123),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_51),
.A2(n_37),
.B1(n_48),
.B2(n_36),
.Y(n_109)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_109),
.A2(n_143),
.B(n_17),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_68),
.A2(n_27),
.B1(n_37),
.B2(n_48),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_116),
.B(n_29),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_56),
.A2(n_27),
.B1(n_37),
.B2(n_33),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_87),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_130),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_72),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_49),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_140),
.A2(n_16),
.B(n_17),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_51),
.A2(n_36),
.B1(n_46),
.B2(n_44),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_57),
.B(n_39),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_155),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_53),
.A2(n_36),
.B1(n_45),
.B2(n_29),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_24),
.B1(n_45),
.B2(n_43),
.Y(n_180)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_58),
.Y(n_153)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_57),
.B(n_43),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_96),
.Y(n_179)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_159),
.A2(n_180),
.B1(n_181),
.B2(n_151),
.Y(n_215)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_119),
.B(n_82),
.CI(n_80),
.CON(n_160),
.SN(n_160)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_160),
.B(n_175),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_99),
.B(n_28),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_161),
.B(n_186),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_176),
.Y(n_214)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_165),
.Y(n_242)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_40),
.B1(n_23),
.B2(n_44),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_168),
.A2(n_191),
.B1(n_112),
.B2(n_124),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_108),
.B(n_74),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_173),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_106),
.B(n_28),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_114),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

NAND2xp67_ASAP7_75t_SL g178 ( 
.A(n_118),
.B(n_41),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_SL g222 ( 
.A1(n_178),
.A2(n_149),
.B(n_156),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_179),
.B(n_185),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_109),
.A2(n_95),
.B1(n_89),
.B2(n_88),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_129),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_187),
.Y(n_221)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_184),
.Y(n_233)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_21),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_129),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_189),
.Y(n_224)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_154),
.A2(n_40),
.B1(n_23),
.B2(n_17),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_152),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_193),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_157),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_150),
.C(n_139),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_195),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_121),
.B(n_86),
.C(n_84),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_102),
.A2(n_78),
.B1(n_76),
.B2(n_69),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_64),
.B1(n_141),
.B2(n_131),
.Y(n_220)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_198),
.Y(n_229)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_110),
.B(n_41),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_202),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_125),
.B(n_24),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_201),
.Y(n_232)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_126),
.B(n_21),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_203),
.B(n_204),
.Y(n_243)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_207),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_126),
.B(n_16),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_206),
.B(n_143),
.Y(n_211)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_172),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_62),
.B1(n_67),
.B2(n_60),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_213),
.A2(n_215),
.B1(n_231),
.B2(n_236),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_160),
.A2(n_134),
.B1(n_151),
.B2(n_149),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_218),
.A2(n_220),
.B1(n_230),
.B2(n_245),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_222),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_159),
.A2(n_104),
.B1(n_131),
.B2(n_127),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_141),
.B1(n_113),
.B2(n_115),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_161),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_235),
.B(n_237),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_186),
.A2(n_124),
.B1(n_132),
.B2(n_103),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_202),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_199),
.A2(n_104),
.B1(n_115),
.B2(n_127),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_246),
.A2(n_275),
.B1(n_276),
.B2(n_220),
.Y(n_288)
);

NOR2x1p5_ASAP7_75t_SL g247 ( 
.A(n_211),
.B(n_208),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_260),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_248),
.B(n_240),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_223),
.B(n_208),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_249),
.A2(n_250),
.B(n_266),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_209),
.A2(n_160),
.B(n_178),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_218),
.A2(n_206),
.B1(n_173),
.B2(n_194),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_251),
.A2(n_263),
.B(n_268),
.Y(n_287)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_221),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_254),
.B(n_255),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_214),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_208),
.B(n_171),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_269),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_173),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_209),
.A2(n_179),
.B1(n_195),
.B2(n_163),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_225),
.Y(n_264)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_265),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_228),
.A2(n_176),
.B(n_188),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_244),
.A2(n_179),
.B(n_158),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_211),
.B(n_185),
.C(n_190),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_234),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_270),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_198),
.B(n_207),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_162),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_274),
.Y(n_300)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_225),
.Y(n_273)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_273),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_215),
.A2(n_117),
.B1(n_113),
.B2(n_162),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_215),
.A2(n_117),
.B1(n_170),
.B2(n_167),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_226),
.Y(n_277)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_277),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_230),
.A2(n_164),
.B1(n_189),
.B2(n_184),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_278),
.A2(n_231),
.B1(n_213),
.B2(n_233),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_214),
.B(n_166),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_279),
.B(n_238),
.Y(n_283)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_224),
.Y(n_280)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_283),
.Y(n_328)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_285),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_288),
.A2(n_302),
.B1(n_305),
.B2(n_261),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_279),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_289),
.B(n_293),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_290),
.A2(n_304),
.B1(n_270),
.B2(n_273),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_274),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_256),
.A2(n_217),
.B1(n_212),
.B2(n_219),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_296),
.A2(n_310),
.B(n_271),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_314),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_275),
.A2(n_276),
.B1(n_246),
.B2(n_262),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_303),
.B(n_239),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_261),
.A2(n_240),
.B1(n_241),
.B2(n_227),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_262),
.A2(n_245),
.B1(n_222),
.B2(n_241),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_267),
.B(n_280),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_306),
.B(n_308),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_249),
.B(n_232),
.Y(n_307)
);

AO21x1_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_250),
.B(n_247),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_232),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_252),
.A2(n_239),
.B1(n_227),
.B2(n_212),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_259),
.B(n_239),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_282),
.C(n_303),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_257),
.B(n_265),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_260),
.B(n_239),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_247),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_316),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_254),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_318),
.B(n_319),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_314),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_255),
.Y(n_320)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_320),
.Y(n_356)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_291),
.Y(n_322)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_322),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_323),
.A2(n_302),
.B1(n_288),
.B2(n_290),
.Y(n_357)
);

AO21x2_ASAP7_75t_L g324 ( 
.A1(n_300),
.A2(n_278),
.B(n_266),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_324),
.A2(n_347),
.B1(n_349),
.B2(n_350),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_306),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_325),
.B(n_326),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_308),
.B(n_248),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_330),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_329),
.A2(n_292),
.B(n_309),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_297),
.B(n_269),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_251),
.Y(n_331)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_331),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_332),
.B(n_333),
.C(n_210),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_282),
.B(n_263),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_291),
.Y(n_334)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_334),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_311),
.B(n_289),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_335),
.B(n_339),
.Y(n_360)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_294),
.Y(n_336)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_336),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_283),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_337),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_311),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_338),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_295),
.B(n_229),
.Y(n_340)
);

AO221x1_ASAP7_75t_L g353 ( 
.A1(n_340),
.A2(n_342),
.B1(n_345),
.B2(n_346),
.C(n_348),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_294),
.B(n_268),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_341),
.B(n_299),
.Y(n_363)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_301),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_295),
.B(n_229),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_301),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_284),
.B(n_277),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_307),
.A2(n_253),
.B1(n_270),
.B2(n_264),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_329),
.A2(n_309),
.B(n_307),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_351),
.A2(n_372),
.B(n_375),
.Y(n_396)
);

FAx1_ASAP7_75t_SL g354 ( 
.A(n_326),
.B(n_298),
.CI(n_315),
.CON(n_354),
.SN(n_354)
);

FAx1_ASAP7_75t_SL g393 ( 
.A(n_354),
.B(n_317),
.CI(n_337),
.CON(n_393),
.SN(n_393)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_355),
.A2(n_132),
.B(n_135),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_357),
.A2(n_384),
.B1(n_324),
.B2(n_382),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_323),
.A2(n_298),
.B1(n_287),
.B2(n_313),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_358),
.A2(n_361),
.B1(n_382),
.B2(n_324),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_319),
.A2(n_287),
.B1(n_310),
.B2(n_305),
.Y(n_361)
);

MAJx2_ASAP7_75t_L g397 ( 
.A(n_362),
.B(n_344),
.C(n_345),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_363),
.B(n_343),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_324),
.A2(n_299),
.B1(n_285),
.B2(n_281),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_365),
.A2(n_383),
.B1(n_322),
.B2(n_336),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_332),
.B(n_233),
.C(n_197),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_371),
.C(n_373),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_333),
.B(n_226),
.C(n_177),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_341),
.A2(n_312),
.B(n_212),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_330),
.B(n_201),
.C(n_234),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_331),
.A2(n_312),
.B(n_216),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_SL g376 ( 
.A(n_344),
.B(n_321),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_376),
.B(n_350),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_234),
.C(n_164),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_378),
.B(n_379),
.C(n_334),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_216),
.C(n_286),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_325),
.A2(n_281),
.B1(n_312),
.B2(n_219),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_324),
.A2(n_182),
.B1(n_203),
.B2(n_219),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_328),
.A2(n_242),
.B1(n_165),
.B2(n_204),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_374),
.Y(n_385)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_385),
.Y(n_423)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_374),
.Y(n_386)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_386),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_360),
.B(n_316),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_388),
.B(n_406),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_389),
.A2(n_398),
.B1(n_370),
.B2(n_384),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_362),
.B(n_316),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_390),
.B(n_408),
.Y(n_419)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_377),
.Y(n_391)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_391),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_397),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_393),
.B(n_409),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_369),
.B(n_335),
.C(n_321),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_394),
.B(n_399),
.C(n_400),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_317),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_395),
.B(n_403),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_347),
.C(n_342),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_346),
.C(n_349),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_401),
.A2(n_402),
.B1(n_404),
.B2(n_365),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_357),
.A2(n_361),
.B1(n_324),
.B2(n_358),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_368),
.B(n_348),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_368),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_405),
.B(n_363),
.Y(n_426)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_377),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_407),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_343),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_359),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_242),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_SL g416 ( 
.A(n_410),
.B(n_411),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_356),
.B(n_242),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_412),
.A2(n_355),
.B(n_372),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_380),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_413),
.Y(n_420)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_353),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_414),
.B(n_367),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_415),
.A2(n_421),
.B1(n_436),
.B2(n_1),
.Y(n_449)
);

FAx1_ASAP7_75t_SL g417 ( 
.A(n_393),
.B(n_354),
.CI(n_352),
.CON(n_417),
.SN(n_417)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_429),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_389),
.A2(n_395),
.B1(n_370),
.B2(n_352),
.Y(n_421)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_424),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_426),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_428),
.A2(n_403),
.B1(n_392),
.B2(n_393),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_387),
.B(n_378),
.C(n_373),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_390),
.B(n_351),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_432),
.B(n_438),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_394),
.B(n_375),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_435),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_396),
.A2(n_366),
.B1(n_383),
.B2(n_354),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_396),
.A2(n_360),
.B(n_105),
.Y(n_437)
);

MAJx2_ASAP7_75t_L g442 ( 
.A(n_437),
.B(n_410),
.C(n_399),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_397),
.B(n_0),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_418),
.Y(n_440)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_440),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_SL g441 ( 
.A1(n_436),
.A2(n_401),
.B1(n_402),
.B2(n_411),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_441),
.A2(n_446),
.B1(n_449),
.B2(n_452),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_442),
.B(n_448),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_418),
.B(n_400),
.Y(n_443)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_443),
.Y(n_475)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_444),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_425),
.C(n_387),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_451),
.C(n_453),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_439),
.A2(n_388),
.B1(n_412),
.B2(n_408),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_406),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_425),
.B(n_1),
.C(n_2),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_439),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_419),
.B(n_2),
.C(n_3),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_432),
.B(n_3),
.C(n_4),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_455),
.B(n_431),
.C(n_433),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_437),
.B(n_3),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_457),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_427),
.B(n_4),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_459),
.B(n_427),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_438),
.B(n_417),
.Y(n_460)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_460),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_461),
.B(n_465),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_458),
.B(n_420),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_464),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_450),
.A2(n_422),
.B(n_428),
.Y(n_464)
);

FAx1_ASAP7_75t_SL g466 ( 
.A(n_447),
.B(n_417),
.CI(n_416),
.CON(n_466),
.SN(n_466)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_467),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_456),
.B(n_433),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_435),
.C(n_430),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_471),
.B(n_472),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_453),
.B(n_430),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_451),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_473),
.B(n_477),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_452),
.B(n_423),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_448),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_487),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_470),
.A2(n_423),
.B1(n_455),
.B2(n_459),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_480),
.B(n_481),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_471),
.B(n_441),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_470),
.A2(n_468),
.B1(n_476),
.B2(n_474),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_491),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_475),
.B(n_454),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_484),
.B(n_485),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_468),
.B(n_442),
.C(n_446),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_469),
.B(n_4),
.Y(n_487)
);

A2O1A1Ixp33_ASAP7_75t_SL g489 ( 
.A1(n_466),
.A2(n_464),
.B(n_476),
.C(n_477),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_489),
.A2(n_472),
.B(n_465),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_463),
.B(n_5),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_5),
.C(n_6),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_7),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_462),
.B(n_5),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_494),
.Y(n_501)
);

OAI21xp33_ASAP7_75t_SL g496 ( 
.A1(n_488),
.A2(n_466),
.B(n_467),
.Y(n_496)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_496),
.Y(n_507)
);

NAND3xp33_ASAP7_75t_SL g514 ( 
.A(n_497),
.B(n_503),
.C(n_7),
.Y(n_514)
);

INVx11_ASAP7_75t_L g498 ( 
.A(n_489),
.Y(n_498)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_498),
.Y(n_512)
);

AOI21xp33_ASAP7_75t_L g502 ( 
.A1(n_482),
.A2(n_486),
.B(n_490),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_502),
.A2(n_497),
.B(n_498),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_489),
.A2(n_478),
.B(n_461),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_504),
.B(n_506),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_491),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_508),
.A2(n_509),
.B(n_510),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_500),
.A2(n_489),
.B(n_479),
.Y(n_509)
);

OAI21xp33_ASAP7_75t_L g510 ( 
.A1(n_503),
.A2(n_493),
.B(n_487),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_478),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_511),
.B(n_7),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_514),
.A2(n_501),
.B(n_499),
.Y(n_515)
);

NOR3xp33_ASAP7_75t_L g521 ( 
.A(n_515),
.B(n_516),
.C(n_518),
.Y(n_521)
);

OAI321xp33_ASAP7_75t_L g516 ( 
.A1(n_512),
.A2(n_507),
.A3(n_513),
.B1(n_514),
.B2(n_505),
.C(n_495),
.Y(n_516)
);

AO21x1_ASAP7_75t_L g517 ( 
.A1(n_512),
.A2(n_7),
.B(n_8),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_517),
.A2(n_8),
.B(n_9),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_519),
.A2(n_7),
.B(n_8),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_520),
.B(n_522),
.C(n_9),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_521),
.C(n_10),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_524),
.A2(n_10),
.B(n_11),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_10),
.Y(n_526)
);


endmodule