module real_aes_7636_n_207 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_174, n_156, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_183, n_205, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_3, n_41, n_140, n_153, n_75, n_178, n_19, n_71, n_180, n_40, n_49, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_81, n_133, n_48, n_204, n_37, n_117, n_97, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_207);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_97;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_207;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_216;
wire n_467;
wire n_327;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_532;
wire n_656;
wire n_316;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_504;
wire n_455;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_649;
wire n_293;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_498;
wire n_481;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_208;
wire n_215;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
wire n_237;
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_0), .A2(n_126), .B1(n_532), .B2(n_568), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_1), .A2(n_66), .B1(n_354), .B2(n_415), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_2), .A2(n_38), .B1(n_245), .B2(n_363), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_3), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_4), .Y(n_333) );
AOI22xp33_ASAP7_75t_SL g358 ( .A1(n_5), .A2(n_201), .B1(n_359), .B2(n_361), .Y(n_358) );
AOI22xp33_ASAP7_75t_SL g497 ( .A1(n_6), .A2(n_87), .B1(n_498), .B2(n_499), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_7), .A2(n_103), .B1(n_245), .B2(n_356), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_8), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_9), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_10), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_11), .A2(n_40), .B1(n_412), .B2(n_414), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_12), .A2(n_160), .B1(n_532), .B2(n_534), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g590 ( .A1(n_13), .A2(n_104), .B1(n_399), .B2(n_555), .Y(n_590) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_14), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_15), .A2(n_168), .B1(n_354), .B2(n_394), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_16), .A2(n_205), .B1(n_246), .B2(n_498), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g335 ( .A(n_17), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_18), .Y(n_462) );
AOI22x1_ASAP7_75t_L g221 ( .A1(n_19), .A2(n_222), .B1(n_327), .B2(n_328), .Y(n_221) );
INVx1_ASAP7_75t_L g327 ( .A(n_19), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_20), .A2(n_200), .B1(n_386), .B2(n_387), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_21), .Y(n_448) );
AO22x2_ASAP7_75t_L g239 ( .A1(n_22), .A2(n_80), .B1(n_231), .B2(n_236), .Y(n_239) );
INVx1_ASAP7_75t_L g669 ( .A(n_22), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_23), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_24), .A2(n_181), .B1(n_245), .B2(n_363), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_25), .A2(n_57), .B1(n_409), .B2(n_410), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_26), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_27), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_28), .A2(n_194), .B1(n_499), .B2(n_541), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_29), .A2(n_118), .B1(n_469), .B2(n_470), .Y(n_468) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_30), .A2(n_41), .B1(n_263), .B2(n_423), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_31), .A2(n_109), .B1(n_412), .B2(n_618), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g302 ( .A(n_32), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_33), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_34), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_35), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_36), .A2(n_89), .B1(n_375), .B2(n_568), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_37), .A2(n_128), .B1(n_246), .B2(n_504), .Y(n_503) );
AO22x2_ASAP7_75t_L g241 ( .A1(n_39), .A2(n_82), .B1(n_231), .B2(n_232), .Y(n_241) );
INVx1_ASAP7_75t_L g670 ( .A(n_39), .Y(n_670) );
INVx1_ASAP7_75t_L g426 ( .A(n_42), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_43), .A2(n_184), .B1(n_476), .B2(n_477), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_44), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_45), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_46), .B(n_382), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g645 ( .A1(n_47), .A2(n_151), .B1(n_351), .B2(n_354), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_48), .A2(n_157), .B1(n_274), .B2(n_618), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_49), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_50), .A2(n_78), .B1(n_252), .B2(n_351), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_51), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_52), .A2(n_94), .B1(n_226), .B2(n_256), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_53), .A2(n_172), .B1(n_310), .B2(n_399), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g691 ( .A1(n_54), .A2(n_175), .B1(n_359), .B2(n_361), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_55), .A2(n_106), .B1(n_250), .B2(n_255), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_56), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_58), .A2(n_135), .B1(n_387), .B2(n_494), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g347 ( .A(n_59), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_60), .A2(n_77), .B1(n_310), .B2(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_61), .A2(n_70), .B1(n_565), .B2(n_566), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_62), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_63), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_64), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_65), .A2(n_108), .B1(n_297), .B2(n_398), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_67), .A2(n_166), .B1(n_418), .B2(n_419), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_68), .A2(n_164), .B1(n_592), .B2(n_594), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g289 ( .A(n_69), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_71), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_72), .A2(n_88), .B1(n_277), .B2(n_422), .Y(n_421) );
AOI222xp33_ASAP7_75t_L g395 ( .A1(n_73), .A2(n_125), .B1(n_132), .B2(n_396), .C1(n_397), .C2(n_399), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_74), .A2(n_76), .B1(n_351), .B2(n_467), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_75), .A2(n_149), .B1(n_354), .B2(n_356), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_79), .A2(n_117), .B1(n_388), .B2(n_455), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_81), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_83), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_84), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g215 ( .A(n_85), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_86), .A2(n_191), .B1(n_473), .B2(n_474), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_90), .A2(n_150), .B1(n_273), .B2(n_277), .Y(n_272) );
INVx1_ASAP7_75t_L g213 ( .A(n_91), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_92), .A2(n_134), .B1(n_351), .B2(n_392), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_93), .A2(n_116), .B1(n_263), .B2(n_603), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_95), .A2(n_197), .B1(n_311), .B2(n_342), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_96), .A2(n_177), .B1(n_469), .B2(n_616), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_97), .A2(n_100), .B1(n_342), .B2(n_387), .Y(n_642) );
OA22x2_ASAP7_75t_L g630 ( .A1(n_98), .A2(n_631), .B1(n_632), .B2(n_651), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_98), .Y(n_631) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_99), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_101), .B(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_102), .B(n_593), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_105), .A2(n_107), .B1(n_374), .B2(n_375), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_110), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_111), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_112), .B(n_489), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_113), .A2(n_176), .B1(n_356), .B2(n_565), .Y(n_598) );
INVx2_ASAP7_75t_L g216 ( .A(n_114), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_115), .B(n_640), .Y(n_639) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_119), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_120), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_121), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_122), .Y(n_557) );
AND2x6_ASAP7_75t_L g212 ( .A(n_123), .B(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_123), .Y(n_663) );
AO22x2_ASAP7_75t_L g230 ( .A1(n_124), .A2(n_167), .B1(n_231), .B2(n_232), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_127), .A2(n_147), .B1(n_467), .B2(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_129), .B(n_491), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_130), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g678 ( .A(n_131), .Y(n_678) );
INVx1_ASAP7_75t_L g542 ( .A(n_133), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_136), .Y(n_514) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_137), .A2(n_192), .B1(n_246), .B2(n_356), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_138), .A2(n_146), .B1(n_388), .B2(n_637), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_139), .B(n_453), .Y(n_452) );
AOI22xp33_ASAP7_75t_SL g648 ( .A1(n_140), .A2(n_188), .B1(n_616), .B2(n_649), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_141), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_142), .A2(n_161), .B1(n_453), .B2(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_143), .A2(n_206), .B1(n_250), .B2(n_688), .Y(n_687) );
AO22x2_ASAP7_75t_L g235 ( .A1(n_144), .A2(n_183), .B1(n_231), .B2(n_236), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_145), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_148), .A2(n_405), .B1(n_440), .B2(n_441), .Y(n_404) );
INVx1_ASAP7_75t_L g440 ( .A(n_148), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g646 ( .A1(n_152), .A2(n_169), .B1(n_423), .B2(n_504), .Y(n_646) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_153), .A2(n_187), .B1(n_398), .B2(n_637), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_154), .A2(n_165), .B1(n_342), .B2(n_398), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_155), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_156), .Y(n_570) );
AOI211xp5_ASAP7_75t_L g207 ( .A1(n_158), .A2(n_208), .B(n_217), .C(n_671), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_159), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_162), .A2(n_190), .B1(n_470), .B2(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_163), .B(n_382), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_167), .B(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_170), .B(n_435), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_171), .Y(n_313) );
INVx1_ASAP7_75t_L g612 ( .A(n_173), .Y(n_612) );
INVx1_ASAP7_75t_L g364 ( .A(n_174), .Y(n_364) );
OA22x2_ASAP7_75t_L g578 ( .A1(n_178), .A2(n_579), .B1(n_580), .B2(n_604), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_178), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_179), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_180), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g283 ( .A(n_182), .Y(n_283) );
INVx1_ASAP7_75t_L g666 ( .A(n_183), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_185), .A2(n_195), .B1(n_351), .B2(n_541), .Y(n_540) );
AOI211xp5_ASAP7_75t_L g547 ( .A1(n_186), .A2(n_548), .B(n_549), .C(n_556), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_189), .A2(n_673), .B1(n_674), .B2(n_693), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_189), .Y(n_693) );
INVx1_ASAP7_75t_L g231 ( .A(n_193), .Y(n_231) );
INVx1_ASAP7_75t_L g233 ( .A(n_193), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_196), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_198), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_199), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_202), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g320 ( .A(n_203), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_204), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_209), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_210), .Y(n_209) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_212), .B(n_214), .Y(n_211) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_213), .Y(n_662) );
OAI21xp5_ASAP7_75t_L g699 ( .A1(n_214), .A2(n_661), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
AOI221xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_507), .B1(n_656), .B2(n_657), .C(n_658), .Y(n_217) );
INVx1_ASAP7_75t_L g656 ( .A(n_218), .Y(n_656) );
XOR2xp5_ASAP7_75t_L g218 ( .A(n_219), .B(n_366), .Y(n_218) );
OAI22xp5_ASAP7_75t_SL g219 ( .A1(n_220), .A2(n_221), .B1(n_329), .B2(n_365), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_SL g328 ( .A(n_222), .Y(n_328) );
AND2x2_ASAP7_75t_SL g222 ( .A(n_223), .B(n_281), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_260), .Y(n_223) );
OAI221xp5_ASAP7_75t_SL g224 ( .A1(n_225), .A2(n_242), .B1(n_243), .B2(n_248), .C(n_249), .Y(n_224) );
INVx2_ASAP7_75t_L g565 ( .A(n_225), .Y(n_565) );
INVx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
BUFx3_ASAP7_75t_L g418 ( .A(n_226), .Y(n_418) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g355 ( .A(n_227), .Y(n_355) );
BUFx2_ASAP7_75t_SL g530 ( .A(n_227), .Y(n_530) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_237), .Y(n_227) );
AND2x6_ASAP7_75t_L g252 ( .A(n_228), .B(n_253), .Y(n_252) );
AND2x4_ASAP7_75t_L g263 ( .A(n_228), .B(n_264), .Y(n_263) );
AND2x6_ASAP7_75t_L g305 ( .A(n_228), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_234), .Y(n_228) );
AND2x2_ASAP7_75t_L g247 ( .A(n_229), .B(n_235), .Y(n_247) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_230), .B(n_235), .Y(n_259) );
AND2x2_ASAP7_75t_L g269 ( .A(n_230), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g301 ( .A(n_230), .B(n_239), .Y(n_301) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g236 ( .A(n_233), .Y(n_236) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g270 ( .A(n_235), .Y(n_270) );
INVx1_ASAP7_75t_L g300 ( .A(n_235), .Y(n_300) );
AND2x4_ASAP7_75t_L g246 ( .A(n_237), .B(n_247), .Y(n_246) );
AND2x4_ASAP7_75t_L g257 ( .A(n_237), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_237), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g352 ( .A(n_237), .B(n_269), .Y(n_352) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_240), .Y(n_237) );
OR2x2_ASAP7_75t_L g254 ( .A(n_238), .B(n_241), .Y(n_254) );
AND2x2_ASAP7_75t_L g264 ( .A(n_238), .B(n_241), .Y(n_264) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g306 ( .A(n_239), .B(n_241), .Y(n_306) );
AND2x2_ASAP7_75t_L g299 ( .A(n_240), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g319 ( .A(n_240), .Y(n_319) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g280 ( .A(n_241), .Y(n_280) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g413 ( .A(n_246), .Y(n_413) );
BUFx3_ASAP7_75t_L g476 ( .A(n_246), .Y(n_476) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_246), .Y(n_539) );
INVx1_ASAP7_75t_L g288 ( .A(n_247), .Y(n_288) );
NAND2x1p5_ASAP7_75t_L g293 ( .A(n_247), .B(n_264), .Y(n_293) );
AND2x4_ASAP7_75t_L g384 ( .A(n_247), .B(n_253), .Y(n_384) );
AND2x6_ASAP7_75t_L g492 ( .A(n_247), .B(n_264), .Y(n_492) );
INVx4_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g392 ( .A(n_251), .Y(n_392) );
INVx5_ASAP7_75t_SL g498 ( .A(n_251), .Y(n_498) );
INVx11_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx11_ASAP7_75t_L g420 ( .A(n_252), .Y(n_420) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g287 ( .A(n_254), .B(n_288), .Y(n_287) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
BUFx2_ASAP7_75t_L g356 ( .A(n_257), .Y(n_356) );
BUFx3_ASAP7_75t_L g394 ( .A(n_257), .Y(n_394) );
BUFx3_ASAP7_75t_L g415 ( .A(n_257), .Y(n_415) );
BUFx2_ASAP7_75t_SL g470 ( .A(n_257), .Y(n_470) );
AND2x2_ASAP7_75t_L g618 ( .A(n_258), .B(n_319), .Y(n_618) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x6_ASAP7_75t_L g279 ( .A(n_259), .B(n_280), .Y(n_279) );
OAI221xp5_ASAP7_75t_SL g260 ( .A1(n_261), .A2(n_265), .B1(n_266), .B2(n_271), .C(n_272), .Y(n_260) );
INVx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx6_ASAP7_75t_L g360 ( .A(n_263), .Y(n_360) );
BUFx3_ASAP7_75t_L g409 ( .A(n_263), .Y(n_409) );
BUFx3_ASAP7_75t_L g541 ( .A(n_263), .Y(n_541) );
AND2x2_ASAP7_75t_L g276 ( .A(n_264), .B(n_269), .Y(n_276) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g573 ( .A(n_267), .Y(n_573) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g326 ( .A(n_270), .Y(n_326) );
BUFx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_274), .Y(n_474) );
INVx5_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx3_ASAP7_75t_L g361 ( .A(n_275), .Y(n_361) );
BUFx3_ASAP7_75t_L g376 ( .A(n_275), .Y(n_376) );
INVx4_ASAP7_75t_L g423 ( .A(n_275), .Y(n_423) );
INVx8_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
BUFx4f_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
BUFx2_ASAP7_75t_L g363 ( .A(n_278), .Y(n_363) );
BUFx2_ASAP7_75t_L g477 ( .A(n_278), .Y(n_477) );
INVx6_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_SL g504 ( .A(n_279), .Y(n_504) );
INVx1_ASAP7_75t_L g534 ( .A(n_279), .Y(n_534) );
INVx1_ASAP7_75t_SL g568 ( .A(n_279), .Y(n_568) );
INVx1_ASAP7_75t_L g389 ( .A(n_280), .Y(n_389) );
NOR3xp33_ASAP7_75t_L g281 ( .A(n_282), .B(n_294), .C(n_314), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B1(n_289), .B2(n_290), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_284), .A2(n_290), .B1(n_457), .B2(n_458), .Y(n_456) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx3_ASAP7_75t_L g334 ( .A(n_287), .Y(n_334) );
INVx2_ASAP7_75t_L g428 ( .A(n_287), .Y(n_428) );
OAI221xp5_ASAP7_75t_L g622 ( .A1(n_287), .A2(n_292), .B1(n_623), .B2(n_624), .C(n_625), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_290), .A2(n_514), .B1(n_515), .B2(n_516), .Y(n_513) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx3_ASAP7_75t_L g551 ( .A(n_292), .Y(n_551) );
BUFx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g337 ( .A(n_293), .Y(n_337) );
OAI222xp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_302), .B1(n_303), .B2(n_307), .C1(n_308), .C2(n_313), .Y(n_294) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_295), .A2(n_431), .B1(n_432), .B2(n_433), .C(n_434), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_295), .A2(n_557), .B1(n_558), .B2(n_559), .Y(n_556) );
INVx2_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_SL g346 ( .A(n_296), .Y(n_346) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g461 ( .A(n_297), .Y(n_461) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_298), .Y(n_386) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_298), .Y(n_494) );
BUFx4f_ASAP7_75t_SL g637 ( .A(n_298), .Y(n_637) );
AND2x4_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g312 ( .A(n_300), .Y(n_312) );
AND2x4_ASAP7_75t_L g311 ( .A(n_301), .B(n_312), .Y(n_311) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_301), .B(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g388 ( .A(n_301), .B(n_389), .Y(n_388) );
OAI222xp33_ASAP7_75t_L g582 ( .A1(n_303), .A2(n_583), .B1(n_584), .B2(n_585), .C1(n_586), .C2(n_588), .Y(n_582) );
INVx2_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g447 ( .A(n_304), .Y(n_447) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx4_ASAP7_75t_L g339 ( .A(n_305), .Y(n_339) );
INVx2_ASAP7_75t_SL g431 ( .A(n_305), .Y(n_431) );
INVx2_ASAP7_75t_L g484 ( .A(n_305), .Y(n_484) );
BUFx3_ASAP7_75t_L g548 ( .A(n_305), .Y(n_548) );
INVx1_ASAP7_75t_L g324 ( .A(n_306), .Y(n_324) );
AND2x4_ASAP7_75t_L g343 ( .A(n_306), .B(n_326), .Y(n_343) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g436 ( .A(n_310), .Y(n_436) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx12f_ASAP7_75t_L g398 ( .A(n_311), .Y(n_398) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_311), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B1(n_320), .B2(n_321), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_316), .A2(n_321), .B1(n_438), .B2(n_439), .Y(n_437) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx3_ASAP7_75t_SL g524 ( .A(n_317), .Y(n_524) );
INVx4_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_318), .A2(n_345), .B1(n_346), .B2(n_347), .Y(n_344) );
BUFx3_ASAP7_75t_L g463 ( .A(n_318), .Y(n_463) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g526 ( .A(n_322), .Y(n_526) );
CKINVDCx16_ASAP7_75t_R g322 ( .A(n_323), .Y(n_322) );
OR2x6_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g365 ( .A(n_329), .Y(n_365) );
XOR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_364), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_348), .Y(n_330) );
NOR3xp33_ASAP7_75t_L g331 ( .A(n_332), .B(n_338), .C(n_344), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_334), .B1(n_335), .B2(n_336), .Y(n_332) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g380 ( .A(n_337), .Y(n_380) );
OAI21xp5_ASAP7_75t_SL g338 ( .A1(n_339), .A2(n_340), .B(n_341), .Y(n_338) );
INVx4_ASAP7_75t_L g396 ( .A(n_339), .Y(n_396) );
BUFx2_ASAP7_75t_L g519 ( .A(n_339), .Y(n_519) );
BUFx2_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_SL g399 ( .A(n_343), .Y(n_399) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_343), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_357), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_353), .Y(n_349) );
BUFx2_ASAP7_75t_L g410 ( .A(n_351), .Y(n_410) );
BUFx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx3_ASAP7_75t_L g499 ( .A(n_352), .Y(n_499) );
BUFx3_ASAP7_75t_L g688 ( .A(n_352), .Y(n_688) );
INVx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx3_ASAP7_75t_L g469 ( .A(n_355), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_362), .Y(n_357) );
INVxp67_ASAP7_75t_L g571 ( .A(n_359), .Y(n_571) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g374 ( .A(n_360), .Y(n_374) );
INVx2_ASAP7_75t_L g473 ( .A(n_360), .Y(n_473) );
INVx3_ASAP7_75t_L g649 ( .A(n_360), .Y(n_649) );
AOI22xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_479), .B1(n_480), .B2(n_506), .Y(n_366) );
INVx1_ASAP7_75t_L g506 ( .A(n_367), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_369), .B1(n_401), .B2(n_402), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
XOR2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_400), .Y(n_370) );
NAND4xp75_ASAP7_75t_L g371 ( .A(n_372), .B(n_378), .C(n_390), .D(n_395), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_377), .Y(n_372) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OA211x2_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B(n_381), .C(n_385), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_380), .A2(n_426), .B1(n_427), .B2(n_429), .Y(n_425) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g489 ( .A(n_383), .Y(n_489) );
INVx5_ASAP7_75t_L g593 ( .A(n_383), .Y(n_593) );
INVx4_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx2_ASAP7_75t_L g555 ( .A(n_388), .Y(n_555) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
BUFx4f_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g561 ( .A(n_398), .Y(n_561) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI22xp5_ASAP7_75t_SL g402 ( .A1(n_403), .A2(n_404), .B1(n_442), .B2(n_443), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g441 ( .A(n_405), .Y(n_441) );
AND2x2_ASAP7_75t_SL g405 ( .A(n_406), .B(n_424), .Y(n_405) );
NOR2xp33_ASAP7_75t_SL g406 ( .A(n_407), .B(n_416), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_411), .Y(n_407) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_413), .A2(n_575), .B1(n_576), .B2(n_577), .Y(n_574) );
INVx1_ASAP7_75t_L g577 ( .A(n_414), .Y(n_577) );
BUFx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_421), .Y(n_416) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_SL g467 ( .A(n_420), .Y(n_467) );
INVx4_ASAP7_75t_L g616 ( .A(n_420), .Y(n_616) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g533 ( .A(n_423), .Y(n_533) );
NOR3xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_430), .C(n_437), .Y(n_424) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g515 ( .A(n_428), .Y(n_515) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
XOR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_478), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_464), .Y(n_444) );
NOR3xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_456), .C(n_459), .Y(n_445) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B1(n_449), .B2(n_451), .C(n_452), .Y(n_446) );
OAI21xp5_ASAP7_75t_L g677 ( .A1(n_447), .A2(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx4f_ASAP7_75t_L g587 ( .A(n_450), .Y(n_587) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_462), .B2(n_463), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_471), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_475), .Y(n_471) );
INVx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
XOR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_505), .Y(n_480) );
NAND2x1_ASAP7_75t_SL g481 ( .A(n_482), .B(n_495), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_487), .Y(n_482) );
OAI21xp5_ASAP7_75t_SL g483 ( .A1(n_484), .A2(n_485), .B(n_486), .Y(n_483) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_490), .C(n_493), .Y(n_487) );
BUFx2_ASAP7_75t_L g553 ( .A(n_489), .Y(n_553) );
BUFx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_SL g595 ( .A(n_492), .Y(n_595) );
BUFx4f_ASAP7_75t_L g683 ( .A(n_492), .Y(n_683) );
BUFx2_ASAP7_75t_L g521 ( .A(n_494), .Y(n_521) );
INVx2_ASAP7_75t_L g583 ( .A(n_494), .Y(n_583) );
NOR2x1_ASAP7_75t_L g495 ( .A(n_496), .B(n_501), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_500), .Y(n_496) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_498), .Y(n_566) );
BUFx3_ASAP7_75t_L g603 ( .A(n_499), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g657 ( .A(n_507), .Y(n_657) );
AOI22xp5_ASAP7_75t_SL g507 ( .A1(n_508), .A2(n_609), .B1(n_654), .B2(n_655), .Y(n_507) );
INVx1_ASAP7_75t_L g654 ( .A(n_508), .Y(n_654) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_543), .B1(n_607), .B2(n_608), .Y(n_509) );
INVx1_ASAP7_75t_L g607 ( .A(n_510), .Y(n_607) );
XOR2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_542), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_527), .Y(n_511) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_517), .C(n_522), .Y(n_512) );
OAI21xp33_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_520), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B1(n_525), .B2(n_526), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_528), .B(n_535), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_540), .Y(n_535) );
INVx4_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx4_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g608 ( .A(n_543), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_578), .B1(n_605), .B2(n_606), .Y(n_543) );
INVx2_ASAP7_75t_L g606 ( .A(n_544), .Y(n_606) );
XNOR2x1_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_562), .Y(n_546) );
INVx3_ASAP7_75t_L g627 ( .A(n_548), .Y(n_627) );
OAI211xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_551), .B(n_552), .C(n_554), .Y(n_549) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NOR3xp33_ASAP7_75t_L g562 ( .A(n_563), .B(n_569), .C(n_574), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_567), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_571), .B1(n_572), .B2(n_573), .Y(n_569) );
INVx1_ASAP7_75t_L g605 ( .A(n_578), .Y(n_605) );
INVx1_ASAP7_75t_SL g604 ( .A(n_580), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_596), .Y(n_580) );
NOR2x1_ASAP7_75t_L g581 ( .A(n_582), .B(n_589), .Y(n_581) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_SL g640 ( .A(n_595), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_600), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g655 ( .A(n_609), .Y(n_655) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_630), .B1(n_652), .B2(n_653), .Y(n_610) );
INVx2_ASAP7_75t_SL g652 ( .A(n_611), .Y(n_652) );
XNOR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
NOR4xp75_ASAP7_75t_L g613 ( .A(n_614), .B(n_619), .C(n_622), .D(n_626), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_615), .B(n_617), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_620), .B(n_621), .Y(n_619) );
OAI21xp5_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_628), .B(n_629), .Y(n_626) );
OAI21xp5_ASAP7_75t_SL g634 ( .A1(n_627), .A2(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g653 ( .A(n_630), .Y(n_653) );
INVx1_ASAP7_75t_L g651 ( .A(n_632), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_643), .Y(n_632) );
NOR2xp67_ASAP7_75t_L g633 ( .A(n_634), .B(n_638), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .C(n_642), .Y(n_638) );
NOR2x1_ASAP7_75t_L g643 ( .A(n_644), .B(n_647), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
NOR2x1_ASAP7_75t_L g659 ( .A(n_660), .B(n_664), .Y(n_659) );
OR2x2_ASAP7_75t_SL g705 ( .A(n_660), .B(n_665), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_662), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_662), .B(n_697), .Y(n_700) );
CKINVDCx16_ASAP7_75t_R g697 ( .A(n_663), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
OAI322xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_694), .A3(n_695), .B1(n_698), .B2(n_701), .C1(n_702), .C2(n_705), .Y(n_671) );
CKINVDCx16_ASAP7_75t_R g673 ( .A(n_674), .Y(n_673) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
XOR2x2_ASAP7_75t_L g704 ( .A(n_675), .B(n_701), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_676), .B(n_685), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_680), .Y(n_676) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .C(n_684), .Y(n_680) );
NOR2x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_690), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_689), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
CKINVDCx16_ASAP7_75t_R g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx3_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
endmodule