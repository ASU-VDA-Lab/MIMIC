module real_aes_539_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g501 ( .A(n_0), .B(n_193), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_1), .B(n_784), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_2), .Y(n_802) );
INVx1_ASAP7_75t_L g127 ( .A(n_3), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_4), .B(n_504), .Y(n_523) );
NAND2xp33_ASAP7_75t_SL g494 ( .A(n_5), .B(n_148), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_6), .B(n_161), .Y(n_184) );
INVx1_ASAP7_75t_L g486 ( .A(n_7), .Y(n_486) );
INVx1_ASAP7_75t_L g218 ( .A(n_8), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g784 ( .A(n_9), .Y(n_784) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_10), .Y(n_235) );
AND2x2_ASAP7_75t_L g521 ( .A(n_11), .B(n_117), .Y(n_521) );
INVx2_ASAP7_75t_L g118 ( .A(n_12), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g472 ( .A(n_13), .Y(n_472) );
INVx1_ASAP7_75t_L g194 ( .A(n_14), .Y(n_194) );
AOI221x1_ASAP7_75t_L g489 ( .A1(n_15), .A2(n_150), .B1(n_490), .B2(n_492), .C(n_493), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_16), .B(n_504), .Y(n_557) );
INVx1_ASAP7_75t_L g475 ( .A(n_17), .Y(n_475) );
INVx1_ASAP7_75t_L g191 ( .A(n_18), .Y(n_191) );
INVx1_ASAP7_75t_SL g139 ( .A(n_19), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_20), .B(n_142), .Y(n_164) );
AOI33xp33_ASAP7_75t_L g209 ( .A1(n_21), .A2(n_49), .A3(n_124), .B1(n_135), .B2(n_210), .B3(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_22), .A2(n_492), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_23), .B(n_193), .Y(n_526) );
AOI221xp5_ASAP7_75t_SL g566 ( .A1(n_24), .A2(n_39), .B1(n_492), .B2(n_504), .C(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g228 ( .A(n_25), .Y(n_228) );
OR2x2_ASAP7_75t_L g119 ( .A(n_26), .B(n_87), .Y(n_119) );
OA21x2_ASAP7_75t_L g152 ( .A1(n_26), .A2(n_87), .B(n_118), .Y(n_152) );
INVxp67_ASAP7_75t_L g488 ( .A(n_27), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_28), .B(n_196), .Y(n_561) );
AND2x2_ASAP7_75t_L g515 ( .A(n_29), .B(n_116), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_30), .B(n_122), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_31), .A2(n_492), .B(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_32), .B(n_196), .Y(n_568) );
AND2x2_ASAP7_75t_L g129 ( .A(n_33), .B(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g134 ( .A(n_33), .Y(n_134) );
AND2x2_ASAP7_75t_L g148 ( .A(n_33), .B(n_127), .Y(n_148) );
OR2x6_ASAP7_75t_L g473 ( .A(n_34), .B(n_474), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_35), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_36), .B(n_122), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g156 ( .A1(n_37), .A2(n_151), .B1(n_157), .B2(n_161), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_38), .B(n_166), .Y(n_165) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_40), .A2(n_79), .B1(n_132), .B2(n_492), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_41), .B(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_42), .B(n_193), .Y(n_513) );
AOI22xp33_ASAP7_75t_SL g770 ( .A1(n_43), .A2(n_769), .B1(n_771), .B2(n_773), .Y(n_770) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_44), .B(n_168), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_45), .B(n_142), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_46), .Y(n_160) );
AND2x2_ASAP7_75t_L g505 ( .A(n_47), .B(n_116), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_48), .B(n_116), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_50), .B(n_142), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_51), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_51), .A2(n_61), .B1(n_407), .B2(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g125 ( .A(n_52), .Y(n_125) );
INVx1_ASAP7_75t_L g144 ( .A(n_52), .Y(n_144) );
AND2x2_ASAP7_75t_L g260 ( .A(n_53), .B(n_116), .Y(n_260) );
AOI221xp5_ASAP7_75t_L g216 ( .A1(n_54), .A2(n_72), .B1(n_122), .B2(n_132), .C(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_55), .B(n_122), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_56), .B(n_504), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_57), .B(n_151), .Y(n_237) );
AOI21xp5_ASAP7_75t_SL g173 ( .A1(n_58), .A2(n_132), .B(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g542 ( .A(n_59), .B(n_116), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_60), .B(n_196), .Y(n_502) );
AOI222xp33_ASAP7_75t_L g99 ( .A1(n_61), .A2(n_100), .B1(n_777), .B2(n_788), .C1(n_803), .C2(n_805), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_61), .Y(n_799) );
INVx1_ASAP7_75t_L g187 ( .A(n_62), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_63), .B(n_193), .Y(n_540) );
AND2x2_ASAP7_75t_SL g562 ( .A(n_64), .B(n_117), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_65), .A2(n_492), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g258 ( .A(n_66), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_67), .B(n_196), .Y(n_527) );
AND2x2_ASAP7_75t_SL g534 ( .A(n_68), .B(n_168), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_69), .A2(n_132), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g130 ( .A(n_70), .Y(n_130) );
INVx1_ASAP7_75t_L g146 ( .A(n_70), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_71), .B(n_122), .Y(n_212) );
AND2x2_ASAP7_75t_L g149 ( .A(n_73), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g188 ( .A(n_74), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_75), .A2(n_132), .B(n_138), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g162 ( .A1(n_76), .A2(n_132), .B(n_163), .C(n_167), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_77), .A2(n_82), .B1(n_122), .B2(n_504), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_78), .B(n_504), .Y(n_541) );
INVx1_ASAP7_75t_L g476 ( .A(n_80), .Y(n_476) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_81), .B(n_150), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_83), .A2(n_132), .B1(n_207), .B2(n_208), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_84), .B(n_193), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_85), .B(n_193), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_86), .A2(n_492), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g175 ( .A(n_88), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_89), .B(n_196), .Y(n_539) );
AND2x2_ASAP7_75t_L g213 ( .A(n_90), .B(n_150), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_91), .A2(n_226), .B(n_227), .C(n_229), .Y(n_225) );
INVxp67_ASAP7_75t_L g491 ( .A(n_92), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_93), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_94), .B(n_196), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_95), .A2(n_492), .B(n_559), .Y(n_558) );
BUFx2_ASAP7_75t_L g785 ( .A(n_96), .Y(n_785) );
BUFx2_ASAP7_75t_SL g809 ( .A(n_96), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_97), .B(n_142), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_98), .Y(n_769) );
HB1xp67_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OAI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_769), .B(n_770), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OAI22x1_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_470), .B1(n_477), .B2(n_765), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_105), .A2(n_470), .B1(n_478), .B2(n_772), .Y(n_771) );
AND3x1_ASAP7_75t_L g105 ( .A(n_106), .B(n_464), .C(n_467), .Y(n_105) );
NAND5xp2_ASAP7_75t_L g106 ( .A(n_107), .B(n_364), .C(n_394), .D(n_408), .E(n_434), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OAI21xp33_ASAP7_75t_L g464 ( .A1(n_108), .A2(n_407), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g795 ( .A(n_108), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_313), .Y(n_108) );
NOR3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_261), .C(n_295), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_178), .B(n_200), .C(n_239), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_153), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_113), .B(n_251), .Y(n_316) );
AND2x2_ASAP7_75t_L g403 ( .A(n_113), .B(n_181), .Y(n_403) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OR2x2_ASAP7_75t_L g199 ( .A(n_114), .B(n_170), .Y(n_199) );
INVx1_ASAP7_75t_L g241 ( .A(n_114), .Y(n_241) );
INVx2_ASAP7_75t_L g246 ( .A(n_114), .Y(n_246) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_114), .Y(n_274) );
INVx1_ASAP7_75t_L g288 ( .A(n_114), .Y(n_288) );
AND2x2_ASAP7_75t_L g292 ( .A(n_114), .B(n_183), .Y(n_292) );
AND2x2_ASAP7_75t_L g373 ( .A(n_114), .B(n_182), .Y(n_373) );
AO21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_149), .Y(n_114) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_115), .A2(n_509), .B(n_515), .Y(n_508) );
AO21x2_ASAP7_75t_L g535 ( .A1(n_115), .A2(n_536), .B(n_542), .Y(n_535) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_115), .A2(n_509), .B(n_515), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
OA21x2_ASAP7_75t_L g565 ( .A1(n_116), .A2(n_566), .B(n_570), .Y(n_565) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_SL g117 ( .A(n_118), .B(n_119), .Y(n_117) );
AND2x4_ASAP7_75t_L g161 ( .A(n_118), .B(n_119), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_131), .Y(n_120) );
INVx1_ASAP7_75t_L g238 ( .A(n_122), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_122), .A2(n_132), .B1(n_485), .B2(n_487), .Y(n_484) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_128), .Y(n_122) );
INVx1_ASAP7_75t_L g158 ( .A(n_123), .Y(n_158) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
OR2x6_ASAP7_75t_L g140 ( .A(n_124), .B(n_136), .Y(n_140) );
INVxp33_ASAP7_75t_L g210 ( .A(n_124), .Y(n_210) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g137 ( .A(n_125), .B(n_127), .Y(n_137) );
AND2x4_ASAP7_75t_L g196 ( .A(n_125), .B(n_145), .Y(n_196) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g159 ( .A(n_128), .Y(n_159) );
BUFx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x6_ASAP7_75t_L g492 ( .A(n_129), .B(n_137), .Y(n_492) );
INVx2_ASAP7_75t_L g136 ( .A(n_130), .Y(n_136) );
AND2x6_ASAP7_75t_L g193 ( .A(n_130), .B(n_143), .Y(n_193) );
INVxp67_ASAP7_75t_L g236 ( .A(n_132), .Y(n_236) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
NOR2x1p5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
INVx1_ASAP7_75t_L g211 ( .A(n_135), .Y(n_211) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
O2A1O1Ixp33_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_140), .B(n_141), .C(n_147), .Y(n_138) );
INVx2_ASAP7_75t_L g166 ( .A(n_140), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_140), .A2(n_147), .B(n_175), .C(n_176), .Y(n_174) );
OAI22xp5_ASAP7_75t_L g186 ( .A1(n_140), .A2(n_187), .B1(n_188), .B2(n_189), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_SL g217 ( .A1(n_140), .A2(n_147), .B(n_218), .C(n_219), .Y(n_217) );
INVxp67_ASAP7_75t_L g226 ( .A(n_140), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_140), .A2(n_147), .B(n_258), .C(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g189 ( .A(n_142), .Y(n_189) );
AND2x4_ASAP7_75t_L g504 ( .A(n_142), .B(n_148), .Y(n_504) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_147), .A2(n_164), .B(n_165), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_147), .B(n_161), .Y(n_197) );
INVx1_ASAP7_75t_L g207 ( .A(n_147), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_147), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_147), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_147), .A2(n_526), .B(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_147), .A2(n_539), .B(n_540), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_147), .A2(n_560), .B(n_561), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_147), .A2(n_568), .B(n_569), .Y(n_567) );
INVx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_148), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g224 ( .A1(n_150), .A2(n_225), .B1(n_230), .B2(n_231), .Y(n_224) );
INVx3_ASAP7_75t_L g231 ( .A(n_150), .Y(n_231) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_151), .B(n_234), .Y(n_233) );
AOI21x1_ASAP7_75t_L g497 ( .A1(n_151), .A2(n_498), .B(n_505), .Y(n_497) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx4f_ASAP7_75t_L g168 ( .A(n_152), .Y(n_168) );
AND2x4_ASAP7_75t_SL g153 ( .A(n_154), .B(n_169), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g198 ( .A(n_155), .Y(n_198) );
AND2x2_ASAP7_75t_L g242 ( .A(n_155), .B(n_183), .Y(n_242) );
AND2x2_ASAP7_75t_L g263 ( .A(n_155), .B(n_170), .Y(n_263) );
INVx1_ASAP7_75t_L g286 ( .A(n_155), .Y(n_286) );
AND2x4_ASAP7_75t_L g353 ( .A(n_155), .B(n_182), .Y(n_353) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_162), .Y(n_155) );
NOR3xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .C(n_160), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_161), .A2(n_173), .B(n_177), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_161), .B(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_161), .B(n_488), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_161), .B(n_491), .Y(n_490) );
NOR3xp33_ASAP7_75t_L g493 ( .A(n_161), .B(n_189), .C(n_494), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_161), .A2(n_523), .B(n_524), .Y(n_522) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_167), .A2(n_205), .B(n_213), .Y(n_204) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_167), .A2(n_205), .B(n_213), .Y(n_268) );
AOI21x1_ASAP7_75t_L g530 ( .A1(n_167), .A2(n_531), .B(n_534), .Y(n_530) );
INVx2_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_168), .A2(n_216), .B(n_220), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_168), .A2(n_557), .B(n_558), .Y(n_556) );
AND2x4_ASAP7_75t_L g369 ( .A(n_169), .B(n_286), .Y(n_369) );
OR2x2_ASAP7_75t_L g410 ( .A(n_169), .B(n_411), .Y(n_410) );
NOR2xp67_ASAP7_75t_SL g429 ( .A(n_169), .B(n_302), .Y(n_429) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_169), .B(n_361), .Y(n_447) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2x1_ASAP7_75t_SL g247 ( .A(n_170), .B(n_183), .Y(n_247) );
AND2x4_ASAP7_75t_L g285 ( .A(n_170), .B(n_286), .Y(n_285) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_170), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_170), .B(n_245), .Y(n_323) );
INVx2_ASAP7_75t_L g337 ( .A(n_170), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_170), .B(n_289), .Y(n_359) );
AND2x2_ASAP7_75t_L g451 ( .A(n_170), .B(n_309), .Y(n_451) );
OR2x6_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2x1_ASAP7_75t_L g179 ( .A(n_180), .B(n_199), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_181), .B(n_288), .Y(n_302) );
AND2x2_ASAP7_75t_SL g311 ( .A(n_181), .B(n_291), .Y(n_311) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_198), .Y(n_181) );
INVx1_ASAP7_75t_L g289 ( .A(n_182), .Y(n_289) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g309 ( .A(n_183), .Y(n_309) );
AND2x4_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_190), .B(n_197), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_189), .B(n_228), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B1(n_194), .B2(n_195), .Y(n_190) );
INVxp67_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVxp67_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g342 ( .A(n_198), .Y(n_342) );
INVx2_ASAP7_75t_SL g387 ( .A(n_199), .Y(n_387) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_221), .Y(n_201) );
NAND2x1p5_ASAP7_75t_L g296 ( .A(n_202), .B(n_297), .Y(n_296) );
BUFx2_ASAP7_75t_L g333 ( .A(n_202), .Y(n_333) );
AND2x2_ASAP7_75t_L g457 ( .A(n_202), .B(n_282), .Y(n_457) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_214), .Y(n_202) );
AND2x4_ASAP7_75t_L g270 ( .A(n_203), .B(n_252), .Y(n_270) );
INVx1_ASAP7_75t_L g281 ( .A(n_203), .Y(n_281) );
AND2x2_ASAP7_75t_L g312 ( .A(n_203), .B(n_267), .Y(n_312) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_204), .B(n_215), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_204), .B(n_253), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_206), .B(n_212), .Y(n_205) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVxp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g250 ( .A(n_215), .Y(n_250) );
AND2x4_ASAP7_75t_L g318 ( .A(n_215), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g330 ( .A(n_215), .Y(n_330) );
INVx1_ASAP7_75t_L g372 ( .A(n_215), .Y(n_372) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_215), .Y(n_384) );
AND2x2_ASAP7_75t_L g400 ( .A(n_215), .B(n_223), .Y(n_400) );
BUFx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g347 ( .A(n_222), .B(n_305), .Y(n_347) );
INVx1_ASAP7_75t_SL g349 ( .A(n_222), .Y(n_349) );
AND2x2_ASAP7_75t_L g370 ( .A(n_222), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x4_ASAP7_75t_L g249 ( .A(n_223), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g277 ( .A(n_223), .Y(n_277) );
INVx2_ASAP7_75t_L g283 ( .A(n_223), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_223), .B(n_253), .Y(n_298) );
OR2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_232), .Y(n_223) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_231), .A2(n_254), .B(n_260), .Y(n_253) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_231), .A2(n_254), .B(n_260), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_236), .B1(n_237), .B2(n_238), .Y(n_232) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_243), .B(n_248), .Y(n_239) );
INVx1_ASAP7_75t_L g379 ( .A(n_240), .Y(n_379) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g299 ( .A(n_242), .Y(n_299) );
AND2x2_ASAP7_75t_L g355 ( .A(n_242), .B(n_291), .Y(n_355) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_247), .Y(n_243) );
INVx1_ASAP7_75t_L g269 ( .A(n_244), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_244), .B(n_285), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_244), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g376 ( .A(n_244), .B(n_369), .Y(n_376) );
AND2x2_ASAP7_75t_L g450 ( .A(n_244), .B(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_245), .Y(n_438) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_246), .Y(n_358) );
AND2x2_ASAP7_75t_L g271 ( .A(n_247), .B(n_272), .Y(n_271) );
OAI21xp33_ASAP7_75t_L g459 ( .A1(n_247), .A2(n_460), .B(n_462), .Y(n_459) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
INVx3_ASAP7_75t_L g345 ( .A(n_249), .Y(n_345) );
NAND2x1_ASAP7_75t_SL g389 ( .A(n_249), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g392 ( .A(n_249), .B(n_270), .Y(n_392) );
AND2x2_ASAP7_75t_L g304 ( .A(n_251), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g441 ( .A(n_251), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g452 ( .A(n_251), .B(n_400), .Y(n_452) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2x1p5_ASAP7_75t_L g328 ( .A(n_252), .B(n_329), .Y(n_328) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g383 ( .A(n_253), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
OAI21xp5_ASAP7_75t_SL g261 ( .A1(n_262), .A2(n_275), .B(n_278), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_264), .B1(n_270), .B2(n_271), .Y(n_262) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_263), .Y(n_320) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_269), .Y(n_264) );
AND2x2_ASAP7_75t_L g293 ( .A(n_265), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g399 ( .A(n_265), .B(n_400), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_265), .A2(n_418), .B1(n_419), .B2(n_420), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_265), .B(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g282 ( .A(n_267), .B(n_283), .Y(n_282) );
NOR2xp67_ASAP7_75t_L g363 ( .A(n_267), .B(n_283), .Y(n_363) );
NOR2x1_ASAP7_75t_L g371 ( .A(n_267), .B(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g319 ( .A(n_268), .Y(n_319) );
AND2x2_ASAP7_75t_L g327 ( .A(n_268), .B(n_283), .Y(n_327) );
INVx1_ASAP7_75t_L g390 ( .A(n_268), .Y(n_390) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2x1_ASAP7_75t_L g308 ( .A(n_273), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g420 ( .A(n_276), .B(n_305), .Y(n_420) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g294 ( .A(n_277), .Y(n_294) );
AND2x2_ASAP7_75t_L g317 ( .A(n_277), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g405 ( .A(n_277), .B(n_312), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_284), .B1(n_290), .B2(n_293), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g413 ( .A(n_280), .B(n_414), .Y(n_413) );
NAND2x1p5_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x2_ASAP7_75t_L g443 ( .A(n_283), .B(n_330), .Y(n_443) );
AND2x2_ASAP7_75t_SL g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx2_ASAP7_75t_L g310 ( .A(n_285), .Y(n_310) );
OAI21xp33_ASAP7_75t_SL g456 ( .A1(n_285), .A2(n_457), .B(n_458), .Y(n_456) );
AND2x4_ASAP7_75t_SL g287 ( .A(n_288), .B(n_289), .Y(n_287) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_288), .Y(n_446) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_SL g388 ( .A1(n_291), .A2(n_389), .B(n_391), .C(n_393), .Y(n_388) );
AND2x2_ASAP7_75t_SL g340 ( .A(n_292), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g393 ( .A(n_292), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_292), .B(n_369), .Y(n_433) );
INVx1_ASAP7_75t_SL g300 ( .A(n_293), .Y(n_300) );
AND2x2_ASAP7_75t_L g381 ( .A(n_294), .B(n_318), .Y(n_381) );
INVx1_ASAP7_75t_L g426 ( .A(n_294), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_299), .B1(n_300), .B2(n_301), .C(n_303), .Y(n_295) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_296), .Y(n_415) );
INVx2_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g463 ( .A(n_298), .B(n_306), .Y(n_463) );
OR2x2_ASAP7_75t_L g322 ( .A(n_299), .B(n_323), .Y(n_322) );
NOR2x1_ASAP7_75t_L g335 ( .A(n_299), .B(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_299), .B(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g461 ( .A(n_299), .B(n_358), .Y(n_461) );
BUFx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AOI32xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_307), .A3(n_310), .B1(n_311), .B2(n_312), .Y(n_303) );
INVx1_ASAP7_75t_L g324 ( .A(n_305), .Y(n_324) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_307), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g419 ( .A(n_308), .Y(n_419) );
OAI22xp33_ASAP7_75t_SL g401 ( .A1(n_310), .A2(n_402), .B1(n_404), .B2(n_406), .Y(n_401) );
INVx1_ASAP7_75t_L g432 ( .A(n_311), .Y(n_432) );
AOI211x1_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_320), .B(n_321), .C(n_338), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_315), .B(n_400), .Y(n_406) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g362 ( .A(n_318), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g428 ( .A(n_318), .Y(n_428) );
OAI222xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_324), .B1(n_325), .B2(n_331), .C1(n_332), .C2(n_334), .Y(n_321) );
INVxp67_ASAP7_75t_L g418 ( .A(n_322), .Y(n_418) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_326), .B(n_411), .Y(n_458) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g374 ( .A(n_327), .B(n_371), .Y(n_374) );
INVx3_ASAP7_75t_L g414 ( .A(n_329), .Y(n_414) );
BUFx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g352 ( .A(n_337), .B(n_353), .Y(n_352) );
OAI221xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_343), .B1(n_346), .B2(n_351), .C(n_354), .Y(n_338) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g396 ( .A1(n_340), .A2(n_397), .B(n_399), .Y(n_396) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g350 ( .A(n_344), .Y(n_350) );
OR2x2_ASAP7_75t_L g454 ( .A(n_345), .B(n_390), .Y(n_454) );
NOR2xp67_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_348), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
OAI21xp5_ASAP7_75t_L g448 ( .A1(n_351), .A2(n_380), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OAI21xp5_ASAP7_75t_L g430 ( .A1(n_352), .A2(n_424), .B(n_431), .Y(n_430) );
INVx4_ASAP7_75t_L g361 ( .A(n_353), .Y(n_361) );
OAI31xp33_ASAP7_75t_SL g354 ( .A1(n_355), .A2(n_356), .A3(n_360), .B(n_362), .Y(n_354) );
INVx1_ASAP7_75t_L g412 ( .A(n_356), .Y(n_412) );
NOR2x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g386 ( .A(n_361), .Y(n_386) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_377), .Y(n_364) );
NAND4xp25_ASAP7_75t_L g465 ( .A(n_365), .B(n_377), .C(n_396), .D(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_375), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_370), .B1(n_373), .B2(n_374), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g437 ( .A(n_369), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_370), .B(n_390), .Y(n_398) );
INVx1_ASAP7_75t_SL g411 ( .A(n_373), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_388), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_382), .B2(n_385), .Y(n_378) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVxp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2x1_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_387), .A2(n_450), .B1(n_452), .B2(n_453), .Y(n_449) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NOR3xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_401), .C(n_407), .Y(n_394) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g466 ( .A(n_401), .Y(n_466) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI21xp33_ASAP7_75t_L g467 ( .A1(n_407), .A2(n_468), .B(n_469), .Y(n_467) );
INVxp33_ASAP7_75t_L g468 ( .A(n_408), .Y(n_468) );
AND2x2_ASAP7_75t_L g794 ( .A(n_408), .B(n_434), .Y(n_794) );
NOR2xp67_ASAP7_75t_L g408 ( .A(n_409), .B(n_416), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B1(n_413), .B2(n_415), .Y(n_409) );
OAI21xp5_ASAP7_75t_L g435 ( .A1(n_413), .A2(n_436), .B(n_439), .Y(n_435) );
INVx2_ASAP7_75t_L g423 ( .A(n_414), .Y(n_423) );
NAND3xp33_ASAP7_75t_SL g416 ( .A(n_417), .B(n_421), .C(n_430), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_424), .B1(n_427), .B2(n_429), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVxp33_ASAP7_75t_SL g469 ( .A(n_434), .Y(n_469) );
NOR3x1_ASAP7_75t_L g434 ( .A(n_435), .B(n_448), .C(n_455), .Y(n_434) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_444), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_456), .B(n_459), .Y(n_455) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g796 ( .A(n_465), .Y(n_796) );
CKINVDCx11_ASAP7_75t_R g470 ( .A(n_471), .Y(n_470) );
AND2x6_ASAP7_75t_SL g471 ( .A(n_472), .B(n_473), .Y(n_471) );
OR2x6_ASAP7_75t_SL g767 ( .A(n_472), .B(n_768), .Y(n_767) );
OR2x2_ASAP7_75t_L g776 ( .A(n_472), .B(n_473), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_472), .B(n_768), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g768 ( .A(n_473), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_479), .B(n_642), .Y(n_478) );
NOR4xp25_ASAP7_75t_L g479 ( .A(n_480), .B(n_585), .C(n_624), .D(n_631), .Y(n_479) );
OAI221xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_506), .B1(n_543), .B2(n_552), .C(n_571), .Y(n_480) );
OR2x2_ASAP7_75t_L g715 ( .A(n_481), .B(n_577), .Y(n_715) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g630 ( .A(n_482), .B(n_555), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_482), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_SL g695 ( .A(n_482), .B(n_696), .Y(n_695) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_495), .Y(n_482) );
AND2x4_ASAP7_75t_SL g554 ( .A(n_483), .B(n_555), .Y(n_554) );
INVx3_ASAP7_75t_L g576 ( .A(n_483), .Y(n_576) );
AND2x2_ASAP7_75t_L g611 ( .A(n_483), .B(n_584), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_483), .B(n_496), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_483), .B(n_578), .Y(n_663) );
OR2x2_ASAP7_75t_L g741 ( .A(n_483), .B(n_555), .Y(n_741) );
AND2x4_ASAP7_75t_L g483 ( .A(n_484), .B(n_489), .Y(n_483) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g563 ( .A(n_496), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_496), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g589 ( .A(n_496), .Y(n_589) );
OR2x2_ASAP7_75t_L g594 ( .A(n_496), .B(n_578), .Y(n_594) );
AND2x2_ASAP7_75t_L g607 ( .A(n_496), .B(n_565), .Y(n_607) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_496), .Y(n_610) );
INVx1_ASAP7_75t_L g622 ( .A(n_496), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_496), .B(n_576), .Y(n_687) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_503), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_507), .B(n_516), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g551 ( .A(n_508), .B(n_535), .Y(n_551) );
AND2x4_ASAP7_75t_L g581 ( .A(n_508), .B(n_520), .Y(n_581) );
INVx2_ASAP7_75t_L g615 ( .A(n_508), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_508), .B(n_535), .Y(n_673) );
AND2x2_ASAP7_75t_L g720 ( .A(n_508), .B(n_549), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_514), .Y(n_509) );
AOI222xp33_ASAP7_75t_L g708 ( .A1(n_516), .A2(n_580), .B1(n_623), .B2(n_683), .C1(n_709), .C2(n_711), .Y(n_708) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_528), .Y(n_517) );
AND2x2_ASAP7_75t_L g627 ( .A(n_518), .B(n_547), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_518), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g756 ( .A(n_518), .B(n_596), .Y(n_756) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_519), .A2(n_587), .B(n_591), .Y(n_586) );
AND2x2_ASAP7_75t_L g667 ( .A(n_519), .B(n_550), .Y(n_667) );
OR2x2_ASAP7_75t_L g692 ( .A(n_519), .B(n_551), .Y(n_692) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx5_ASAP7_75t_L g546 ( .A(n_520), .Y(n_546) );
AND2x2_ASAP7_75t_L g633 ( .A(n_520), .B(n_615), .Y(n_633) );
AND2x2_ASAP7_75t_L g659 ( .A(n_520), .B(n_535), .Y(n_659) );
OR2x2_ASAP7_75t_L g662 ( .A(n_520), .B(n_549), .Y(n_662) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_520), .Y(n_680) );
AND2x4_ASAP7_75t_SL g737 ( .A(n_520), .B(n_614), .Y(n_737) );
OR2x2_ASAP7_75t_L g746 ( .A(n_520), .B(n_573), .Y(n_746) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g579 ( .A(n_528), .Y(n_579) );
AOI221xp5_ASAP7_75t_SL g697 ( .A1(n_528), .A2(n_581), .B1(n_698), .B2(n_700), .C(n_701), .Y(n_697) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_535), .Y(n_528) );
OR2x2_ASAP7_75t_L g636 ( .A(n_529), .B(n_606), .Y(n_636) );
OR2x2_ASAP7_75t_L g646 ( .A(n_529), .B(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g672 ( .A(n_529), .B(n_673), .Y(n_672) );
AND2x4_ASAP7_75t_L g678 ( .A(n_529), .B(n_597), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_529), .B(n_661), .Y(n_690) );
INVx2_ASAP7_75t_L g703 ( .A(n_529), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_529), .B(n_581), .Y(n_724) );
AND2x2_ASAP7_75t_L g728 ( .A(n_529), .B(n_550), .Y(n_728) );
AND2x2_ASAP7_75t_L g736 ( .A(n_529), .B(n_737), .Y(n_736) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g549 ( .A(n_530), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_535), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g580 ( .A(n_535), .B(n_549), .Y(n_580) );
INVx2_ASAP7_75t_L g597 ( .A(n_535), .Y(n_597) );
AND2x4_ASAP7_75t_L g614 ( .A(n_535), .B(n_615), .Y(n_614) );
HB1xp67_ASAP7_75t_L g719 ( .A(n_535), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_541), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_547), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g726 ( .A(n_545), .B(n_548), .Y(n_726) );
AND2x4_ASAP7_75t_L g572 ( .A(n_546), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g613 ( .A(n_546), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g640 ( .A(n_546), .B(n_580), .Y(n_640) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
AND2x2_ASAP7_75t_L g744 ( .A(n_548), .B(n_745), .Y(n_744) );
BUFx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g596 ( .A(n_549), .B(n_597), .Y(n_596) );
OAI21xp5_ASAP7_75t_SL g616 ( .A1(n_550), .A2(n_617), .B(n_623), .Y(n_616) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_563), .Y(n_553) );
INVx1_ASAP7_75t_SL g670 ( .A(n_554), .Y(n_670) );
AND2x2_ASAP7_75t_L g700 ( .A(n_554), .B(n_610), .Y(n_700) );
AND2x4_ASAP7_75t_L g711 ( .A(n_554), .B(n_712), .Y(n_711) );
OR2x2_ASAP7_75t_L g577 ( .A(n_555), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g584 ( .A(n_555), .Y(n_584) );
AND2x4_ASAP7_75t_L g590 ( .A(n_555), .B(n_576), .Y(n_590) );
INVx2_ASAP7_75t_L g601 ( .A(n_555), .Y(n_601) );
INVx1_ASAP7_75t_L g650 ( .A(n_555), .Y(n_650) );
OR2x2_ASAP7_75t_L g671 ( .A(n_555), .B(n_655), .Y(n_671) );
OR2x2_ASAP7_75t_L g685 ( .A(n_555), .B(n_565), .Y(n_685) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_555), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_555), .B(n_607), .Y(n_757) );
OR2x6_ASAP7_75t_L g555 ( .A(n_556), .B(n_562), .Y(n_555) );
INVx1_ASAP7_75t_L g602 ( .A(n_563), .Y(n_602) );
AND2x2_ASAP7_75t_L g735 ( .A(n_563), .B(n_601), .Y(n_735) );
AND2x2_ASAP7_75t_L g760 ( .A(n_563), .B(n_590), .Y(n_760) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g578 ( .A(n_565), .Y(n_578) );
BUFx3_ASAP7_75t_L g620 ( .A(n_565), .Y(n_620) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_565), .Y(n_647) );
INVx1_ASAP7_75t_L g656 ( .A(n_565), .Y(n_656) );
AOI33xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_574), .A3(n_579), .B1(n_580), .B2(n_581), .B3(n_582), .Y(n_571) );
AOI21x1_ASAP7_75t_SL g674 ( .A1(n_572), .A2(n_596), .B(n_658), .Y(n_674) );
INVx2_ASAP7_75t_L g704 ( .A(n_572), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_572), .B(n_703), .Y(n_710) );
AND2x2_ASAP7_75t_L g658 ( .A(n_573), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g621 ( .A(n_576), .B(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g722 ( .A(n_577), .Y(n_722) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_578), .Y(n_712) );
OAI32xp33_ASAP7_75t_L g761 ( .A1(n_579), .A2(n_581), .A3(n_757), .B1(n_762), .B2(n_764), .Y(n_761) );
AND2x2_ASAP7_75t_L g679 ( .A(n_580), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_SL g669 ( .A(n_581), .Y(n_669) );
AND2x2_ASAP7_75t_L g734 ( .A(n_581), .B(n_678), .Y(n_734) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OAI221xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_595), .B1(n_598), .B2(n_612), .C(n_616), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_589), .B(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_590), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_590), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_590), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g639 ( .A(n_594), .Y(n_639) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NOR3xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_603), .C(n_608), .Y(n_598) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_600), .A2(n_662), .B1(n_702), .B2(n_705), .Y(n_701) );
OR2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g605 ( .A(n_601), .Y(n_605) );
NOR2x1p5_ASAP7_75t_L g619 ( .A(n_601), .B(n_620), .Y(n_619) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_601), .Y(n_641) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI322xp33_ASAP7_75t_L g668 ( .A1(n_604), .A2(n_646), .A3(n_669), .B1(n_670), .B2(n_671), .C1(n_672), .C2(n_674), .Y(n_668) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g624 ( .A1(n_606), .A2(n_625), .B(n_626), .C(n_628), .Y(n_624) );
OR2x2_ASAP7_75t_L g716 ( .A(n_606), .B(n_670), .Y(n_716) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g623 ( .A(n_607), .B(n_611), .Y(n_623) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g629 ( .A(n_613), .B(n_630), .Y(n_629) );
INVx3_ASAP7_75t_SL g661 ( .A(n_614), .Y(n_661) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_618), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVx1_ASAP7_75t_SL g665 ( .A(n_621), .Y(n_665) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_622), .Y(n_707) );
OR2x6_ASAP7_75t_SL g762 ( .A(n_625), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVxp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI211xp5_ASAP7_75t_L g752 ( .A1(n_630), .A2(n_753), .B(n_754), .C(n_761), .Y(n_752) );
O2A1O1Ixp33_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_634), .B(n_637), .C(n_641), .Y(n_631) );
OAI211xp5_ASAP7_75t_SL g643 ( .A1(n_632), .A2(n_644), .B(n_651), .C(n_675), .Y(n_643) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVxp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
NOR3xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_688), .C(n_732), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_648), .Y(n_644) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_647), .Y(n_739) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g694 ( .A(n_650), .Y(n_694) );
NOR3xp33_ASAP7_75t_SL g651 ( .A(n_652), .B(n_664), .C(n_668), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_657), .B1(n_660), .B2(n_663), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g696 ( .A(n_656), .Y(n_696) );
INVxp67_ASAP7_75t_SL g763 ( .A(n_656), .Y(n_763) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_SL g749 ( .A(n_662), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
OR2x2_ASAP7_75t_L g699 ( .A(n_665), .B(n_685), .Y(n_699) );
OR2x2_ASAP7_75t_L g750 ( .A(n_665), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g748 ( .A(n_673), .Y(n_748) );
OR2x2_ASAP7_75t_L g764 ( .A(n_673), .B(n_703), .Y(n_764) );
OAI21xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_679), .B(n_681), .Y(n_675) );
OAI31xp33_ASAP7_75t_L g689 ( .A1(n_676), .A2(n_690), .A3(n_691), .B(n_693), .Y(n_689) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
INVx1_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
AND2x4_ASAP7_75t_L g721 ( .A(n_686), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND4xp25_ASAP7_75t_SL g688 ( .A(n_689), .B(n_697), .C(n_708), .D(n_713), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_696), .Y(n_731) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
INVxp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_717), .B1(n_721), .B2(n_723), .C(n_725), .Y(n_713) );
NAND2xp33_ASAP7_75t_SL g714 ( .A(n_715), .B(n_716), .Y(n_714) );
INVx1_ASAP7_75t_L g758 ( .A(n_717), .Y(n_758) );
AND2x2_ASAP7_75t_SL g717 ( .A(n_718), .B(n_720), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AOI21xp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B(n_729), .Y(n_725) );
INVx1_ASAP7_75t_L g753 ( .A(n_727), .Y(n_753) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g732 ( .A(n_733), .B(n_752), .Y(n_732) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B1(n_736), .B2(n_738), .C(n_742), .Y(n_733) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
AOI21xp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_747), .B(n_750), .Y(n_742) );
INVxp33_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_757), .B1(n_758), .B2(n_759), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
CKINVDCx5p33_ASAP7_75t_R g765 ( .A(n_766), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_766), .Y(n_772) );
CKINVDCx11_ASAP7_75t_R g766 ( .A(n_767), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g773 ( .A(n_774), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g774 ( .A(n_775), .Y(n_774) );
INVx3_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_786), .Y(n_779) );
INVxp67_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND2xp5_ASAP7_75t_SL g781 ( .A(n_782), .B(n_785), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
OR2x2_ASAP7_75t_SL g804 ( .A(n_783), .B(n_785), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g806 ( .A1(n_783), .A2(n_807), .B(n_810), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_786), .A2(n_790), .B(n_800), .Y(n_789) );
BUFx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
BUFx2_ASAP7_75t_R g801 ( .A(n_787), .Y(n_801) );
BUFx2_ASAP7_75t_L g811 ( .A(n_787), .Y(n_811) );
INVxp67_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OAI22xp33_ASAP7_75t_SL g790 ( .A1(n_791), .A2(n_792), .B1(n_797), .B2(n_798), .Y(n_790) );
INVxp67_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND3x1_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .C(n_796), .Y(n_793) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NOR2xp33_ASAP7_75t_SL g800 ( .A(n_801), .B(n_802), .Y(n_800) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
CKINVDCx11_ASAP7_75t_R g807 ( .A(n_808), .Y(n_807) );
CKINVDCx8_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
endmodule