module fake_jpeg_13018_n_177 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

OR2x2_ASAP7_75t_SL g55 ( 
.A(n_21),
.B(n_6),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_12),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_27),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_30),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_78),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_62),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_58),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_68),
.B1(n_58),
.B2(n_60),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_83),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_57),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_76),
.Y(n_97)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_86),
.Y(n_91)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_101),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_62),
.B(n_56),
.Y(n_106)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_97),
.Y(n_118)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_70),
.Y(n_117)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_39),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_111),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_75),
.C(n_69),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_113),
.C(n_9),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_108),
.B1(n_15),
.B2(n_16),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_110),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_68),
.B1(n_67),
.B2(n_61),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_74),
.Y(n_110)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_26),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_65),
.C(n_71),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_72),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_121),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_SL g115 ( 
.A1(n_101),
.A2(n_64),
.B(n_65),
.C(n_67),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_4),
.B(n_5),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_10),
.Y(n_138)
);

INVx4_ASAP7_75t_SL g119 ( 
.A(n_92),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_87),
.Y(n_121)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_51),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_123),
.B(n_132),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_116),
.A2(n_63),
.B1(n_52),
.B2(n_64),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_131),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_1),
.B(n_3),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_128),
.B(n_29),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_18),
.B1(n_48),
.B2(n_43),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_134),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_7),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_8),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_8),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_137),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_24),
.C(n_25),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_9),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_141),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_13),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_140),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_14),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_115),
.B(n_17),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_144),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_23),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_155),
.C(n_157),
.Y(n_165)
);

A2O1A1O1Ixp25_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_126),
.B(n_153),
.C(n_146),
.D(n_136),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_32),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_37),
.C(n_41),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_162),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_159),
.B(n_129),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_127),
.B1(n_128),
.B2(n_42),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_169),
.B(n_149),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_168),
.A2(n_164),
.B(n_162),
.C(n_160),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_171),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_152),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_155),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_156),
.Y(n_175)
);

OA21x2_ASAP7_75t_SL g176 ( 
.A1(n_175),
.A2(n_167),
.B(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);


endmodule