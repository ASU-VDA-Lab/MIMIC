module real_jpeg_33474_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_698, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_698;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_578;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_611;
wire n_221;
wire n_489;
wire n_393;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_411;
wire n_382;
wire n_278;
wire n_689;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_642;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_400;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_694;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_468;
wire n_133;
wire n_447;
wire n_257;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_0),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_0),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g274 ( 
.A(n_0),
.Y(n_274)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_0),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_1),
.A2(n_178),
.B1(n_179),
.B2(n_184),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_1),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_1),
.A2(n_178),
.B1(n_237),
.B2(n_242),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_1),
.A2(n_178),
.B1(n_390),
.B2(n_394),
.Y(n_389)
);

OAI22xp33_ASAP7_75t_SL g641 ( 
.A1(n_1),
.A2(n_178),
.B1(n_642),
.B2(n_644),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_3),
.A2(n_126),
.B1(n_129),
.B2(n_130),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_3),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_3),
.A2(n_129),
.B1(n_290),
.B2(n_294),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_3),
.A2(n_129),
.B1(n_401),
.B2(n_403),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_3),
.A2(n_129),
.B1(n_266),
.B2(n_500),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_4),
.A2(n_163),
.B1(n_168),
.B2(n_169),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_4),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_4),
.A2(n_168),
.B1(n_336),
.B2(n_340),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_4),
.A2(n_168),
.B1(n_447),
.B2(n_449),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g637 ( 
.A1(n_4),
.A2(n_168),
.B1(n_200),
.B2(n_638),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_5),
.B(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_5),
.A2(n_55),
.B(n_218),
.Y(n_287)
);

INVx2_ASAP7_75t_R g325 ( 
.A(n_5),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_5),
.A2(n_325),
.B1(n_516),
.B2(n_518),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_5),
.B(n_112),
.Y(n_532)
);

OAI22xp33_ASAP7_75t_SL g587 ( 
.A1(n_5),
.A2(n_188),
.B1(n_588),
.B2(n_592),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_6),
.A2(n_67),
.B1(n_71),
.B2(n_74),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_6),
.A2(n_74),
.B1(n_351),
.B2(n_354),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_6),
.A2(n_74),
.B1(n_438),
.B2(n_442),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g627 ( 
.A1(n_6),
.A2(n_74),
.B1(n_628),
.B2(n_631),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_8),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_8),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_9),
.Y(n_167)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_9),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_9),
.Y(n_192)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_9),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_10),
.A2(n_55),
.B1(n_60),
.B2(n_64),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_10),
.A2(n_64),
.B1(n_265),
.B2(n_270),
.Y(n_264)
);

AOI22x1_ASAP7_75t_L g415 ( 
.A1(n_10),
.A2(n_64),
.B1(n_416),
.B2(n_418),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_10),
.A2(n_64),
.B1(n_366),
.B2(n_623),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_11),
.A2(n_135),
.B1(n_141),
.B2(n_145),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_11),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_11),
.A2(n_145),
.B1(n_373),
.B2(n_375),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_11),
.A2(n_145),
.B1(n_479),
.B2(n_484),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_11),
.A2(n_145),
.B1(n_529),
.B2(n_531),
.Y(n_528)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_12),
.Y(n_229)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_12),
.Y(n_235)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_13),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_14),
.A2(n_257),
.B1(n_260),
.B2(n_261),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_14),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_14),
.A2(n_260),
.B1(n_318),
.B2(n_322),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_14),
.A2(n_260),
.B1(n_365),
.B2(n_368),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_14),
.A2(n_61),
.B1(n_94),
.B2(n_260),
.Y(n_456)
);

AOI22x1_ASAP7_75t_SL g92 ( 
.A1(n_15),
.A2(n_93),
.B1(n_97),
.B2(n_100),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_15),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_15),
.A2(n_100),
.B1(n_278),
.B2(n_283),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_15),
.A2(n_100),
.B1(n_242),
.B2(n_510),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_SL g579 ( 
.A1(n_15),
.A2(n_100),
.B1(n_580),
.B2(n_582),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_16),
.B(n_689),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_16),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_17),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_17),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_17),
.A2(n_106),
.B1(n_307),
.B2(n_313),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_17),
.A2(n_106),
.B1(n_257),
.B2(n_537),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_17),
.A2(n_106),
.B1(n_589),
.B2(n_591),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_18),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_18),
.Y(n_124)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_18),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_18),
.Y(n_512)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_19),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_19),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_19),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_691),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_81),
.B(n_688),
.Y(n_21)
);

INVxp33_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_76),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_24),
.B(n_680),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_24),
.B(n_680),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_25),
.B(n_77),
.Y(n_690)
);

NAND4xp25_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_53),
.C(n_65),
.D(n_75),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_49),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_L g65 ( 
.A(n_27),
.B(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_27),
.A2(n_49),
.B1(n_637),
.B2(n_640),
.Y(n_636)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_28),
.A2(n_50),
.B1(n_456),
.B2(n_641),
.Y(n_653)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_29),
.A2(n_51),
.B1(n_103),
.B2(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_29),
.A2(n_51),
.B1(n_92),
.B2(n_372),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_29),
.A2(n_51),
.B1(n_372),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_41),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_34),
.Y(n_203)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_34),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_36),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_36),
.Y(n_212)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_37),
.Y(n_402)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_37),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_37),
.Y(n_645)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_41)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_42),
.Y(n_393)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_43),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_43),
.Y(n_634)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_46),
.Y(n_151)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_46),
.Y(n_626)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_66),
.B(n_78),
.Y(n_77)
);

OAI21x1_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_90),
.B(n_101),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g649 ( 
.A1(n_49),
.A2(n_54),
.B1(n_78),
.B2(n_637),
.Y(n_649)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22x1_ASAP7_75t_L g455 ( 
.A1(n_50),
.A2(n_79),
.B1(n_400),
.B2(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2x1_ASAP7_75t_R g324 ( 
.A(n_51),
.B(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_56),
.Y(n_219)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_58),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_59),
.Y(n_374)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_63),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_616),
.B(n_681),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_468),
.B(n_611),
.Y(n_83)
);

NAND4xp25_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_328),
.C(n_425),
.D(n_460),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_298),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_86),
.B(n_298),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_220),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_87),
.A2(n_462),
.B(n_463),
.Y(n_461)
);

XNOR2x1_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_158),
.Y(n_87)
);

XNOR2x1_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_110),
.Y(n_88)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_89),
.Y(n_331)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_110),
.B(n_158),
.C(n_331),
.Y(n_330)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_125),
.B1(n_134),
.B2(n_146),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_111),
.A2(n_134),
.B1(n_146),
.B2(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_111),
.A2(n_277),
.B(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_111),
.A2(n_125),
.B1(n_146),
.B2(n_364),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_111),
.A2(n_146),
.B1(n_306),
.B2(n_515),
.Y(n_514)
);

OAI22xp33_ASAP7_75t_SL g621 ( 
.A1(n_111),
.A2(n_146),
.B1(n_622),
.B2(n_627),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_SL g654 ( 
.A1(n_111),
.A2(n_146),
.B1(n_622),
.B2(n_655),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22x1_ASAP7_75t_SL g387 ( 
.A1(n_112),
.A2(n_304),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_112),
.A2(n_304),
.B1(n_389),
.B2(n_446),
.Y(n_445)
);

OAI21xp33_ASAP7_75t_SL g647 ( 
.A1(n_112),
.A2(n_304),
.B(n_648),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AO21x2_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_147),
.B(n_152),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_117),
.B1(n_120),
.B2(n_123),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_118),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_118),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_119),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_119),
.Y(n_342)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_119),
.Y(n_441)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_123),
.B(n_253),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_123),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_123),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_124),
.Y(n_241)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_124),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_124),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_124),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_128),
.Y(n_450)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_133),
.Y(n_285)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_133),
.Y(n_630)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_140),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_140),
.Y(n_282)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_143),
.Y(n_448)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_144),
.Y(n_519)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_146),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_152),
.A2(n_489),
.B(n_494),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_154),
.Y(n_313)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_194),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_159),
.A2(n_160),
.B1(n_194),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_171),
.B1(n_177),
.B2(n_187),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_162),
.A2(n_188),
.B1(n_264),
.B2(n_272),
.Y(n_263)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_167),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_167),
.Y(n_530)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_170),
.Y(n_271)
);

BUFx2_ASAP7_75t_SL g323 ( 
.A(n_170),
.Y(n_323)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_172),
.B(n_325),
.Y(n_594)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_176),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_176),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_177),
.A2(n_187),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_183),
.Y(n_561)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx2_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

AO22x1_ASAP7_75t_L g498 ( 
.A1(n_187),
.A2(n_317),
.B1(n_499),
.B2(n_503),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_187),
.A2(n_345),
.B1(n_577),
.B2(n_578),
.Y(n_576)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_188),
.A2(n_264),
.B(n_344),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_188),
.A2(n_350),
.B(n_411),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_188),
.A2(n_524),
.B1(n_527),
.B2(n_528),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_188),
.A2(n_524),
.B1(n_579),
.B2(n_588),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_191),
.Y(n_583)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_192),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_193),
.Y(n_503)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_193),
.Y(n_592)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_194),
.Y(n_327)
);

OAI22x1_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_204),
.B1(n_207),
.B2(n_217),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx11_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_216),
.Y(n_396)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_275),
.B1(n_296),
.B2(n_297),
.Y(n_220)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_221),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_263),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_222),
.B(n_263),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_236),
.B1(n_245),
.B2(n_256),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_223),
.A2(n_236),
.B1(n_245),
.B2(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_223),
.A2(n_245),
.B1(n_509),
.B2(n_535),
.Y(n_534)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_225),
.Y(n_295)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AO21x2_ASAP7_75t_L g245 ( 
.A1(n_226),
.A2(n_246),
.B(n_252),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_229),
.Y(n_563)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_245),
.A2(n_256),
.B1(n_289),
.B2(n_295),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_245),
.A2(n_295),
.B1(n_335),
.B2(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_245),
.Y(n_435)
);

AO21x1_ASAP7_75t_L g635 ( 
.A1(n_245),
.A2(n_295),
.B(n_437),
.Y(n_635)
);

AOI21xp33_ASAP7_75t_SL g652 ( 
.A1(n_245),
.A2(n_295),
.B(n_437),
.Y(n_652)
);

NAND2xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_250),
.Y(n_485)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_250),
.Y(n_554)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_251),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_251),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_252),
.Y(n_567)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_259),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_269),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_269),
.Y(n_356)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_269),
.Y(n_502)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_269),
.Y(n_597)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_270),
.Y(n_531)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_272),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_275),
.Y(n_297)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_286),
.C(n_288),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_288),
.Y(n_300)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_282),
.Y(n_517)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_300),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_289),
.A2(n_295),
.B1(n_477),
.B2(n_486),
.Y(n_476)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_295),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g600 ( 
.A(n_295),
.B(n_325),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_R g462 ( 
.A(n_296),
.B(n_297),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_R g463 ( 
.A(n_296),
.B(n_297),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.C(n_326),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g607 ( 
.A(n_299),
.B(n_608),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_301),
.B(n_326),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_314),
.C(n_324),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_302),
.B(n_473),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_309),
.Y(n_497)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_311),
.Y(n_369)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_312),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_314),
.A2(n_315),
.B1(n_324),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_324),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_325),
.B(n_490),
.Y(n_489)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_325),
.B(n_495),
.C(n_497),
.Y(n_494)
);

OAI21xp33_ASAP7_75t_SL g548 ( 
.A1(n_325),
.A2(n_549),
.B(n_551),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_325),
.B(n_552),
.Y(n_551)
);

A2O1A1O1Ixp25_ASAP7_75t_L g611 ( 
.A1(n_328),
.A2(n_425),
.B(n_612),
.C(n_614),
.D(n_615),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_381),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_329),
.B(n_381),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_332),
.C(n_357),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_330),
.B(n_465),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_333),
.A2(n_358),
.B1(n_359),
.B2(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_333),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_343),
.Y(n_333)
);

NAND2xp33_ASAP7_75t_SL g384 ( 
.A(n_334),
.B(n_343),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_349),
.Y(n_344)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_352),
.Y(n_566)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_356),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_359),
.B1(n_360),
.B2(n_380),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_358),
.B(n_362),
.C(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_360),
.B(n_466),
.Y(n_465)
);

AO21x1_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_370),
.B(n_379),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_370),
.Y(n_379)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_364),
.Y(n_388)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_370),
.Y(n_424)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_374),
.Y(n_373)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_407),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_383),
.B(n_408),
.C(n_427),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_384),
.A2(n_385),
.B1(n_405),
.B2(n_406),
.Y(n_383)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_384),
.Y(n_406)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_385),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_386),
.A2(n_387),
.B1(n_397),
.B2(n_398),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_386),
.B(n_406),
.C(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_398),
.Y(n_430)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_423),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_413),
.B(n_422),
.Y(n_408)
);

NAND2xp33_ASAP7_75t_SL g422 ( 
.A(n_409),
.B(n_414),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_409),
.A2(n_410),
.B1(n_454),
.B2(n_455),
.Y(n_453)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_410),
.B(n_414),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_410),
.Y(n_667)
);

INVx8_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_415),
.Y(n_434)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx2_ASAP7_75t_SL g418 ( 
.A(n_419),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx5_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_423),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_428),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_426),
.B(n_428),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_431),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g671 ( 
.A(n_429),
.B(n_459),
.C(n_672),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_452),
.B1(n_458),
.B2(n_459),
.Y(n_431)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_432),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_445),
.B(n_451),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_445),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_435),
.B1(n_436),
.B2(n_444),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_435),
.Y(n_486)
);

AOI22x1_ASAP7_75t_L g507 ( 
.A1(n_435),
.A2(n_444),
.B1(n_478),
.B2(n_508),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_435),
.A2(n_444),
.B1(n_536),
.B2(n_548),
.Y(n_547)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_440),
.Y(n_550)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_441),
.Y(n_538)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_446),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx8_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_451),
.Y(n_663)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_452),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_452),
.Y(n_672)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_457),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_455),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_457),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_464),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_461),
.B(n_464),
.C(n_613),
.Y(n_612)
);

AOI21x1_ASAP7_75t_SL g468 ( 
.A1(n_469),
.A2(n_606),
.B(n_610),
.Y(n_468)
);

OAI21x1_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_520),
.B(n_605),
.Y(n_469)
);

NOR2x1_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_504),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_471),
.B(n_504),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_475),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_472),
.B(n_476),
.C(n_487),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_487),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_498),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_488),
.B(n_498),
.Y(n_505)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_493),
.Y(n_496)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_499),
.Y(n_527)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_501),
.Y(n_591)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_502),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_506),
.C(n_513),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_505),
.B(n_540),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

OA21x2_ASAP7_75t_L g540 ( 
.A1(n_507),
.A2(n_513),
.B(n_541),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_507),
.B(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_514),
.Y(n_542)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

AOI31xp67_ASAP7_75t_L g520 ( 
.A1(n_521),
.A2(n_543),
.A3(n_571),
.B(n_604),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_539),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_522),
.B(n_539),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_532),
.C(n_533),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_523),
.B(n_569),
.Y(n_568)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVxp33_ASAP7_75t_L g577 ( 
.A(n_528),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_530),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_532),
.B(n_534),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_570),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_568),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_545),
.B(n_568),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_546),
.B(n_555),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_546),
.B(n_556),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_546),
.A2(n_556),
.B(n_575),
.Y(n_603)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_547),
.B(n_555),
.Y(n_575)
);

INVxp67_ASAP7_75t_SL g549 ( 
.A(n_550),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_551),
.Y(n_564)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_557),
.A2(n_564),
.B1(n_565),
.B2(n_567),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_SL g557 ( 
.A(n_558),
.B(n_562),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

NAND3xp33_ASAP7_75t_L g571 ( 
.A(n_570),
.B(n_572),
.C(n_584),
.Y(n_571)
);

AO21x1_ASAP7_75t_L g572 ( 
.A1(n_573),
.A2(n_574),
.B(n_576),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_576),
.B(n_603),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_585),
.B(n_602),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_586),
.A2(n_598),
.B(n_601),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_587),
.B(n_593),
.Y(n_586)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_594),
.B(n_595),
.Y(n_593)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

BUFx12f_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_599),
.B(n_600),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_599),
.B(n_600),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_607),
.B(n_609),
.Y(n_606)
);

NOR2x1_ASAP7_75t_L g610 ( 
.A(n_607),
.B(n_609),
.Y(n_610)
);

NAND3xp33_ASAP7_75t_L g616 ( 
.A(n_617),
.B(n_659),
.C(n_679),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_SL g682 ( 
.A1(n_618),
.A2(n_683),
.B(n_686),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_619),
.B(n_650),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_619),
.B(n_650),
.Y(n_686)
);

XNOR2xp5_ASAP7_75t_SL g619 ( 
.A(n_620),
.B(n_646),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g680 ( 
.A(n_620),
.B(n_647),
.C(n_649),
.Y(n_680)
);

MAJx2_ASAP7_75t_L g620 ( 
.A(n_621),
.B(n_635),
.C(n_636),
.Y(n_620)
);

OA22x2_ASAP7_75t_L g657 ( 
.A1(n_621),
.A2(n_635),
.B1(n_652),
.B2(n_658),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_621),
.Y(n_658)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_624),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_626),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_627),
.Y(n_648)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_629),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_632),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_633),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_634),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_SL g669 ( 
.A1(n_635),
.A2(n_652),
.B1(n_654),
.B2(n_670),
.Y(n_669)
);

XNOR2xp5_ASAP7_75t_L g656 ( 
.A(n_636),
.B(n_657),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g678 ( 
.A(n_636),
.B(n_653),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_641),
.Y(n_640)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_643),
.Y(n_642)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_647),
.B(n_649),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_651),
.B(n_653),
.C(n_656),
.Y(n_650)
);

XNOR2xp5_ASAP7_75t_L g676 ( 
.A(n_651),
.B(n_677),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_652),
.B(n_653),
.C(n_654),
.Y(n_651)
);

XNOR2xp5_ASAP7_75t_L g668 ( 
.A(n_653),
.B(n_669),
.Y(n_668)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_654),
.Y(n_670)
);

XNOR2xp5_ASAP7_75t_L g677 ( 
.A(n_657),
.B(n_678),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_SL g659 ( 
.A(n_660),
.B(n_673),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_661),
.B(n_671),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_661),
.B(n_671),
.Y(n_684)
);

XOR2xp5_ASAP7_75t_L g661 ( 
.A(n_662),
.B(n_668),
.Y(n_661)
);

XOR2xp5_ASAP7_75t_L g662 ( 
.A(n_663),
.B(n_664),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_663),
.B(n_664),
.C(n_668),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_SL g664 ( 
.A1(n_665),
.A2(n_666),
.B1(n_667),
.B2(n_698),
.Y(n_664)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_674),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_SL g683 ( 
.A1(n_674),
.A2(n_684),
.B(n_685),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_675),
.B(n_676),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_675),
.B(n_676),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_679),
.A2(n_682),
.B(n_687),
.Y(n_681)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_690),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_692),
.B(n_696),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_693),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_694),
.Y(n_693)
);

BUFx12f_ASAP7_75t_SL g694 ( 
.A(n_695),
.Y(n_694)
);


endmodule