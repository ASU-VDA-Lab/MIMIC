module fake_jpeg_26014_n_199 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_199);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_28),
.B1(n_26),
.B2(n_24),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_53),
.B1(n_31),
.B2(n_37),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_40),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_28),
.B1(n_26),
.B2(n_29),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_54),
.B1(n_19),
.B2(n_18),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_25),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_25),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_28),
.B1(n_26),
.B2(n_17),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_21),
.B1(n_29),
.B2(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_57),
.Y(n_84)
);

BUFx2_ASAP7_75t_SL g56 ( 
.A(n_42),
.Y(n_56)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_63),
.Y(n_79)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_31),
.B1(n_47),
.B2(n_41),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_73),
.B1(n_74),
.B2(n_70),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_30),
.B1(n_22),
.B2(n_20),
.Y(n_100)
);

OR2x4_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_38),
.Y(n_66)
);

AO21x1_ASAP7_75t_L g99 ( 
.A1(n_66),
.A2(n_36),
.B(n_33),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_72),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_27),
.C(n_30),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_32),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_21),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_38),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_43),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_27),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_66),
.A2(n_38),
.B(n_34),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_99),
.B(n_33),
.Y(n_116)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_68),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_34),
.B1(n_40),
.B2(n_36),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_94),
.B1(n_74),
.B2(n_73),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_40),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_57),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_98),
.C(n_61),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_55),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_61),
.B(n_36),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_76),
.B1(n_77),
.B2(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_109),
.C(n_112),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_105),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_95),
.B(n_69),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

XNOR2x2_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_72),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_116),
.B(n_84),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_79),
.A2(n_67),
.B1(n_33),
.B2(n_20),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_58),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_79),
.A2(n_20),
.B1(n_22),
.B2(n_4),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_98),
.B1(n_90),
.B2(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_86),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_91),
.C(n_109),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_128),
.C(n_98),
.Y(n_149)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_138),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_80),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_137),
.B(n_80),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_132),
.B(n_139),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_133),
.A2(n_120),
.B(n_112),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_104),
.A2(n_84),
.B(n_88),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_87),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_136),
.Y(n_162)
);

AOI221xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_105),
.B1(n_113),
.B2(n_116),
.C(n_120),
.Y(n_143)
);

AOI321xp33_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_144),
.A3(n_156),
.B1(n_123),
.B2(n_126),
.C(n_136),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_107),
.B1(n_117),
.B2(n_110),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_146),
.B1(n_153),
.B2(n_142),
.Y(n_163)
);

OAI22x1_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_99),
.B1(n_86),
.B2(n_122),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_151),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_152),
.C(n_154),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_155),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_93),
.C(n_97),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_99),
.C(n_85),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

OAI322xp33_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_22),
.A3(n_20),
.B1(n_14),
.B2(n_13),
.C1(n_85),
.C2(n_7),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_166),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_152),
.B(n_128),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_162),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_165),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_127),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_141),
.C(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_144),
.B(n_14),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_149),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_170),
.C(n_171),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_154),
.C(n_146),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_141),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_176),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_111),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_158),
.C(n_167),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_181),
.C(n_177),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_129),
.C(n_161),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_180),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_173),
.A2(n_96),
.B1(n_20),
.B2(n_4),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_175),
.B(n_168),
.Y(n_187)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_174),
.Y(n_182)
);

AOI31xp67_ASAP7_75t_SL g188 ( 
.A1(n_182),
.A2(n_96),
.A3(n_4),
.B(n_5),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_1),
.B(n_3),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_183),
.A2(n_1),
.B(n_3),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_188),
.C(n_1),
.Y(n_191)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_187),
.Y(n_192)
);

A2O1A1O1Ixp25_ASAP7_75t_L g189 ( 
.A1(n_185),
.A2(n_10),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_189),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_8),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_9),
.C(n_6),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_8),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_195),
.A2(n_192),
.B1(n_8),
.B2(n_9),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_197),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_193),
.Y(n_199)
);


endmodule