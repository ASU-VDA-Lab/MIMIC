module fake_jpeg_29667_n_316 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_21),
.B(n_6),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_31),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_31),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_33),
.B1(n_28),
.B2(n_17),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_60),
.B1(n_15),
.B2(n_17),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_25),
.B1(n_28),
.B2(n_15),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_50),
.B1(n_57),
.B2(n_43),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_62),
.A2(n_81),
.B1(n_88),
.B2(n_93),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_63),
.B(n_83),
.Y(n_104)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_68),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_18),
.B1(n_36),
.B2(n_29),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_40),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_37),
.B1(n_43),
.B2(n_28),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_70),
.A2(n_27),
.B1(n_22),
.B2(n_23),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_24),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_86),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

NAND2x1_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_40),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_73),
.B(n_79),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_46),
.Y(n_95)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

NAND2x1p5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_37),
.B1(n_18),
.B2(n_27),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_85),
.B1(n_54),
.B2(n_68),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_29),
.B1(n_34),
.B2(n_20),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_48),
.A2(n_15),
.B1(n_17),
.B2(n_22),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_55),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_30),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_94),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_44),
.B1(n_45),
.B2(n_22),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_105),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_60),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_120),
.C(n_73),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_23),
.B(n_20),
.C(n_30),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_60),
.Y(n_105)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_111),
.B1(n_73),
.B2(n_83),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_55),
.B1(n_44),
.B2(n_54),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_31),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_31),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_67),
.B(n_76),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_41),
.C(n_27),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_90),
.B1(n_87),
.B2(n_84),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_125),
.B(n_131),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_63),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_126),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_133),
.B1(n_149),
.B2(n_111),
.Y(n_153)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_112),
.B(n_79),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_130),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_97),
.B(n_80),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_119),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_140),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_105),
.A2(n_93),
.B1(n_75),
.B2(n_86),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_134),
.B(n_141),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_113),
.Y(n_162)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_89),
.C(n_64),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_144),
.C(n_147),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_145),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_114),
.B(n_16),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_103),
.B(n_78),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_142),
.B(n_148),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_94),
.C(n_72),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_92),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_31),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_121),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_41),
.C(n_16),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_108),
.B(n_32),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_113),
.A2(n_77),
.B1(n_32),
.B2(n_16),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_153),
.A2(n_16),
.B1(n_7),
.B2(n_8),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_100),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_155),
.B(n_156),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_100),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_109),
.C(n_120),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_158),
.B(n_160),
.C(n_161),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_109),
.C(n_101),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_101),
.C(n_106),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_136),
.B1(n_116),
.B2(n_102),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_177),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_98),
.B1(n_106),
.B2(n_121),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_165),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_200)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_149),
.A2(n_136),
.B1(n_132),
.B2(n_133),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_129),
.B(n_11),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_135),
.A2(n_122),
.B(n_118),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_138),
.B(n_144),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_147),
.A2(n_102),
.B(n_116),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_139),
.B(n_130),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_183),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_189),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_185),
.A2(n_187),
.B(n_195),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_167),
.B1(n_178),
.B2(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_150),
.B1(n_99),
.B2(n_123),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_196),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_200),
.B1(n_202),
.B2(n_171),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_0),
.B(n_1),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_6),
.B1(n_13),
.B2(n_11),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_161),
.A2(n_5),
.B(n_13),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_197),
.B(n_205),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_0),
.B(n_1),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_7),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_152),
.C(n_160),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_151),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_159),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_153),
.A2(n_8),
.B1(n_4),
.B2(n_5),
.Y(n_202)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_158),
.B(n_7),
.CI(n_8),
.CON(n_205),
.SN(n_205)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_154),
.B(n_2),
.Y(n_208)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_168),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_165),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_216),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_188),
.Y(n_216)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_218),
.B(n_222),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_179),
.B1(n_181),
.B2(n_174),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_219),
.A2(n_223),
.B(n_224),
.Y(n_248)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_195),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_198),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_230),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_154),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_226),
.B(n_227),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_189),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_234),
.C(n_152),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_206),
.C(n_207),
.Y(n_233)
);

FAx1_ASAP7_75t_SL g241 ( 
.A(n_233),
.B(n_202),
.CI(n_208),
.CON(n_241),
.SN(n_241)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_173),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_210),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_246),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_236),
.B(n_239),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_210),
.C(n_205),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_184),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_243),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_249),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_183),
.C(n_185),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_247),
.C(n_246),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_199),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_182),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_197),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_251),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_231),
.C(n_209),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_187),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_186),
.C(n_204),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_224),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_215),
.B(n_193),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_228),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_244),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_254),
.Y(n_271)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g256 ( 
.A(n_241),
.Y(n_256)
);

OAI21x1_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_264),
.B(n_258),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_248),
.A2(n_229),
.B(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_217),
.B1(n_215),
.B2(n_225),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_269),
.B1(n_166),
.B2(n_157),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_267),
.Y(n_278)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_227),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_200),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_242),
.A2(n_223),
.B1(n_229),
.B2(n_213),
.Y(n_269)
);

AOI21xp33_ASAP7_75t_L g272 ( 
.A1(n_263),
.A2(n_213),
.B(n_251),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_272),
.A2(n_261),
.B(n_257),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_279),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_268),
.A2(n_253),
.B1(n_240),
.B2(n_192),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_274),
.B(n_275),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_243),
.C(n_222),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_169),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_281),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_166),
.Y(n_282)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_275),
.B(n_270),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_294),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_288),
.Y(n_296)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_293),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_261),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_292),
.Y(n_295)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_157),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_279),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_278),
.C(n_257),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_277),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_298),
.B(n_301),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_287),
.A2(n_282),
.B(n_280),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_299),
.B(n_296),
.Y(n_308)
);

NOR2x1_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_278),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_304),
.B(n_305),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_286),
.C(n_176),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_176),
.Y(n_306)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_9),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_307),
.A2(n_308),
.B(n_299),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_309),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_311),
.A2(n_303),
.B(n_14),
.Y(n_312)
);

MAJx2_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_310),
.C(n_303),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_314),
.A2(n_313),
.B(n_2),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);


endmodule