module fake_jpeg_7877_n_30 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_30);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_30;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_29;
wire n_15;

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_1),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_13),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_10),
.A2(n_6),
.B1(n_3),
.B2(n_12),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_7),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_15),
.B(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_19),
.B(n_6),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_17),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_21),
.B(n_22),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_14),
.A2(n_4),
.B(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_5),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_25),
.C(n_26),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_21),
.C(n_7),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_8),
.B(n_27),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_8),
.Y(n_30)
);


endmodule