module real_jpeg_6250_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_1),
.B(n_147),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_1),
.A2(n_62),
.B1(n_134),
.B2(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_1),
.B(n_248),
.C(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_1),
.B(n_23),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_1),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_1),
.B(n_136),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_2),
.A2(n_125),
.B1(n_126),
.B2(n_130),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_2),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_2),
.A2(n_130),
.B1(n_139),
.B2(n_220),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_2),
.A2(n_92),
.B1(n_130),
.B2(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_3),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_4),
.A2(n_90),
.B1(n_91),
.B2(n_96),
.Y(n_89)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_4),
.Y(n_96)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_6),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_6),
.Y(n_156)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_6),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_6),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_7),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_8),
.A2(n_38),
.B1(n_47),
.B2(n_52),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_8),
.A2(n_52),
.B1(n_125),
.B2(n_133),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_8),
.A2(n_52),
.B1(n_159),
.B2(n_162),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_8),
.A2(n_52),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_10),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_10),
.Y(n_183)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_10),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_10),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_10),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_11),
.A2(n_76),
.B1(n_80),
.B2(n_81),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_11),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_11),
.A2(n_80),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_12),
.A2(n_191),
.B1(n_195),
.B2(n_196),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_12),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_13),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_13),
.A2(n_43),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_13),
.A2(n_43),
.B1(n_159),
.B2(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_14),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_14),
.Y(n_110)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_14),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_14),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_232),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_230),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_163),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_18),
.B(n_163),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_99),
.C(n_137),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_19),
.A2(n_20),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_60),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_21),
.B(n_61),
.C(n_74),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_36),
.B(n_44),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_22),
.A2(n_36),
.B1(n_54),
.B2(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_22),
.B(n_46),
.Y(n_312)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_55),
.Y(n_54)
);

AO22x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_24),
.A2(n_48),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_26),
.Y(n_145)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_31),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_31),
.Y(n_125)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_31),
.Y(n_129)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_31),
.Y(n_135)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_41),
.Y(n_149)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_41),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_53),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_51),
.Y(n_168)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_51),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_53),
.A2(n_309),
.B(n_312),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_56),
.Y(n_153)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_74),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_62),
.B(n_180),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_SL g208 ( 
.A1(n_62),
.A2(n_179),
.B(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_62),
.A2(n_186),
.B(n_257),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_SL g309 ( 
.A1(n_62),
.A2(n_310),
.B(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_64),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_65),
.B(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_68),
.Y(n_175)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_84),
.B1(n_89),
.B2(n_97),
.Y(n_74)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_78),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_79),
.Y(n_194)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_84),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_84),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_84),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_85),
.Y(n_287)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_86),
.Y(n_296)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_89),
.Y(n_187)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_95),
.Y(n_285)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_97),
.Y(n_188)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_99),
.B(n_137),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_124),
.B(n_131),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_100),
.A2(n_131),
.B(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_100),
.A2(n_124),
.B1(n_223),
.B2(n_262),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_101),
.B(n_132),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_113),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_105),
.B1(n_108),
.B2(n_111),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g227 ( 
.A(n_103),
.Y(n_227)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_113),
.A2(n_228),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_126),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_129),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_129),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_129),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_136),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_154),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_138),
.B(n_154),
.Y(n_313)
);

AOI32xp33_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_141),
.A3(n_144),
.B1(n_146),
.B2(n_150),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx5_ASAP7_75t_SL g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_146),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_152),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B(n_157),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_157),
.A2(n_282),
.B(n_286),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_158),
.B(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_200),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_164)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_184),
.B2(n_185),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI32xp33_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.A3(n_171),
.B1(n_174),
.B2(n_179),
.Y(n_167)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_173),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_204)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_186),
.A2(n_254),
.B(n_257),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_194),
.Y(n_256)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_217),
.B2(n_229),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_208),
.B(n_210),
.Y(n_202)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_217),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B(n_228),
.Y(n_222)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_315),
.B(n_320),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_301),
.B(n_314),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_269),
.B(n_300),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_252),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_236),
.B(n_252),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_242),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_237),
.A2(n_242),
.B1(n_243),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_259),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_253),
.B(n_260),
.C(n_268),
.Y(n_302)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_254),
.Y(n_293)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_267),
.B2(n_268),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx11_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_290),
.B(n_299),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_280),
.B(n_289),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_279),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_277),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_288),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_288),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_297),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_297),
.Y(n_299)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_303),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_313),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_307),
.C(n_313),
.Y(n_316)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_316),
.B(n_317),
.Y(n_320)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);


endmodule