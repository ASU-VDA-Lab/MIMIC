module fake_jpeg_6395_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_21),
.B(n_23),
.C(n_20),
.Y(n_35)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_26),
.B(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_17),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_14),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_13),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_43),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_38),
.B1(n_40),
.B2(n_18),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_21),
.B1(n_20),
.B2(n_15),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_29),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_23),
.B1(n_15),
.B2(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_12),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_50),
.B(n_52),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_53),
.B(n_57),
.Y(n_65)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_60),
.C(n_61),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_46),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_37),
.C(n_36),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_71),
.C(n_49),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_36),
.C(n_35),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_78),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_60),
.B1(n_53),
.B2(n_59),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_22),
.B1(n_54),
.B2(n_30),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_51),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_71),
.A2(n_53),
.B(n_63),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_77),
.A2(n_79),
.B(n_80),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_25),
.C(n_30),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_22),
.Y(n_81)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_25),
.B1(n_31),
.B2(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_81),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_89),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_64),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_33),
.B(n_8),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_10),
.Y(n_95)
);

AOI322xp5_ASAP7_75t_SL g91 ( 
.A1(n_84),
.A2(n_85),
.A3(n_82),
.B1(n_87),
.B2(n_3),
.C1(n_4),
.C2(n_6),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_0),
.B(n_1),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_92),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_96),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_2),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_70),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_99),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_2),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_44),
.B(n_33),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_100),
.C(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_47),
.Y(n_104)
);


endmodule