module fake_jpeg_8305_n_278 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_278);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_37),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_15),
.B(n_26),
.Y(n_41)
);

OR2x2_ASAP7_75t_SL g74 ( 
.A(n_41),
.B(n_21),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_22),
.B1(n_15),
.B2(n_24),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_28),
.B1(n_22),
.B2(n_15),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_35),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_27),
.B1(n_21),
.B2(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_29),
.Y(n_72)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_51),
.B(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_58),
.B(n_66),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_67),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_28),
.B1(n_22),
.B2(n_36),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_68),
.B1(n_40),
.B2(n_43),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_69),
.B1(n_14),
.B2(n_20),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_37),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_37),
.B1(n_29),
.B2(n_20),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_18),
.B1(n_13),
.B2(n_21),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_32),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_88),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_35),
.C(n_31),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_83),
.C(n_90),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_61),
.B(n_33),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_86),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_35),
.C(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_35),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_35),
.C(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_31),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_101),
.B(n_102),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_58),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_106),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_65),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_81),
.C(n_78),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_76),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_113),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_71),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_25),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_66),
.B1(n_56),
.B2(n_46),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_110),
.A2(n_112),
.B1(n_27),
.B2(n_53),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_77),
.A2(n_64),
.B1(n_55),
.B2(n_38),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_79),
.B1(n_88),
.B2(n_78),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_47),
.B1(n_54),
.B2(n_55),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_71),
.Y(n_113)
);

OAI32xp33_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_27),
.A3(n_24),
.B1(n_33),
.B2(n_16),
.Y(n_114)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_63),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_115),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_60),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_33),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_96),
.B1(n_90),
.B2(n_91),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_140),
.B(n_104),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_129),
.B1(n_106),
.B2(n_100),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_93),
.B1(n_82),
.B2(n_80),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_125),
.B1(n_126),
.B2(n_117),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_116),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_122),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_89),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_87),
.C(n_52),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_86),
.B1(n_38),
.B2(n_95),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_95),
.B1(n_60),
.B2(n_49),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_128),
.A2(n_131),
.B(n_137),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_19),
.B1(n_13),
.B2(n_87),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_113),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_17),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_59),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_105),
.Y(n_147)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_136),
.Y(n_149)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_145),
.B1(n_159),
.B2(n_138),
.Y(n_166)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_146),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_130),
.A2(n_115),
.B1(n_97),
.B2(n_104),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_154),
.C(n_158),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_118),
.B(n_134),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_109),
.B(n_108),
.Y(n_150)
);

NOR4xp25_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_120),
.C(n_132),
.D(n_135),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_163),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_100),
.B1(n_111),
.B2(n_97),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_109),
.B1(n_102),
.B2(n_13),
.Y(n_153)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_157),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_48),
.C(n_33),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_127),
.A2(n_59),
.B1(n_14),
.B2(n_23),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_16),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_166),
.A2(n_16),
.B1(n_25),
.B2(n_17),
.Y(n_200)
);

AO21x1_ASAP7_75t_L g191 ( 
.A1(n_168),
.A2(n_170),
.B(n_164),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_162),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_171),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_156),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_122),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_181),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_127),
.B(n_131),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_176),
.B(n_23),
.Y(n_198)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_175),
.A2(n_186),
.B1(n_142),
.B2(n_160),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_143),
.A2(n_128),
.B1(n_59),
.B2(n_24),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_156),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_177),
.A2(n_183),
.B(n_169),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_143),
.A2(n_62),
.B1(n_23),
.B2(n_73),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_159),
.B1(n_155),
.B2(n_161),
.Y(n_192)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_48),
.C(n_62),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_154),
.C(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_167),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_190),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_200),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_141),
.B1(n_163),
.B2(n_157),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_189),
.A2(n_191),
.B1(n_192),
.B2(n_176),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_145),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_201),
.Y(n_211)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_199),
.B(n_177),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_48),
.C(n_62),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_62),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_203),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_62),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_186),
.Y(n_209)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_210),
.A2(n_25),
.B(n_1),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_218),
.Y(n_227)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_214),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_182),
.B1(n_165),
.B2(n_173),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_219),
.B1(n_7),
.B2(n_12),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_192),
.A2(n_165),
.B1(n_166),
.B2(n_173),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_216),
.A2(n_25),
.B1(n_17),
.B2(n_2),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_196),
.B1(n_180),
.B2(n_202),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_217),
.A2(n_188),
.B1(n_25),
.B2(n_8),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_198),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_193),
.A2(n_175),
.B1(n_181),
.B2(n_185),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_25),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_17),
.C(n_1),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_207),
.A2(n_203),
.B(n_201),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_223),
.Y(n_246)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_222),
.A2(n_8),
.B(n_12),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_229),
.C(n_233),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_6),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_11),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_231),
.Y(n_238)
);

NOR3xp33_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_11),
.C(n_10),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_208),
.C(n_220),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_212),
.C(n_11),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_235),
.A2(n_217),
.B1(n_212),
.B2(n_220),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_236),
.B(n_221),
.Y(n_243)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_229),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_228),
.B(n_10),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_17),
.C(n_1),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_0),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_256),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_254),
.C(n_239),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_241),
.A2(n_237),
.B1(n_223),
.B2(n_227),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_252),
.A2(n_254),
.B(n_17),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_224),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_232),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_242),
.B(n_226),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_257),
.A2(n_258),
.B(n_244),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_233),
.Y(n_258)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_260),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_262),
.B(n_264),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_253),
.A2(n_246),
.B(n_249),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_255),
.A2(n_245),
.B1(n_239),
.B2(n_247),
.Y(n_264)
);

OA21x2_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_9),
.B(n_10),
.Y(n_265)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_9),
.C(n_3),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_266),
.A2(n_252),
.B(n_3),
.Y(n_268)
);

NOR2x1_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_270),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_269),
.B(n_263),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_273),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_271),
.A3(n_267),
.B1(n_4),
.B2(n_5),
.C1(n_3),
.C2(n_2),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_275),
.A2(n_2),
.B(n_5),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_2),
.C(n_5),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_5),
.Y(n_278)
);


endmodule