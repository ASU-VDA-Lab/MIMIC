module fake_jpeg_26461_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_11),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_20),
.B(n_26),
.Y(n_31)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_23),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_19),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_17),
.C(n_15),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_37),
.Y(n_48)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR3xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_14),
.C(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_9),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_45),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_27),
.A2(n_22),
.B(n_12),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_25),
.B1(n_19),
.B2(n_18),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_25),
.B1(n_18),
.B2(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_54),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_6),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_36),
.C(n_44),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_53),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_36),
.B(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_56),
.Y(n_67)
);

OAI321xp33_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_64),
.A3(n_63),
.B1(n_13),
.B2(n_12),
.C(n_8),
.Y(n_70)
);

AO221x1_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_45),
.B1(n_37),
.B2(n_12),
.C(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_71),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_7),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_72),
.A2(n_69),
.B(n_8),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_74),
.B(n_13),
.C(n_12),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_13),
.B(n_71),
.Y(n_77)
);


endmodule