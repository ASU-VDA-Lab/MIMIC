module fake_jpeg_9315_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_12),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_35),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_24),
.Y(n_43)
);

AO22x1_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_22),
.B1(n_21),
.B2(n_20),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_26),
.Y(n_39)
);

INVxp33_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_29),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_22),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_22),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_35),
.B1(n_31),
.B2(n_25),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_46),
.B(n_37),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_34),
.B(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_36),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_50),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_51),
.C(n_19),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_36),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_55),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_58),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_33),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_25),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_49),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_33),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_52),
.B1(n_9),
.B2(n_17),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_62),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_16),
.C(n_11),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_16),
.C(n_13),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NAND4xp25_ASAP7_75t_SL g66 ( 
.A(n_64),
.B(n_13),
.C(n_9),
.D(n_11),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_66),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_68),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_60),
.B1(n_62),
.B2(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_61),
.Y(n_72)
);

AOI322xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_73),
.A3(n_70),
.B1(n_71),
.B2(n_6),
.C1(n_8),
.C2(n_2),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_67),
.C(n_5),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

AOI322xp5_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_0),
.A3(n_1),
.B1(n_4),
.B2(n_6),
.C1(n_8),
.C2(n_64),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_76),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_75),
.Y(n_78)
);


endmodule