module fake_jpeg_5396_n_257 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_225;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_7),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_36),
.B(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_38),
.B(n_40),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_23),
.B(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_39),
.B(n_21),
.Y(n_77)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_15),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_20),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_48),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_45),
.Y(n_96)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_46),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_8),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_47),
.B(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_13),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_27),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_55),
.Y(n_102)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_18),
.B1(n_29),
.B2(n_32),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_54),
.A2(n_75),
.B1(n_83),
.B2(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_47),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_59),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_15),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_79),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_66),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_31),
.B1(n_23),
.B2(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_63),
.A2(n_72),
.B1(n_82),
.B2(n_98),
.Y(n_112)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_31),
.B1(n_29),
.B2(n_33),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_74),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_40),
.A2(n_33),
.B1(n_21),
.B2(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_78),
.Y(n_116)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_22),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_39),
.A2(n_26),
.B1(n_16),
.B2(n_25),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_80),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_34),
.B1(n_16),
.B2(n_25),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_22),
.B1(n_25),
.B2(n_24),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_36),
.B(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_22),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_89),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_35),
.B(n_27),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_50),
.B(n_22),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_16),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_93),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_45),
.B(n_30),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_39),
.B(n_30),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_42),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_24),
.B1(n_9),
.B2(n_10),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_30),
.B(n_25),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_114),
.B(n_120),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_55),
.A2(n_51),
.B(n_58),
.C(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_108),
.B(n_123),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_64),
.B1(n_78),
.B2(n_84),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_30),
.B1(n_24),
.B2(n_2),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_114),
.A2(n_61),
.B1(n_76),
.B2(n_52),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_24),
.B(n_1),
.C(n_2),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_0),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_60),
.B1(n_87),
.B2(n_76),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_81),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_130),
.B(n_135),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_134),
.B1(n_154),
.B2(n_157),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_69),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_145),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_99),
.C(n_62),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_141),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_116),
.B(n_53),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_136),
.Y(n_166)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_73),
.B1(n_64),
.B2(n_71),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_104),
.A2(n_119),
.B1(n_53),
.B2(n_112),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_139),
.A2(n_142),
.B1(n_123),
.B2(n_113),
.Y(n_180)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_94),
.C(n_86),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_68),
.C(n_91),
.Y(n_143)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_143),
.B(n_152),
.CI(n_107),
.CON(n_161),
.SN(n_161)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_110),
.B(n_67),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_151),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_106),
.A2(n_65),
.B1(n_59),
.B2(n_56),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_149),
.A2(n_126),
.B1(n_115),
.B2(n_103),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_70),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_156),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_66),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_88),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_95),
.Y(n_153)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_108),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_9),
.Y(n_155)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_125),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_12),
.Y(n_159)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_161),
.B(n_177),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_120),
.B(n_118),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_168),
.A2(n_156),
.B(n_145),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_118),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_177),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_107),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_179),
.Y(n_188)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_184),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_101),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_185),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_128),
.B(n_101),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_182),
.B(n_187),
.Y(n_203)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_129),
.B(n_125),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_141),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_202),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_158),
.B(n_139),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_195),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_147),
.B(n_133),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_205),
.B(n_209),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_143),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_161),
.Y(n_213)
);

NAND2xp67_ASAP7_75t_SL g197 ( 
.A(n_168),
.B(n_147),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_198),
.B(n_171),
.Y(n_212)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_207),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_134),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_201),
.A2(n_169),
.B(n_166),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_157),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_111),
.B(n_103),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_146),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_208),
.C(n_162),
.Y(n_211)
);

INVxp33_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_122),
.C(n_121),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_122),
.B(n_121),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_206),
.C(n_208),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_198),
.B1(n_178),
.B2(n_204),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_214),
.A2(n_216),
.B1(n_217),
.B2(n_220),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_171),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_160),
.B1(n_184),
.B2(n_164),
.Y(n_217)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_193),
.B(n_162),
.CI(n_160),
.CON(n_219),
.SN(n_219)
);

OAI321xp33_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_223),
.A3(n_224),
.B1(n_201),
.B2(n_209),
.C(n_203),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_166),
.B1(n_182),
.B2(n_169),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_191),
.B(n_180),
.Y(n_223)
);

OAI321xp33_ASAP7_75t_L g224 ( 
.A1(n_197),
.A2(n_173),
.A3(n_167),
.B1(n_174),
.B2(n_126),
.C(n_111),
.Y(n_224)
);

XOR2x2_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_167),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_221),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_228),
.C(n_230),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_196),
.C(n_190),
.Y(n_228)
);

AOI321xp33_ASAP7_75t_L g240 ( 
.A1(n_229),
.A2(n_221),
.A3(n_222),
.B1(n_219),
.B2(n_218),
.C(n_224),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_190),
.C(n_189),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_223),
.A2(n_201),
.B1(n_191),
.B2(n_202),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_231),
.A2(n_234),
.B1(n_212),
.B2(n_210),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_233),
.B(n_215),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_174),
.B(n_170),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_163),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_226),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_240),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_239),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_232),
.B1(n_234),
.B2(n_228),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_238),
.B(n_186),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_242),
.Y(n_245)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_245),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_241),
.A2(n_239),
.B(n_238),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_246),
.A2(n_247),
.B(n_249),
.Y(n_250)
);

AOI31xp67_ASAP7_75t_SL g247 ( 
.A1(n_244),
.A2(n_12),
.A3(n_5),
.B(n_6),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_186),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_109),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_246),
.A2(n_137),
.B(n_140),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_4),
.C(n_250),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_144),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_255),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_253),
.Y(n_257)
);


endmodule