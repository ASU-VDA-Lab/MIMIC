module fake_jpeg_7138_n_274 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_274);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_220;
wire n_74;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx12f_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_41),
.B(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_6),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_50),
.Y(n_70)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_24),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_47),
.B(n_52),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_24),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_53),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_31),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_37),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_34),
.A2(n_19),
.B1(n_30),
.B2(n_26),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_16),
.B1(n_21),
.B2(n_25),
.Y(n_83)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_37),
.C(n_15),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_40),
.B(n_38),
.C(n_36),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_71),
.B1(n_86),
.B2(n_23),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_40),
.B(n_38),
.C(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_30),
.B1(n_27),
.B2(n_64),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_19),
.B1(n_27),
.B2(n_18),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_81),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_19),
.B1(n_18),
.B2(n_20),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_56),
.A2(n_20),
.B1(n_26),
.B2(n_21),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_85),
.B1(n_29),
.B2(n_57),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_51),
.B1(n_52),
.B2(n_46),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_25),
.B1(n_16),
.B2(n_57),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_40),
.B1(n_38),
.B2(n_29),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_55),
.Y(n_98)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_92),
.Y(n_118)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_93),
.A2(n_88),
.B1(n_107),
.B2(n_108),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

FAx1_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_48),
.CI(n_53),
.CON(n_95),
.SN(n_95)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_100),
.C(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_97),
.Y(n_124)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_99),
.A2(n_106),
.B1(n_109),
.B2(n_65),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_46),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_70),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_76),
.B1(n_66),
.B2(n_65),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_11),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_0),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_37),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_111),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_55),
.B1(n_37),
.B2(n_32),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_55),
.B1(n_37),
.B2(n_23),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_0),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_10),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_63),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_112),
.A2(n_114),
.B1(n_92),
.B2(n_66),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_89),
.A2(n_65),
.B1(n_73),
.B2(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_103),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_121),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_126),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_70),
.C(n_73),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_109),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_122),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_87),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_91),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_67),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_123),
.A2(n_135),
.B(n_1),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_67),
.B(n_65),
.C(n_63),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_134),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_97),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_97),
.B1(n_90),
.B2(n_82),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_60),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_106),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_89),
.A2(n_0),
.B(n_1),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_95),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_159),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_142),
.B(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_147),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_94),
.Y(n_144)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_151),
.C(n_119),
.Y(n_162)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_101),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_150),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_94),
.Y(n_149)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_131),
.B(n_110),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_104),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_128),
.B1(n_113),
.B2(n_129),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_156),
.B(n_129),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_112),
.B1(n_123),
.B2(n_114),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_131),
.B(n_1),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_134),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_90),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_82),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_158),
.B(n_118),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_115),
.B(n_121),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_149),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_160),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_145),
.C(n_159),
.Y(n_193)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_165),
.B(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_169),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_117),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_170),
.B(n_136),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_152),
.A2(n_128),
.B1(n_130),
.B2(n_133),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_176),
.B1(n_182),
.B2(n_140),
.Y(n_199)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_174),
.B(n_177),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_138),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_155),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_123),
.Y(n_181)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_148),
.A2(n_117),
.B1(n_135),
.B2(n_127),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_169),
.A2(n_173),
.B1(n_170),
.B2(n_160),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_198),
.Y(n_205)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_192),
.Y(n_209)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_136),
.C(n_171),
.Y(n_204)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_127),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_196),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_151),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_143),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_162),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_146),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_172),
.Y(n_208)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_202),
.B1(n_147),
.B2(n_166),
.Y(n_213)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_204),
.C(n_211),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_182),
.B1(n_140),
.B2(n_154),
.Y(n_206)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_187),
.A2(n_174),
.B1(n_181),
.B2(n_163),
.Y(n_207)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_213),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_161),
.C(n_166),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_214),
.C(n_186),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_156),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_150),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_180),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_216),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_196),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_164),
.B1(n_141),
.B2(n_168),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_219),
.B(n_191),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_210),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_224),
.A2(n_226),
.B(n_232),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_217),
.A2(n_183),
.B(n_200),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_198),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_10),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_229),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_SL g229 ( 
.A(n_218),
.B(n_201),
.C(n_192),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_217),
.B(n_188),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_204),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_188),
.C(n_202),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_164),
.B1(n_167),
.B2(n_185),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_205),
.Y(n_238)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_239),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_194),
.Y(n_236)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_240),
.C(n_242),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_221),
.B(n_212),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_245),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_190),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_227),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_244),
.Y(n_250)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g246 ( 
.A(n_242),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_7),
.Y(n_257)
);

NAND4xp25_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_232),
.C(n_223),
.D(n_225),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_254),
.B(n_60),
.Y(n_260)
);

OAI321xp33_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_11),
.A3(n_14),
.B1(n_12),
.B2(n_9),
.C(n_5),
.Y(n_251)
);

OAI21x1_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_9),
.B(n_14),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_74),
.C(n_82),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_248),
.A2(n_234),
.B1(n_241),
.B2(n_74),
.Y(n_255)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_255),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_256),
.B(n_258),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_12),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_5),
.B(n_12),
.C(n_11),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_60),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_260),
.C(n_261),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_249),
.B(n_1),
.Y(n_261)
);

NAND4xp25_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_254),
.C(n_252),
.D(n_4),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_266),
.C(n_2),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_262),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_63),
.B(n_3),
.Y(n_269)
);

AOI31xp33_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_264),
.A3(n_3),
.B(n_4),
.Y(n_270)
);

AOI211xp5_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_264),
.B(n_3),
.C(n_2),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_271),
.C(n_2),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_3),
.Y(n_274)
);


endmodule