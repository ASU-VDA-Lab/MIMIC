module real_jpeg_1644_n_30 (n_17, n_8, n_0, n_21, n_2, n_29, n_180, n_10, n_175, n_9, n_178, n_12, n_24, n_170, n_176, n_6, n_28, n_171, n_177, n_179, n_23, n_11, n_14, n_172, n_25, n_7, n_22, n_18, n_3, n_174, n_5, n_4, n_173, n_1, n_26, n_27, n_20, n_19, n_16, n_15, n_13, n_30);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_29;
input n_180;
input n_10;
input n_175;
input n_9;
input n_178;
input n_12;
input n_24;
input n_170;
input n_176;
input n_6;
input n_28;
input n_171;
input n_177;
input n_179;
input n_23;
input n_11;
input n_14;
input n_172;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_174;
input n_5;
input n_4;
input n_173;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_30;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_150;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

AND2x2_ASAP7_75t_L g80 ( 
.A(n_0),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_2),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_3),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_4),
.B(n_73),
.C(n_98),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_5),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_6),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_7),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_8),
.A2(n_34),
.B1(n_146),
.B2(n_148),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_8),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_8),
.B(n_36),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_8),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_8),
.B(n_154),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_8),
.A2(n_141),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_9),
.B(n_54),
.Y(n_139)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_10),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_11),
.B(n_75),
.C(n_90),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g83 ( 
.A(n_13),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

BUFx16f_ASAP7_75t_L g92 ( 
.A(n_13),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_14),
.A2(n_71),
.B1(n_104),
.B2(n_107),
.Y(n_70)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_14),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_15),
.B(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_15),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_17),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_18),
.A2(n_76),
.B1(n_78),
.B2(n_89),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_19),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_20),
.A2(n_80),
.B(n_84),
.Y(n_79)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_22),
.Y(n_144)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_25),
.B(n_66),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_26),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_27),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_28),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_163),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_157),
.B(n_162),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_153),
.B(n_156),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_43),
.B(n_145),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_39),
.B(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_39),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_39),
.B(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_39),
.Y(n_152)
);

BUFx4f_ASAP7_75t_SL g161 ( 
.A(n_39),
.Y(n_161)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx6p67_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_77),
.Y(n_76)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_42),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_42),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_141),
.C(n_142),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_51),
.B(n_140),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_46),
.B(n_50),
.Y(n_140)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_49),
.B(n_155),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B(n_56),
.C(n_139),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_135),
.C(n_136),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_64),
.B(n_134),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_59),
.B(n_63),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_103),
.Y(n_102)
);

OAI221xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_69),
.B1(n_70),
.B2(n_110),
.C(n_124),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_100),
.C(n_101),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_93),
.C(n_94),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_87),
.C(n_88),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_87),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_84),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_119),
.Y(n_110)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_125),
.A3(n_126),
.B1(n_129),
.B2(n_130),
.C1(n_133),
.C2(n_180),
.Y(n_124)
);

NOR3xp33_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_113),
.C(n_116),
.Y(n_111)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_141),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_158),
.Y(n_162)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

BUFx4f_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_170),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_171),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_172),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_173),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_174),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_175),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_176),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_177),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_178),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_179),
.Y(n_123)
);


endmodule