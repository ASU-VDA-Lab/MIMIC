module fake_jpeg_26404_n_67 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_67);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_67;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;
wire n_66;

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_0),
.B(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g37 ( 
.A1(n_24),
.A2(n_7),
.B1(n_30),
.B2(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_40),
.Y(n_54)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_23),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_45),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_56),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_54),
.A2(n_51),
.B1(n_37),
.B2(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_49),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_44),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_58),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_60),
.A2(n_48),
.B(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_61),
.B(n_62),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_60),
.A2(n_50),
.B1(n_52),
.B2(n_42),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

BUFx24_ASAP7_75t_SL g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_66),
.B(n_46),
.Y(n_67)
);


endmodule