module real_jpeg_23470_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_288;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_249;
wire n_286;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_1),
.A2(n_70),
.B(n_158),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_1),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_1),
.B(n_58),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_L g226 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_160),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_1),
.B(n_29),
.C(n_46),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_1),
.B(n_79),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_1),
.A2(n_94),
.B1(n_245),
.B2(n_252),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g61 ( 
.A(n_4),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_5),
.A2(n_71),
.B1(n_75),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_5),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_5),
.A2(n_59),
.B1(n_62),
.B2(n_116),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_116),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_5),
.A2(n_29),
.B1(n_31),
.B2(n_116),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_6),
.A2(n_30),
.B1(n_70),
.B2(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_6),
.A2(n_30),
.B1(n_59),
.B2(n_62),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_6),
.A2(n_30),
.B1(n_41),
.B2(n_42),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_7),
.A2(n_29),
.B1(n_31),
.B2(n_52),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_7),
.A2(n_52),
.B1(n_59),
.B2(n_62),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_10),
.A2(n_65),
.B1(n_75),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_10),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_10),
.A2(n_59),
.B1(n_62),
.B2(n_163),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_163),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_10),
.A2(n_29),
.B1(n_31),
.B2(n_163),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_11),
.A2(n_43),
.B1(n_59),
.B2(n_62),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_11),
.A2(n_29),
.B1(n_31),
.B2(n_43),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_13),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_13),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_13),
.A2(n_59),
.B1(n_62),
.B2(n_68),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_68),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_13),
.A2(n_29),
.B1(n_31),
.B2(n_68),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_14),
.A2(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_14),
.A2(n_34),
.B1(n_59),
.B2(n_62),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_14),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_14),
.A2(n_34),
.B1(n_65),
.B2(n_75),
.Y(n_134)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_15),
.Y(n_246)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_15),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_143),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_141),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_117),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_19),
.B(n_117),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_87),
.C(n_99),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_20),
.A2(n_21),
.B1(n_87),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_22),
.B(n_55),
.C(n_76),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_23),
.A2(n_24),
.B1(n_37),
.B2(n_38),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_32),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_25),
.A2(n_94),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_29),
.A2(n_31),
.B1(n_46),
.B2(n_48),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_31),
.B(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_32),
.A2(n_179),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_33),
.B(n_36),
.Y(n_104)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_35),
.A2(n_103),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_35),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_50),
.B2(n_51),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_40),
.A2(n_49),
.B(n_106),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_42),
.B1(n_46),
.B2(n_48),
.Y(n_45)
);

AO22x1_ASAP7_75t_L g79 ( 
.A1(n_41),
.A2(n_42),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_41),
.B(n_81),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_42),
.A2(n_62),
.A3(n_80),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_42),
.B(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_44),
.A2(n_51),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_44),
.B(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_44),
.A2(n_90),
.B(n_125),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_44),
.A2(n_50),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_44),
.A2(n_123),
.B(n_209),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_44),
.A2(n_50),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_44),
.A2(n_50),
.B1(n_208),
.B2(n_227),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_49),
.B(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_49),
.B(n_160),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_76),
.B2(n_77),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_67),
.B(n_73),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_56),
.A2(n_58),
.B1(n_67),
.B2(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_56),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_56),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_56),
.A2(n_58),
.B1(n_115),
.B2(n_162),
.Y(n_169)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_64),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_57),
.B(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_57),
.A2(n_156),
.B1(n_157),
.B2(n_161),
.Y(n_155)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_59),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_62),
.B1(n_80),
.B2(n_81),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_59),
.A2(n_63),
.B(n_159),
.C(n_175),
.Y(n_174)
);

HAxp5_ASAP7_75t_SL g203 ( 
.A(n_59),
.B(n_160),
.CON(n_203),
.SN(n_203)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_61),
.B(n_62),
.C(n_72),
.Y(n_175)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_66),
.B(n_160),
.Y(n_159)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_82),
.B(n_83),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_78),
.A2(n_82),
.B1(n_112),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_78),
.A2(n_112),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_78),
.A2(n_112),
.B1(n_153),
.B2(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_79),
.B(n_86),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_79),
.B(n_111),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_79),
.A2(n_84),
.B1(n_194),
.B2(n_203),
.Y(n_206)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_87),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_92),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_93),
.B1(n_131),
.B2(n_135),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B(n_98),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_94),
.A2(n_98),
.B(n_104),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_94),
.A2(n_95),
.B1(n_242),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_97),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_99),
.B(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_108),
.C(n_114),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_100),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_105),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_108),
.A2(n_109),
.B1(n_114),
.B2(n_280),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_112),
.B(n_113),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_112),
.A2(n_154),
.B(n_172),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_114),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_139),
.B2(n_140),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_129),
.B1(n_137),
.B2(n_138),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_126),
.B(n_128),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_126),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_136),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_284),
.B(n_289),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_195),
.B(n_272),
.C(n_283),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_181),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_181),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_166),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_164),
.B2(n_165),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_148),
.B(n_165),
.C(n_166),
.Y(n_273)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_155),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_184),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_155),
.B(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_160),
.B(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_173),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_169),
.B(n_170),
.C(n_173),
.Y(n_281)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_176),
.B1(n_177),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.C(n_187),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_182),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_185),
.B(n_187),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_192),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_190),
.B1(n_191),
.B2(n_214),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_188),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_267),
.B(n_271),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_221),
.B(n_266),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_210),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_200),
.B(n_210),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_206),
.C(n_207),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_201),
.B(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_205),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_206),
.B(n_207),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_215),
.B2(n_216),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_211),
.B(n_218),
.C(n_220),
.Y(n_268)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_217),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_261),
.B(n_265),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_238),
.B(n_260),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_230),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_224),
.B(n_230),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_228),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_235),
.C(n_236),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_234),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_248),
.B(n_259),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_247),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_247),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_253),
.B(n_258),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_250),
.B(n_251),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_262),
.B(n_263),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_274),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_281),
.B2(n_282),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_278),
.C(n_282),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_281),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);


endmodule