module fake_jpeg_22833_n_32 (n_3, n_2, n_1, n_0, n_4, n_32);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_32;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx13_ASAP7_75t_L g5 ( 
.A(n_2),
.Y(n_5)
);

INVx3_ASAP7_75t_SL g6 ( 
.A(n_1),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

BUFx10_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_7),
.B(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_9),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_12),
.A2(n_14),
.B1(n_6),
.B2(n_5),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_0),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_6),
.A2(n_9),
.B1(n_5),
.B2(n_3),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_6),
.C(n_8),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_11),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_16),
.A2(n_9),
.B1(n_11),
.B2(n_3),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_18),
.A2(n_13),
.B(n_12),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_22),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_21),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_25),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_24),
.A2(n_16),
.B1(n_8),
.B2(n_4),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_24),
.B1(n_27),
.B2(n_8),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_27),
.B(n_8),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_29),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_29),
.B(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_4),
.Y(n_32)
);


endmodule