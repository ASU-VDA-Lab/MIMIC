module fake_ariane_606_n_1863 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_172, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1863);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1863;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_15),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_31),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_165),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_9),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_67),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_59),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_90),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_81),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_6),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_116),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_96),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_7),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_157),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_15),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_43),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_144),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_86),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_42),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_18),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_38),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_78),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_71),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_139),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_82),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_72),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_146),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_99),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_80),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_102),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_20),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_25),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_62),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_33),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_47),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_79),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_100),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_28),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_88),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_91),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_138),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_110),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_38),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_6),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_11),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_137),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_147),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_69),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_135),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_19),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_106),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_160),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_9),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_127),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_18),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_34),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_141),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_51),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_117),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_43),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_151),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_149),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_159),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_109),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_1),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_108),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_140),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_112),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_64),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_12),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_53),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_118),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_85),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_56),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_107),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_129),
.Y(n_256)
);

BUFx2_ASAP7_75t_SL g257 ( 
.A(n_105),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_56),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_52),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_46),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_40),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_130),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_83),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_23),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_2),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_89),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_47),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_39),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_154),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_8),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_122),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_17),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_155),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_60),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_115),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_3),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_8),
.Y(n_277)
);

BUFx5_ASAP7_75t_L g278 ( 
.A(n_62),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_16),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_143),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_49),
.Y(n_281)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_142),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_30),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_93),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_168),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_51),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_84),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_68),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_5),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_113),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_163),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_21),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_31),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_2),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_104),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_19),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_14),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_30),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_145),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_75),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_60),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_14),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_26),
.Y(n_303)
);

BUFx2_ASAP7_75t_SL g304 ( 
.A(n_5),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_125),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_33),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_70),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_1),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_134),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_32),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_87),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_3),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_37),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_54),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_103),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_50),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_28),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_119),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_4),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_52),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_59),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_66),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_169),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_162),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_136),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_57),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_55),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_7),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_153),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_120),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_76),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_25),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_10),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_21),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_114),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_4),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_10),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_97),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_121),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_57),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_46),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_50),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_27),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_36),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_98),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_20),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_22),
.Y(n_347)
);

NOR2xp67_ASAP7_75t_L g348 ( 
.A(n_292),
.B(n_0),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_340),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_278),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_278),
.B(n_0),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_220),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_279),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_278),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_278),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_278),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_239),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_R g358 ( 
.A(n_237),
.B(n_123),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_278),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_278),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_278),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_333),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_333),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_242),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_230),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_233),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_333),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_333),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_261),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_236),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_261),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_333),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_189),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_195),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_333),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_223),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_208),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_209),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_187),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_194),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_210),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_238),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_246),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_219),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_250),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_258),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_223),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_283),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_246),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_283),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_288),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_288),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_261),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_240),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_317),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_267),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_281),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_277),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_317),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_320),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_221),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_320),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_245),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_249),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_327),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_181),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_251),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_181),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_285),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_319),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_198),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_198),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_305),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_174),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_206),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_259),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_175),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_260),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_206),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_264),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_213),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_205),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_175),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_213),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_265),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_226),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_176),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_270),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_226),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_289),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_272),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_350),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_354),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_417),
.B(n_315),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_350),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_354),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_355),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_358),
.B(n_188),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_355),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_401),
.B(n_292),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_417),
.B(n_188),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_433),
.B(n_296),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_376),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_400),
.A2(n_347),
.B1(n_346),
.B2(n_328),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_376),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_356),
.B(n_184),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_356),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_297),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_359),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_359),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_360),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_360),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_361),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_361),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_362),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_362),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_363),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_363),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_367),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_351),
.B(n_266),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_367),
.B(n_192),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_368),
.Y(n_465)
);

OA21x2_ASAP7_75t_L g466 ( 
.A1(n_409),
.A2(n_204),
.B(n_193),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_368),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_372),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_372),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_413),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_373),
.B(n_216),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_373),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_377),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_377),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_409),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_411),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_411),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_365),
.Y(n_478)
);

BUFx8_ASAP7_75t_L g479 ( 
.A(n_414),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_414),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_415),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_415),
.B(n_218),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_418),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_348),
.B(n_366),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_418),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_422),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_353),
.B(n_207),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_422),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_424),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_424),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_379),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_427),
.Y(n_492)
);

NAND2x1p5_ASAP7_75t_L g493 ( 
.A(n_427),
.B(n_266),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_429),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_429),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_432),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_432),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_378),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_378),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_389),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_389),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_381),
.B(n_301),
.Y(n_502)
);

BUFx12f_ASAP7_75t_L g503 ( 
.A(n_370),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_390),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_390),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_382),
.B(n_222),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_392),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_392),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_397),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_397),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_402),
.B(n_303),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_478),
.B(n_384),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_450),
.Y(n_513)
);

CKINVDCx11_ASAP7_75t_R g514 ( 
.A(n_503),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_444),
.B(n_383),
.Y(n_515)
);

BUFx4f_ASAP7_75t_L g516 ( 
.A(n_466),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_450),
.Y(n_517)
);

OR2x6_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_304),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_444),
.A2(n_425),
.B1(n_412),
.B2(n_416),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_450),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_470),
.Y(n_521)
);

INVx5_ASAP7_75t_L g522 ( 
.A(n_463),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_462),
.B(n_396),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_462),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_450),
.Y(n_525)
);

BUFx4f_ASAP7_75t_L g526 ( 
.A(n_466),
.Y(n_526)
);

OR2x6_ASAP7_75t_L g527 ( 
.A(n_503),
.B(n_444),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_454),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_462),
.B(n_405),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_454),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_454),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_462),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_L g533 ( 
.A(n_463),
.B(n_406),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_463),
.Y(n_534)
);

NOR2x1p5_ASAP7_75t_L g535 ( 
.A(n_503),
.B(n_352),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_454),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_479),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_455),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_462),
.B(n_410),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_455),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_462),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_435),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_455),
.Y(n_543)
);

INVx3_ASAP7_75t_SL g544 ( 
.A(n_487),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_455),
.Y(n_545)
);

NAND3xp33_ASAP7_75t_L g546 ( 
.A(n_436),
.B(n_316),
.C(n_310),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_478),
.B(n_419),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_443),
.B(n_421),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_456),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_491),
.B(n_374),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_456),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_456),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_456),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_460),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g555 ( 
.A(n_479),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_458),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_441),
.B(n_423),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_447),
.A2(n_235),
.B1(n_254),
.B2(n_430),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_463),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_460),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_441),
.B(n_428),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_484),
.B(n_431),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_484),
.B(n_434),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_444),
.A2(n_403),
.B1(n_394),
.B2(n_393),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_443),
.B(n_369),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_479),
.Y(n_566)
);

OAI22xp33_ASAP7_75t_L g567 ( 
.A1(n_447),
.A2(n_371),
.B1(n_426),
.B2(n_420),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_435),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_457),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_463),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_457),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_457),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_457),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_444),
.B(n_448),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_469),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_491),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_439),
.B(n_385),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_469),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_469),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_SL g580 ( 
.A1(n_487),
.A2(n_349),
.B1(n_357),
.B2(n_364),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_469),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_472),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_487),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_439),
.B(n_391),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_437),
.B(n_386),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_470),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_472),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_472),
.Y(n_588)
);

AND2x2_ASAP7_75t_SL g589 ( 
.A(n_466),
.B(n_266),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_472),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_474),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_474),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_474),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_444),
.B(n_177),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_474),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_479),
.A2(n_332),
.B1(n_334),
.B2(n_336),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_448),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_436),
.B(n_341),
.C(n_322),
.Y(n_598)
);

NAND3xp33_ASAP7_75t_L g599 ( 
.A(n_436),
.B(n_294),
.C(n_229),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_448),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_440),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_448),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_479),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_460),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_435),
.Y(n_605)
);

CKINVDCx16_ASAP7_75t_R g606 ( 
.A(n_502),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_440),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_437),
.B(n_387),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_460),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_502),
.B(n_388),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_440),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_L g612 ( 
.A1(n_506),
.A2(n_211),
.B1(n_196),
.B2(n_190),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_479),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_460),
.Y(n_614)
);

NAND3xp33_ASAP7_75t_L g615 ( 
.A(n_442),
.B(n_231),
.C(n_227),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_442),
.B(n_398),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_442),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_452),
.B(n_399),
.Y(n_618)
);

BUFx4f_ASAP7_75t_L g619 ( 
.A(n_466),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_452),
.B(n_185),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_473),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_445),
.B(n_402),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_473),
.Y(n_623)
);

INVxp33_ASAP7_75t_L g624 ( 
.A(n_445),
.Y(n_624)
);

AND2x2_ASAP7_75t_SL g625 ( 
.A(n_466),
.B(n_266),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_452),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_453),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_502),
.A2(n_176),
.B1(n_214),
.B2(n_211),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_502),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_473),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_453),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_453),
.B(n_395),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_463),
.Y(n_633)
);

NOR2x1p5_ASAP7_75t_L g634 ( 
.A(n_445),
.B(n_178),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_459),
.B(n_461),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_459),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_466),
.Y(n_637)
);

INVx4_ASAP7_75t_SL g638 ( 
.A(n_463),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_459),
.B(n_199),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_461),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_502),
.A2(n_217),
.B1(n_256),
.B2(n_408),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_461),
.B(n_266),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_502),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_451),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_473),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_463),
.A2(n_408),
.B1(n_407),
.B2(n_404),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_473),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_458),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_465),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_463),
.A2(n_407),
.B1(n_404),
.B2(n_257),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_458),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_465),
.B(n_177),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_458),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_465),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_506),
.B(n_182),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_467),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_463),
.A2(n_274),
.B1(n_276),
.B2(n_286),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_451),
.B(n_178),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_468),
.A2(n_326),
.B1(n_196),
.B2(n_190),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_451),
.B(n_179),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_468),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_585),
.B(n_608),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_606),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_644),
.B(n_468),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_644),
.B(n_485),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_576),
.B(n_511),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_577),
.B(n_375),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_597),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_597),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_611),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_584),
.B(n_544),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_596),
.A2(n_463),
.B1(n_486),
.B2(n_464),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_L g673 ( 
.A(n_632),
.B(n_464),
.C(n_449),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_544),
.B(n_380),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_548),
.B(n_485),
.Y(n_675)
);

OAI22xp33_ASAP7_75t_L g676 ( 
.A1(n_606),
.A2(n_268),
.B1(n_179),
.B2(n_326),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_583),
.B(n_565),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_SL g678 ( 
.A(n_643),
.B(n_449),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_643),
.B(n_485),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_600),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_565),
.B(n_511),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_516),
.B(n_458),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_516),
.B(n_458),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_516),
.B(n_458),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_521),
.B(n_511),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_521),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_600),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_617),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_L g689 ( 
.A(n_613),
.B(n_458),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_526),
.B(n_471),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_526),
.B(n_435),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_616),
.B(n_485),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_601),
.Y(n_693)
);

O2A1O1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_635),
.A2(n_480),
.B(n_490),
.C(n_483),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_544),
.B(n_482),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_629),
.B(n_476),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_601),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_629),
.B(n_476),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_574),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_620),
.B(n_476),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_557),
.B(n_486),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_526),
.B(n_435),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_639),
.B(n_477),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_550),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_562),
.B(n_622),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_619),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_607),
.Y(n_707)
);

NAND2xp33_ASAP7_75t_SL g708 ( 
.A(n_535),
.B(n_180),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_622),
.B(n_477),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_515),
.B(n_477),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_619),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_515),
.B(n_480),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_613),
.B(n_537),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_574),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_515),
.B(n_480),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_515),
.B(n_483),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_619),
.B(n_435),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_607),
.Y(n_718)
);

NAND2xp33_ASAP7_75t_L g719 ( 
.A(n_537),
.B(n_435),
.Y(n_719)
);

NAND2x1p5_ASAP7_75t_L g720 ( 
.A(n_534),
.B(n_490),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_554),
.B(n_435),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_602),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_554),
.B(n_560),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_586),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_554),
.B(n_492),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_586),
.B(n_498),
.Y(n_726)
);

NOR2xp67_ASAP7_75t_L g727 ( 
.A(n_615),
.B(n_492),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_560),
.B(n_438),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_626),
.Y(n_729)
);

NOR2xp67_ASAP7_75t_SL g730 ( 
.A(n_566),
.B(n_180),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_560),
.B(n_438),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_614),
.B(n_524),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_614),
.B(n_510),
.Y(n_733)
);

NAND2x1_ASAP7_75t_L g734 ( 
.A(n_534),
.B(n_438),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_624),
.B(n_498),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_614),
.B(n_510),
.Y(n_736)
);

NOR2xp67_ASAP7_75t_L g737 ( 
.A(n_615),
.B(n_482),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_523),
.B(n_498),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_558),
.A2(n_518),
.B1(n_527),
.B2(n_610),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_512),
.B(n_183),
.Y(n_740)
);

OR2x6_ASAP7_75t_L g741 ( 
.A(n_527),
.B(n_499),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_626),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_602),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_529),
.B(n_499),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_539),
.B(n_499),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_517),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_524),
.B(n_438),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_604),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_524),
.B(n_438),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_542),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_L g751 ( 
.A(n_566),
.B(n_438),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_547),
.B(n_214),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_517),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_532),
.B(n_504),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_550),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_L g756 ( 
.A(n_603),
.B(n_438),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_520),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_532),
.B(n_504),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_574),
.A2(n_318),
.B1(n_191),
.B2(n_197),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_627),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_520),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_660),
.B(n_504),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_657),
.B(n_308),
.C(n_268),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_631),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_525),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_532),
.B(n_438),
.Y(n_766)
);

BUFx8_ASAP7_75t_L g767 ( 
.A(n_660),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_631),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_541),
.B(n_510),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_541),
.B(n_508),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_589),
.A2(n_495),
.B1(n_481),
.B2(n_489),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_541),
.B(n_508),
.Y(n_772)
);

OR2x6_ASAP7_75t_L g773 ( 
.A(n_527),
.B(n_518),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_564),
.B(n_508),
.Y(n_774)
);

NAND2xp33_ASAP7_75t_L g775 ( 
.A(n_603),
.B(n_446),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_561),
.B(n_308),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_574),
.B(n_509),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_534),
.B(n_446),
.Y(n_778)
);

BUFx8_ASAP7_75t_L g779 ( 
.A(n_658),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_658),
.B(n_509),
.Y(n_780)
);

INVx8_ASAP7_75t_L g781 ( 
.A(n_574),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_604),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_574),
.B(n_618),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_636),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_652),
.B(n_509),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_527),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_L g787 ( 
.A(n_567),
.B(n_313),
.C(n_312),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_589),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_563),
.B(n_312),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_514),
.Y(n_790)
);

NOR3xp33_ASAP7_75t_L g791 ( 
.A(n_612),
.B(n_314),
.C(n_313),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_636),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_519),
.B(n_314),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_640),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_640),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_649),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_589),
.A2(n_481),
.B1(n_489),
.B2(n_495),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_610),
.B(n_475),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_649),
.Y(n_799)
);

NAND3xp33_ASAP7_75t_L g800 ( 
.A(n_659),
.B(n_328),
.C(n_321),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_525),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_518),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_661),
.B(n_475),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_SL g804 ( 
.A(n_535),
.B(n_634),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_634),
.A2(n_212),
.B1(n_215),
.B2(n_202),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_625),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_661),
.B(n_475),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_580),
.B(n_518),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_528),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_518),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_655),
.Y(n_811)
);

O2A1O1Ixp5_ASAP7_75t_L g812 ( 
.A1(n_556),
.A2(n_507),
.B(n_501),
.C(n_500),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_609),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_654),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_528),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_594),
.B(n_321),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_656),
.B(n_488),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_542),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_543),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_599),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_527),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_628),
.B(n_337),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_543),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_625),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_663),
.B(n_534),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_662),
.A2(n_533),
.B1(n_641),
.B2(n_625),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_705),
.B(n_656),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_724),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_682),
.A2(n_621),
.B(n_609),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_682),
.A2(n_623),
.B(n_621),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_701),
.A2(n_623),
.B(n_630),
.C(n_645),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_781),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_683),
.A2(n_645),
.B(n_630),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_R g834 ( 
.A(n_714),
.B(n_522),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_762),
.B(n_555),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_666),
.B(n_513),
.Y(n_836)
);

AOI21xp33_ASAP7_75t_L g837 ( 
.A1(n_822),
.A2(n_637),
.B(n_530),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_671),
.B(n_513),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_677),
.B(n_599),
.Y(n_839)
);

BUFx2_ASAP7_75t_SL g840 ( 
.A(n_663),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_813),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_726),
.B(n_500),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_699),
.B(n_559),
.Y(n_843)
);

AOI22x1_ASAP7_75t_L g844 ( 
.A1(n_693),
.A2(n_647),
.B1(n_530),
.B2(n_553),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_812),
.A2(n_647),
.B(n_536),
.Y(n_845)
);

NOR2xp67_ASAP7_75t_L g846 ( 
.A(n_674),
.B(n_546),
.Y(n_846)
);

NAND2x1_ASAP7_75t_L g847 ( 
.A(n_699),
.B(n_559),
.Y(n_847)
);

O2A1O1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_709),
.A2(n_579),
.B(n_536),
.C(n_538),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_699),
.B(n_559),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_735),
.B(n_531),
.Y(n_850)
);

NAND2x1_ASAP7_75t_L g851 ( 
.A(n_741),
.B(n_559),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_798),
.A2(n_700),
.B(n_703),
.C(n_664),
.Y(n_852)
);

NOR2x1_ASAP7_75t_L g853 ( 
.A(n_673),
.B(n_546),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_681),
.B(n_531),
.Y(n_854)
);

NOR2xp67_ASAP7_75t_L g855 ( 
.A(n_686),
.B(n_598),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_690),
.A2(n_540),
.B(n_538),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_781),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_695),
.B(n_556),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_683),
.A2(n_653),
.B(n_651),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_684),
.A2(n_653),
.B(n_651),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_820),
.B(n_540),
.Y(n_861)
);

NOR3xp33_ASAP7_75t_L g862 ( 
.A(n_667),
.B(n_598),
.C(n_298),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_697),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_707),
.Y(n_864)
);

OR2x6_ASAP7_75t_L g865 ( 
.A(n_773),
.B(n_570),
.Y(n_865)
);

AO21x1_ASAP7_75t_L g866 ( 
.A1(n_690),
.A2(n_551),
.B(n_545),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_684),
.A2(n_637),
.B(n_556),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_738),
.A2(n_648),
.B(n_553),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_685),
.B(n_500),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_739),
.B(n_570),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_813),
.Y(n_871)
);

O2A1O1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_692),
.A2(n_578),
.B(n_551),
.C(n_579),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_718),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_696),
.A2(n_578),
.B(n_581),
.C(n_582),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_675),
.B(n_581),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_744),
.A2(n_648),
.B(n_591),
.Y(n_876)
);

NAND2xp33_ASAP7_75t_L g877 ( 
.A(n_781),
.B(n_582),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_767),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_745),
.A2(n_648),
.B(n_592),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_698),
.A2(n_591),
.B(n_592),
.C(n_593),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_811),
.B(n_676),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_747),
.A2(n_593),
.B(n_552),
.Y(n_882)
);

AND2x2_ASAP7_75t_SL g883 ( 
.A(n_808),
.B(n_650),
.Y(n_883)
);

INVx4_ASAP7_75t_L g884 ( 
.A(n_781),
.Y(n_884)
);

O2A1O1Ixp5_ASAP7_75t_L g885 ( 
.A1(n_678),
.A2(n_575),
.B(n_549),
.C(n_552),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_780),
.B(n_549),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_747),
.A2(n_571),
.B(n_569),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_749),
.A2(n_571),
.B(n_569),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_710),
.B(n_712),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_767),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_749),
.A2(n_573),
.B(n_572),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_678),
.A2(n_573),
.B(n_572),
.C(n_595),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_729),
.A2(n_575),
.B1(n_595),
.B2(n_590),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_715),
.B(n_587),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_766),
.A2(n_588),
.B(n_587),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_716),
.B(n_737),
.Y(n_896)
);

AO21x2_ASAP7_75t_L g897 ( 
.A1(n_691),
.A2(n_590),
.B(n_588),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_766),
.A2(n_702),
.B(n_691),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_702),
.A2(n_568),
.B(n_542),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_774),
.B(n_570),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_668),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_783),
.A2(n_488),
.B(n_494),
.C(n_497),
.Y(n_902)
);

NOR3xp33_ASAP7_75t_L g903 ( 
.A(n_791),
.B(n_302),
.C(n_293),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_788),
.A2(n_633),
.B1(n_570),
.B2(n_605),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_741),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_732),
.A2(n_633),
.B(n_646),
.Y(n_906)
);

BUFx8_ASAP7_75t_L g907 ( 
.A(n_793),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_717),
.A2(n_568),
.B(n_542),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_785),
.B(n_633),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_732),
.A2(n_723),
.B(n_778),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_767),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_742),
.A2(n_633),
.B1(n_542),
.B2(n_605),
.Y(n_912)
);

OAI21xp33_ASAP7_75t_L g913 ( 
.A1(n_740),
.A2(n_752),
.B(n_816),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_SL g914 ( 
.A1(n_721),
.A2(n_247),
.B(n_252),
.C(n_269),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_788),
.A2(n_568),
.B1(n_605),
.B2(n_638),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_714),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_760),
.A2(n_494),
.B(n_497),
.C(n_500),
.Y(n_917)
);

BUFx8_ASAP7_75t_SL g918 ( 
.A(n_790),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_764),
.B(n_568),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_787),
.B(n_501),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_778),
.A2(n_522),
.B(n_493),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_721),
.A2(n_605),
.B(n_568),
.Y(n_922)
);

O2A1O1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_803),
.A2(n_507),
.B(n_501),
.C(n_493),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_768),
.B(n_605),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_728),
.A2(n_522),
.B(n_446),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_784),
.A2(n_343),
.B1(n_346),
.B2(n_337),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_728),
.A2(n_522),
.B(n_446),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_806),
.B(n_342),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_731),
.A2(n_522),
.B(n_446),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_792),
.A2(n_501),
.B(n_507),
.C(n_335),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_777),
.A2(n_522),
.B(n_493),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_794),
.B(n_507),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_789),
.B(n_342),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_790),
.Y(n_934)
);

O2A1O1Ixp33_ASAP7_75t_SL g935 ( 
.A1(n_731),
.A2(n_290),
.B(n_311),
.C(n_329),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_741),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_741),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_821),
.B(n_638),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_795),
.B(n_505),
.Y(n_939)
);

NAND2x1_ASAP7_75t_L g940 ( 
.A(n_748),
.B(n_642),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_750),
.Y(n_941)
);

NAND3xp33_ASAP7_75t_L g942 ( 
.A(n_763),
.B(n_343),
.C(n_344),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_669),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_786),
.B(n_638),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_754),
.A2(n_446),
.B(n_186),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_758),
.A2(n_446),
.B(n_186),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_796),
.A2(n_344),
.B(n_347),
.C(n_496),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_750),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_773),
.B(n_802),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_679),
.A2(n_493),
.B(n_642),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_750),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_799),
.B(n_505),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_769),
.A2(n_446),
.B(n_201),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_770),
.A2(n_772),
.B(n_733),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_669),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_814),
.B(n_505),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_773),
.B(n_505),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_670),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_725),
.A2(n_191),
.B(n_197),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_665),
.B(n_505),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_779),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_806),
.B(n_306),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_779),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_688),
.B(n_779),
.Y(n_964)
);

NOR3xp33_ASAP7_75t_L g965 ( 
.A(n_800),
.B(n_345),
.C(n_215),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_736),
.A2(n_200),
.B(n_212),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_750),
.Y(n_967)
);

AND2x6_ASAP7_75t_L g968 ( 
.A(n_810),
.B(n_338),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_824),
.B(n_505),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_805),
.B(n_200),
.Y(n_970)
);

AO21x1_ASAP7_75t_L g971 ( 
.A1(n_719),
.A2(n_282),
.B(n_203),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_807),
.A2(n_201),
.B(n_202),
.Y(n_972)
);

BUFx2_ASAP7_75t_SL g973 ( 
.A(n_727),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_824),
.B(n_505),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_776),
.B(n_481),
.Y(n_975)
);

BUFx4f_ASAP7_75t_L g976 ( 
.A(n_773),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_706),
.B(n_481),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_818),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_748),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_817),
.A2(n_307),
.B(n_309),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_734),
.A2(n_323),
.B(n_324),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_694),
.A2(n_481),
.B(n_489),
.C(n_495),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_748),
.B(n_481),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_782),
.A2(n_324),
.B(n_325),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_782),
.A2(n_489),
.B(n_495),
.C(n_496),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_704),
.B(n_489),
.Y(n_986)
);

AO21x1_ASAP7_75t_L g987 ( 
.A1(n_719),
.A2(n_203),
.B(n_282),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_782),
.A2(n_325),
.B(n_330),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_672),
.B(n_489),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_706),
.B(n_330),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_755),
.Y(n_991)
);

O2A1O1Ixp5_ASAP7_75t_L g992 ( 
.A1(n_730),
.A2(n_496),
.B(n_495),
.C(n_642),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_746),
.A2(n_331),
.B(n_339),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_823),
.B(n_819),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_823),
.B(n_496),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_711),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_746),
.A2(n_331),
.B(n_339),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_753),
.A2(n_345),
.B(n_273),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_818),
.Y(n_999)
);

AOI21x1_ASAP7_75t_L g1000 ( 
.A1(n_753),
.A2(n_642),
.B(n_496),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_757),
.B(n_642),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_708),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_757),
.B(n_642),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_761),
.A2(n_262),
.B(n_228),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_913),
.A2(n_804),
.B(n_711),
.C(n_708),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_909),
.A2(n_751),
.B(n_756),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_828),
.Y(n_1007)
);

OAI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_933),
.A2(n_759),
.B1(n_720),
.B2(n_815),
.Y(n_1008)
);

INVx4_ASAP7_75t_L g1009 ( 
.A(n_936),
.Y(n_1009)
);

NAND3xp33_ASAP7_75t_SL g1010 ( 
.A(n_862),
.B(n_287),
.C(n_225),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_954),
.A2(n_756),
.B(n_775),
.Y(n_1011)
);

INVx5_ASAP7_75t_L g1012 ( 
.A(n_865),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_827),
.B(n_765),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_862),
.A2(n_689),
.B(n_713),
.C(n_751),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_991),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_838),
.A2(n_775),
.B(n_689),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_852),
.A2(n_818),
.B(n_720),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_835),
.B(n_881),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_889),
.B(n_819),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_852),
.A2(n_818),
.B(n_809),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_839),
.B(n_765),
.Y(n_1021)
);

BUFx8_ASAP7_75t_L g1022 ( 
.A(n_890),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_949),
.B(n_801),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_869),
.B(n_680),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_963),
.B(n_687),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_970),
.B(n_687),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_863),
.Y(n_1027)
);

INVx2_ASAP7_75t_SL g1028 ( 
.A(n_934),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_864),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_961),
.B(n_722),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_875),
.A2(n_898),
.B(n_877),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_826),
.A2(n_771),
.B1(n_797),
.B2(n_743),
.Y(n_1032)
);

AO21x1_ASAP7_75t_L g1033 ( 
.A1(n_975),
.A2(n_282),
.B(n_203),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_854),
.A2(n_224),
.B1(n_232),
.B2(n_234),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_846),
.A2(n_642),
.B1(n_275),
.B2(n_300),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_842),
.B(n_11),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_1002),
.B(n_241),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_878),
.B(n_12),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_903),
.A2(n_13),
.B(n_16),
.C(n_17),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_918),
.Y(n_1040)
);

NOR2x1_ASAP7_75t_L g1041 ( 
.A(n_840),
.B(n_964),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_899),
.A2(n_271),
.B(n_299),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_908),
.A2(n_263),
.B(n_295),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_R g1044 ( 
.A(n_911),
.B(n_243),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_905),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_836),
.B(n_13),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_928),
.B(n_22),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_855),
.B(n_23),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_905),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_941),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_901),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_928),
.B(n_244),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_949),
.B(n_24),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_SL g1054 ( 
.A1(n_982),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_1054)
);

INVxp67_ASAP7_75t_L g1055 ( 
.A(n_986),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_962),
.B(n_873),
.Y(n_1056)
);

AOI21x1_ASAP7_75t_L g1057 ( 
.A1(n_971),
.A2(n_203),
.B(n_282),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_903),
.A2(n_29),
.B(n_32),
.C(n_34),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_975),
.A2(n_280),
.B(n_291),
.C(n_284),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_958),
.B(n_248),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_861),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_965),
.A2(n_958),
.B(n_947),
.C(n_896),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_962),
.B(n_253),
.Y(n_1063)
);

OAI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_886),
.A2(n_255),
.B1(n_338),
.B2(n_36),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_853),
.A2(n_338),
.B(n_282),
.C(n_203),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_907),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_850),
.A2(n_338),
.B1(n_35),
.B2(n_37),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_943),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_926),
.B(n_29),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_858),
.B(n_35),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_858),
.B(n_39),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_883),
.B(n_900),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_907),
.Y(n_1073)
);

NAND2x1p5_ASAP7_75t_L g1074 ( 
.A(n_976),
.B(n_338),
.Y(n_1074)
);

OAI21xp33_ASAP7_75t_SL g1075 ( 
.A1(n_870),
.A2(n_894),
.B(n_919),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_973),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_883),
.B(n_40),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_955),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_920),
.B(n_41),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_957),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_941),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_859),
.A2(n_282),
.B(n_203),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_916),
.B(n_41),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_916),
.B(n_42),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_936),
.B(n_44),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_996),
.B(n_44),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_937),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_996),
.B(n_45),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_941),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_932),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_874),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_874),
.A2(n_282),
.B(n_203),
.C(n_55),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_917),
.Y(n_1093)
);

AOI221xp5_ASAP7_75t_L g1094 ( 
.A1(n_965),
.A2(n_48),
.B1(n_54),
.B2(n_58),
.C(n_61),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_841),
.A2(n_282),
.B1(n_203),
.B2(n_63),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_832),
.B(n_58),
.Y(n_1096)
);

OAI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_937),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_860),
.A2(n_872),
.B(n_830),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_957),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_871),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_979),
.B(n_65),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_994),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_884),
.B(n_65),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_939),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_942),
.B(n_66),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_952),
.Y(n_1106)
);

OR2x6_ASAP7_75t_L g1107 ( 
.A(n_865),
.B(n_67),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_956),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_829),
.A2(n_73),
.B(n_74),
.Y(n_1109)
);

INVxp67_ASAP7_75t_L g1110 ( 
.A(n_990),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_832),
.B(n_77),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_976),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_833),
.A2(n_92),
.B(n_94),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_865),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_880),
.A2(n_95),
.B(n_101),
.C(n_111),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_880),
.A2(n_124),
.B1(n_131),
.B2(n_133),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_884),
.B(n_832),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_848),
.A2(n_148),
.B(n_150),
.C(n_156),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_948),
.B(n_166),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_848),
.A2(n_167),
.B1(n_171),
.B2(n_172),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_SL g1121 ( 
.A1(n_968),
.A2(n_173),
.B1(n_906),
.B2(n_832),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_995),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_857),
.B(n_910),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_857),
.B(n_837),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_948),
.B(n_951),
.Y(n_1125)
);

O2A1O1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_831),
.A2(n_930),
.B(n_892),
.C(n_902),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_941),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_967),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_951),
.B(n_999),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_999),
.B(n_944),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_984),
.B(n_988),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_868),
.A2(n_879),
.B(n_876),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_SL g1133 ( 
.A1(n_851),
.A2(n_940),
.B1(n_978),
.B2(n_967),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_867),
.A2(n_922),
.B(n_924),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_967),
.B(n_978),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_912),
.A2(n_895),
.B(n_888),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_982),
.A2(n_923),
.B(n_985),
.C(n_885),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_967),
.B(n_978),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_978),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_844),
.A2(n_893),
.B1(n_989),
.B2(n_856),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_SL g1141 ( 
.A1(n_845),
.A2(n_953),
.B(n_946),
.C(n_945),
.Y(n_1141)
);

NOR3xp33_ASAP7_75t_SL g1142 ( 
.A(n_959),
.B(n_966),
.C(n_972),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_969),
.B(n_974),
.Y(n_1143)
);

OR2x6_ASAP7_75t_L g1144 ( 
.A(n_938),
.B(n_825),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_866),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_968),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_977),
.B(n_960),
.Y(n_1147)
);

CKINVDCx14_ASAP7_75t_R g1148 ( 
.A(n_968),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_968),
.Y(n_1149)
);

NOR2xp67_ASAP7_75t_SL g1150 ( 
.A(n_980),
.B(n_981),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_887),
.B(n_983),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_968),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_993),
.B(n_997),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_977),
.B(n_882),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_998),
.B(n_915),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_891),
.B(n_985),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1001),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_897),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_885),
.A2(n_923),
.B(n_843),
.Y(n_1159)
);

AO31x2_ASAP7_75t_L g1160 ( 
.A1(n_1033),
.A2(n_987),
.A3(n_1003),
.B(n_929),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1007),
.B(n_1004),
.Y(n_1161)
);

O2A1O1Ixp5_ASAP7_75t_SL g1162 ( 
.A1(n_1067),
.A2(n_950),
.B(n_921),
.C(n_931),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1047),
.A2(n_1070),
.B1(n_1071),
.B2(n_1056),
.Y(n_1163)
);

OA21x2_ASAP7_75t_L g1164 ( 
.A1(n_1132),
.A2(n_992),
.B(n_1000),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1015),
.B(n_897),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1011),
.A2(n_849),
.B(n_992),
.Y(n_1166)
);

AO32x2_ASAP7_75t_L g1167 ( 
.A1(n_1091),
.A2(n_914),
.A3(n_935),
.B1(n_925),
.B2(n_927),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1077),
.A2(n_904),
.B1(n_847),
.B2(n_834),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1137),
.A2(n_1075),
.B(n_1140),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1061),
.B(n_1018),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1021),
.B(n_1026),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1053),
.B(n_1025),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1158),
.A2(n_1145),
.A3(n_1140),
.B(n_1159),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_1032),
.A2(n_1134),
.A3(n_1020),
.B(n_1065),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1082),
.A2(n_1098),
.B(n_1136),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_1022),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1052),
.A2(n_1063),
.B1(n_1072),
.B2(n_1079),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1027),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1031),
.A2(n_1017),
.B(n_1016),
.Y(n_1179)
);

AO21x2_ASAP7_75t_L g1180 ( 
.A1(n_1124),
.A2(n_1057),
.B(n_1156),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_1045),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1006),
.A2(n_1147),
.B(n_1154),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1010),
.A2(n_1069),
.B1(n_1107),
.B2(n_1078),
.Y(n_1183)
);

INVxp67_ASAP7_75t_SL g1184 ( 
.A(n_1024),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_1022),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1049),
.B(n_1029),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1147),
.A2(n_1008),
.B(n_1013),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1126),
.A2(n_1109),
.B(n_1113),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1050),
.Y(n_1189)
);

NAND3xp33_ASAP7_75t_L g1190 ( 
.A(n_1094),
.B(n_1091),
.C(n_1092),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1068),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_SL g1192 ( 
.A1(n_1116),
.A2(n_1120),
.B(n_1013),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1039),
.A2(n_1058),
.B(n_1105),
.C(n_1067),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1116),
.A2(n_1131),
.A3(n_1120),
.B(n_1122),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1123),
.A2(n_1093),
.B(n_1155),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1037),
.B(n_1060),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1019),
.A2(n_1141),
.B(n_1014),
.Y(n_1197)
);

AO21x1_ASAP7_75t_L g1198 ( 
.A1(n_1064),
.A2(n_1062),
.B(n_1046),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1112),
.B(n_1053),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1028),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1080),
.B(n_1099),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1012),
.B(n_1114),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1076),
.B(n_1023),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1157),
.A2(n_1151),
.B(n_1135),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_1107),
.Y(n_1205)
);

OA21x2_ASAP7_75t_L g1206 ( 
.A1(n_1115),
.A2(n_1118),
.B(n_1143),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1090),
.B(n_1102),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1048),
.A2(n_1005),
.B(n_1059),
.C(n_1036),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1121),
.A2(n_1153),
.B(n_1110),
.C(n_1095),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1100),
.Y(n_1210)
);

BUFx12f_ASAP7_75t_L g1211 ( 
.A(n_1066),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1107),
.B(n_1038),
.Y(n_1212)
);

NAND3xp33_ASAP7_75t_SL g1213 ( 
.A(n_1044),
.B(n_1040),
.C(n_1073),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1086),
.A2(n_1088),
.B1(n_1103),
.B2(n_1104),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_SL g1215 ( 
.A(n_1149),
.B(n_1012),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_1041),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1103),
.A2(n_1142),
.B(n_1119),
.C(n_1083),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1050),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_1050),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1148),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1085),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1084),
.A2(n_1108),
.B(n_1106),
.C(n_1035),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1101),
.A2(n_1097),
.B1(n_1034),
.B2(n_1143),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1030),
.B(n_1009),
.Y(n_1224)
);

BUFx10_ASAP7_75t_L g1225 ( 
.A(n_1081),
.Y(n_1225)
);

AO32x2_ASAP7_75t_L g1226 ( 
.A1(n_1133),
.A2(n_1009),
.A3(n_1034),
.B1(n_1054),
.B2(n_1055),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1051),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1023),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1096),
.A2(n_1144),
.B1(n_1101),
.B2(n_1130),
.Y(n_1229)
);

BUFx10_ASAP7_75t_L g1230 ( 
.A(n_1081),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1012),
.Y(n_1231)
);

OR2x6_ASAP7_75t_L g1232 ( 
.A(n_1146),
.B(n_1144),
.Y(n_1232)
);

INVx5_ASAP7_75t_L g1233 ( 
.A(n_1146),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1138),
.A2(n_1129),
.B(n_1117),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_SL g1235 ( 
.A(n_1042),
.B(n_1043),
.C(n_1129),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1117),
.A2(n_1111),
.B(n_1074),
.Y(n_1236)
);

O2A1O1Ixp5_ASAP7_75t_SL g1237 ( 
.A1(n_1087),
.A2(n_1150),
.B(n_1125),
.C(n_1144),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1081),
.B(n_1128),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1089),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1012),
.A2(n_1074),
.B1(n_1146),
.B2(n_1152),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_SL g1241 ( 
.A(n_1089),
.B(n_1139),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1089),
.Y(n_1242)
);

AO32x2_ASAP7_75t_L g1243 ( 
.A1(n_1127),
.A2(n_1091),
.A3(n_1067),
.B1(n_1140),
.B2(n_1032),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1139),
.A2(n_1127),
.B(n_1128),
.Y(n_1244)
);

NAND3xp33_ASAP7_75t_L g1245 ( 
.A(n_1127),
.B(n_1128),
.C(n_1139),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1052),
.A2(n_933),
.B(n_913),
.C(n_662),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1017),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1047),
.A2(n_662),
.B1(n_826),
.B2(n_827),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1053),
.B(n_677),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1052),
.A2(n_933),
.B(n_913),
.C(n_662),
.Y(n_1250)
);

OAI22x1_ASAP7_75t_L g1251 ( 
.A1(n_1077),
.A2(n_558),
.B1(n_808),
.B2(n_550),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1040),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_1040),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1017),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1017),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1027),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1047),
.A2(n_662),
.B1(n_826),
.B2(n_827),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1017),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1017),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1077),
.A2(n_667),
.B1(n_787),
.B2(n_883),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1050),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1017),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1061),
.B(n_662),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1082),
.A2(n_1098),
.B(n_1136),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1017),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1077),
.A2(n_933),
.B1(n_913),
.B2(n_667),
.Y(n_1266)
);

NOR2x1_ASAP7_75t_R g1267 ( 
.A(n_1066),
.B(n_514),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1082),
.A2(n_1098),
.B(n_1136),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1017),
.Y(n_1269)
);

O2A1O1Ixp5_ASAP7_75t_L g1270 ( 
.A1(n_1063),
.A2(n_933),
.B(n_1052),
.C(n_671),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1027),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1061),
.B(n_662),
.Y(n_1272)
);

INVx5_ASAP7_75t_L g1273 ( 
.A(n_1107),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1137),
.A2(n_1075),
.B(n_885),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1056),
.B(n_671),
.Y(n_1275)
);

BUFx8_ASAP7_75t_L g1276 ( 
.A(n_1028),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_1007),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1082),
.A2(n_1098),
.B(n_1136),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1082),
.A2(n_1098),
.B(n_1136),
.Y(n_1279)
);

CKINVDCx16_ASAP7_75t_R g1280 ( 
.A(n_1040),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1027),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1022),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1077),
.A2(n_667),
.B1(n_787),
.B2(n_883),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1040),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1017),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1015),
.Y(n_1286)
);

BUFx8_ASAP7_75t_L g1287 ( 
.A(n_1028),
.Y(n_1287)
);

BUFx2_ASAP7_75t_SL g1288 ( 
.A(n_1040),
.Y(n_1288)
);

AO22x1_ASAP7_75t_L g1289 ( 
.A1(n_1063),
.A2(n_767),
.B1(n_907),
.B2(n_787),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1027),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1047),
.A2(n_662),
.B1(n_826),
.B2(n_827),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1061),
.B(n_662),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1082),
.A2(n_1098),
.B(n_1136),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1015),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1015),
.Y(n_1295)
);

OR2x2_ASAP7_75t_L g1296 ( 
.A(n_1007),
.B(n_677),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1077),
.A2(n_667),
.B1(n_787),
.B2(n_883),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1022),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1027),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1007),
.B(n_677),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1082),
.A2(n_1098),
.B(n_1136),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1017),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1027),
.Y(n_1303)
);

INVx3_ASAP7_75t_SL g1304 ( 
.A(n_1066),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1017),
.Y(n_1305)
);

NAND2x1p5_ASAP7_75t_L g1306 ( 
.A(n_1012),
.B(n_976),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1052),
.A2(n_933),
.B(n_913),
.C(n_662),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1017),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1082),
.A2(n_1098),
.B(n_1136),
.Y(n_1309)
);

NAND3x1_ASAP7_75t_L g1310 ( 
.A(n_1041),
.B(n_787),
.C(n_808),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1017),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1082),
.A2(n_1098),
.B(n_1136),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1137),
.A2(n_1075),
.B(n_885),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1015),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1011),
.A2(n_1031),
.B(n_1017),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1061),
.B(n_662),
.Y(n_1316)
);

AO31x2_ASAP7_75t_L g1317 ( 
.A1(n_1033),
.A2(n_1158),
.A3(n_1145),
.B(n_866),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1251),
.A2(n_1260),
.B1(n_1297),
.B2(n_1283),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1184),
.B(n_1187),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1190),
.A2(n_1273),
.B1(n_1196),
.B2(n_1163),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1178),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1190),
.A2(n_1266),
.B1(n_1177),
.B2(n_1163),
.Y(n_1322)
);

BUFx4f_ASAP7_75t_SL g1323 ( 
.A(n_1211),
.Y(n_1323)
);

NAND2x1p5_ASAP7_75t_L g1324 ( 
.A(n_1273),
.B(n_1233),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1266),
.A2(n_1307),
.B1(n_1250),
.B2(n_1246),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1189),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1273),
.A2(n_1205),
.B1(n_1223),
.B2(n_1214),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1181),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1252),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1198),
.A2(n_1249),
.B1(n_1291),
.B2(n_1257),
.Y(n_1330)
);

CKINVDCx11_ASAP7_75t_R g1331 ( 
.A(n_1304),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1248),
.A2(n_1257),
.B1(n_1291),
.B2(n_1214),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1248),
.A2(n_1223),
.B1(n_1183),
.B2(n_1171),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1225),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1275),
.A2(n_1228),
.B1(n_1227),
.B2(n_1172),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1256),
.Y(n_1336)
);

INVx6_ASAP7_75t_L g1337 ( 
.A(n_1276),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1192),
.A2(n_1169),
.B1(n_1263),
.B2(n_1272),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1165),
.A2(n_1316),
.B1(n_1292),
.B2(n_1212),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1296),
.A2(n_1300),
.B1(n_1210),
.B2(n_1191),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1271),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1169),
.A2(n_1193),
.B1(n_1229),
.B2(n_1217),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1201),
.A2(n_1161),
.B1(n_1207),
.B2(n_1221),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1207),
.A2(n_1229),
.B1(n_1170),
.B2(n_1206),
.Y(n_1344)
);

CKINVDCx11_ASAP7_75t_R g1345 ( 
.A(n_1280),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1310),
.A2(n_1224),
.B1(n_1289),
.B2(n_1213),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1206),
.A2(n_1281),
.B1(n_1303),
.B2(n_1299),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1290),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1232),
.A2(n_1277),
.B1(n_1181),
.B2(n_1294),
.Y(n_1349)
);

BUFx8_ASAP7_75t_L g1350 ( 
.A(n_1185),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1186),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1239),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1204),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1209),
.A2(n_1277),
.B1(n_1274),
.B2(n_1313),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1232),
.A2(n_1286),
.B1(n_1314),
.B2(n_1295),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1242),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1199),
.A2(n_1202),
.B1(n_1203),
.B2(n_1240),
.Y(n_1357)
);

BUFx4f_ASAP7_75t_SL g1358 ( 
.A(n_1176),
.Y(n_1358)
);

INVx1_ASAP7_75t_SL g1359 ( 
.A(n_1218),
.Y(n_1359)
);

INVx3_ASAP7_75t_SL g1360 ( 
.A(n_1253),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1225),
.Y(n_1361)
);

CKINVDCx11_ASAP7_75t_R g1362 ( 
.A(n_1282),
.Y(n_1362)
);

INVx4_ASAP7_75t_L g1363 ( 
.A(n_1189),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1276),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_SL g1365 ( 
.A1(n_1215),
.A2(n_1270),
.B1(n_1274),
.B2(n_1313),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1240),
.A2(n_1235),
.B1(n_1220),
.B2(n_1215),
.Y(n_1366)
);

NAND2x1p5_ASAP7_75t_L g1367 ( 
.A(n_1233),
.B(n_1231),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1195),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1245),
.Y(n_1369)
);

OAI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1298),
.A2(n_1200),
.B1(n_1168),
.B2(n_1241),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1243),
.A2(n_1233),
.B1(n_1216),
.B2(n_1306),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1287),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1241),
.A2(n_1243),
.B1(n_1234),
.B2(n_1168),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1287),
.Y(n_1374)
);

OAI22x1_ASAP7_75t_L g1375 ( 
.A1(n_1243),
.A2(n_1245),
.B1(n_1284),
.B2(n_1267),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_1230),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1219),
.Y(n_1377)
);

CKINVDCx20_ASAP7_75t_R g1378 ( 
.A(n_1288),
.Y(n_1378)
);

INVx4_ASAP7_75t_L g1379 ( 
.A(n_1261),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1261),
.Y(n_1380)
);

BUFx10_ASAP7_75t_L g1381 ( 
.A(n_1238),
.Y(n_1381)
);

INVx4_ASAP7_75t_SL g1382 ( 
.A(n_1194),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1244),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1236),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1226),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1180),
.A2(n_1197),
.B1(n_1188),
.B2(n_1182),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_1267),
.Y(n_1387)
);

BUFx12f_ASAP7_75t_L g1388 ( 
.A(n_1237),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_1180),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1208),
.A2(n_1222),
.B(n_1258),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1247),
.A2(n_1265),
.B1(n_1302),
.B2(n_1269),
.Y(n_1391)
);

INVx4_ASAP7_75t_L g1392 ( 
.A(n_1164),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1254),
.A2(n_1285),
.B1(n_1305),
.B2(n_1308),
.Y(n_1393)
);

CKINVDCx11_ASAP7_75t_R g1394 ( 
.A(n_1226),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1166),
.A2(n_1194),
.B1(n_1164),
.B2(n_1179),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1255),
.A2(n_1262),
.B1(n_1311),
.B2(n_1315),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1259),
.A2(n_1162),
.B1(n_1226),
.B2(n_1268),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1173),
.B(n_1317),
.Y(n_1398)
);

OAI21xp33_ASAP7_75t_L g1399 ( 
.A1(n_1175),
.A2(n_1279),
.B(n_1309),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1264),
.A2(n_1293),
.B1(n_1312),
.B2(n_1278),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1317),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1167),
.A2(n_1174),
.B1(n_1317),
.B2(n_1160),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1167),
.A2(n_1174),
.B1(n_1160),
.B2(n_1301),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1167),
.A2(n_1266),
.B1(n_1190),
.B2(n_1260),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1174),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1251),
.A2(n_667),
.B1(n_787),
.B2(n_883),
.Y(n_1406)
);

CKINVDCx11_ASAP7_75t_R g1407 ( 
.A(n_1304),
.Y(n_1407)
);

INVx6_ASAP7_75t_L g1408 ( 
.A(n_1276),
.Y(n_1408)
);

OAI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1266),
.A2(n_1196),
.B1(n_1107),
.B2(n_558),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1266),
.A2(n_667),
.B1(n_933),
.B2(n_913),
.Y(n_1410)
);

BUFx8_ASAP7_75t_SL g1411 ( 
.A(n_1252),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1178),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1266),
.A2(n_667),
.B1(n_933),
.B2(n_913),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1178),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1184),
.B(n_1187),
.Y(n_1415)
);

CKINVDCx11_ASAP7_75t_R g1416 ( 
.A(n_1304),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1252),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1178),
.Y(n_1418)
);

BUFx12f_ASAP7_75t_L g1419 ( 
.A(n_1252),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1280),
.Y(n_1420)
);

CKINVDCx8_ASAP7_75t_R g1421 ( 
.A(n_1288),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1178),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1266),
.A2(n_1196),
.B1(n_1107),
.B2(n_558),
.Y(n_1423)
);

INVx6_ASAP7_75t_L g1424 ( 
.A(n_1276),
.Y(n_1424)
);

BUFx12f_ASAP7_75t_L g1425 ( 
.A(n_1252),
.Y(n_1425)
);

CKINVDCx6p67_ASAP7_75t_R g1426 ( 
.A(n_1304),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1178),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1266),
.A2(n_1190),
.B1(n_1283),
.B2(n_1260),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1190),
.A2(n_667),
.B1(n_808),
.B2(n_375),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1251),
.A2(n_667),
.B1(n_787),
.B2(n_883),
.Y(n_1430)
);

INVx11_ASAP7_75t_L g1431 ( 
.A(n_1276),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1266),
.A2(n_1190),
.B1(n_1283),
.B2(n_1260),
.Y(n_1432)
);

NAND2x1p5_ASAP7_75t_L g1433 ( 
.A(n_1273),
.B(n_1012),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1266),
.A2(n_1190),
.B1(n_1283),
.B2(n_1260),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1266),
.A2(n_1190),
.B1(n_1283),
.B2(n_1260),
.Y(n_1435)
);

INVxp67_ASAP7_75t_SL g1436 ( 
.A(n_1184),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1251),
.A2(n_667),
.B1(n_787),
.B2(n_883),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1251),
.A2(n_667),
.B1(n_787),
.B2(n_883),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1266),
.A2(n_1190),
.B1(n_1283),
.B2(n_1260),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1266),
.A2(n_1190),
.B1(n_1283),
.B2(n_1260),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1178),
.Y(n_1441)
);

BUFx10_ASAP7_75t_L g1442 ( 
.A(n_1252),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1181),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1178),
.Y(n_1444)
);

INVx6_ASAP7_75t_L g1445 ( 
.A(n_1276),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1178),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_SL g1447 ( 
.A(n_1428),
.B(n_1432),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1368),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1319),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1436),
.B(n_1332),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1319),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1415),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_1392),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1397),
.A2(n_1396),
.B(n_1386),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1385),
.B(n_1321),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1415),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1351),
.B(n_1328),
.Y(n_1457)
);

NOR2xp67_ASAP7_75t_L g1458 ( 
.A(n_1390),
.B(n_1375),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1410),
.A2(n_1413),
.B(n_1325),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1336),
.B(n_1341),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1353),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1328),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1443),
.B(n_1338),
.Y(n_1463)
);

BUFx4f_ASAP7_75t_SL g1464 ( 
.A(n_1419),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1398),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1398),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1412),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1446),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1443),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1414),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1418),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1382),
.B(n_1384),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1422),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1394),
.A2(n_1429),
.B1(n_1438),
.B2(n_1430),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1427),
.B(n_1441),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1444),
.B(n_1348),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1405),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1391),
.A2(n_1393),
.B(n_1400),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_SL g1479 ( 
.A1(n_1428),
.A2(n_1439),
.B1(n_1434),
.B2(n_1432),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1338),
.B(n_1354),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1391),
.A2(n_1393),
.B(n_1395),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1401),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1399),
.A2(n_1403),
.B(n_1402),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1354),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1359),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1403),
.A2(n_1402),
.B(n_1342),
.Y(n_1486)
);

INVx2_ASAP7_75t_SL g1487 ( 
.A(n_1381),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1343),
.B(n_1404),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1404),
.B(n_1339),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1347),
.B(n_1365),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1369),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1352),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1388),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1330),
.B(n_1322),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1359),
.Y(n_1495)
);

AOI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1325),
.A2(n_1342),
.B(n_1439),
.Y(n_1496)
);

INVxp67_ASAP7_75t_SL g1497 ( 
.A(n_1344),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1389),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1381),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1326),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1373),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1356),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1383),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_SL g1504 ( 
.A1(n_1434),
.A2(n_1435),
.B1(n_1440),
.B2(n_1409),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1333),
.B(n_1320),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1435),
.A2(n_1440),
.B(n_1423),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1377),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1371),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1380),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1370),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1327),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1340),
.B(n_1349),
.Y(n_1512)
);

AO21x2_ASAP7_75t_L g1513 ( 
.A1(n_1346),
.A2(n_1318),
.B(n_1366),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1367),
.A2(n_1324),
.B(n_1433),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1367),
.A2(n_1324),
.B(n_1433),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1335),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1363),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1406),
.A2(n_1437),
.B(n_1357),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1420),
.A2(n_1387),
.B1(n_1355),
.B2(n_1378),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1379),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1411),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1334),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1361),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1376),
.B(n_1374),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1364),
.B(n_1372),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1337),
.B(n_1408),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1421),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1350),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1337),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1472),
.B(n_1417),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1486),
.B(n_1445),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1462),
.B(n_1445),
.Y(n_1532)
);

AOI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1447),
.A2(n_1479),
.B1(n_1504),
.B2(n_1506),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1467),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1447),
.B(n_1424),
.Y(n_1535)
);

NAND2x1_ASAP7_75t_L g1536 ( 
.A(n_1500),
.B(n_1408),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1457),
.B(n_1469),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1485),
.B(n_1424),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1467),
.Y(n_1539)
);

OA21x2_ASAP7_75t_L g1540 ( 
.A1(n_1478),
.A2(n_1329),
.B(n_1408),
.Y(n_1540)
);

OA21x2_ASAP7_75t_L g1541 ( 
.A1(n_1478),
.A2(n_1424),
.B(n_1337),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1459),
.A2(n_1426),
.B1(n_1431),
.B2(n_1358),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1459),
.A2(n_1360),
.B1(n_1323),
.B2(n_1425),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1495),
.B(n_1442),
.Y(n_1544)
);

NOR2x1_ASAP7_75t_R g1545 ( 
.A(n_1528),
.B(n_1345),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1457),
.B(n_1331),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1455),
.B(n_1407),
.Y(n_1547)
);

NAND2xp33_ASAP7_75t_L g1548 ( 
.A(n_1480),
.B(n_1506),
.Y(n_1548)
);

AOI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1458),
.A2(n_1416),
.B(n_1350),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1507),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1480),
.A2(n_1362),
.B1(n_1458),
.B2(n_1496),
.Y(n_1551)
);

NAND2xp33_ASAP7_75t_L g1552 ( 
.A(n_1484),
.B(n_1450),
.Y(n_1552)
);

AOI221xp5_ASAP7_75t_L g1553 ( 
.A1(n_1494),
.A2(n_1505),
.B1(n_1501),
.B2(n_1488),
.C(n_1490),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1455),
.B(n_1460),
.Y(n_1554)
);

A2O1A1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1505),
.A2(n_1494),
.B(n_1490),
.C(n_1488),
.Y(n_1555)
);

A2O1A1Ixp33_ASAP7_75t_L g1556 ( 
.A1(n_1474),
.A2(n_1489),
.B(n_1511),
.C(n_1463),
.Y(n_1556)
);

A2O1A1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1489),
.A2(n_1511),
.B(n_1450),
.C(n_1497),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1496),
.B(n_1487),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1509),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1518),
.A2(n_1491),
.B(n_1493),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1460),
.B(n_1475),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1487),
.B(n_1499),
.Y(n_1562)
);

OAI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1481),
.A2(n_1515),
.B(n_1514),
.Y(n_1563)
);

A2O1A1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1501),
.A2(n_1510),
.B(n_1508),
.C(n_1512),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1475),
.B(n_1468),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1499),
.B(n_1493),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1470),
.B(n_1471),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1518),
.A2(n_1491),
.B(n_1493),
.Y(n_1568)
);

AO21x1_ASAP7_75t_L g1569 ( 
.A1(n_1492),
.A2(n_1449),
.B(n_1451),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1449),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1473),
.B(n_1451),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1498),
.B(n_1476),
.Y(n_1572)
);

OA21x2_ASAP7_75t_L g1573 ( 
.A1(n_1481),
.A2(n_1456),
.B(n_1452),
.Y(n_1573)
);

OAI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1518),
.A2(n_1493),
.B(n_1503),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1498),
.B(n_1476),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1452),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1456),
.A2(n_1454),
.B(n_1513),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1503),
.A2(n_1453),
.B(n_1482),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1492),
.Y(n_1579)
);

O2A1O1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1513),
.A2(n_1510),
.B(n_1529),
.C(n_1527),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1522),
.A2(n_1523),
.B(n_1454),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1513),
.A2(n_1516),
.B1(n_1512),
.B2(n_1466),
.C(n_1465),
.Y(n_1582)
);

AOI221xp5_ASAP7_75t_L g1583 ( 
.A1(n_1513),
.A2(n_1516),
.B1(n_1465),
.B2(n_1466),
.C(n_1519),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1522),
.Y(n_1584)
);

OAI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1523),
.A2(n_1454),
.B(n_1520),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1536),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1561),
.B(n_1483),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1537),
.B(n_1483),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1570),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1554),
.B(n_1483),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1576),
.B(n_1571),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1554),
.B(n_1483),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1565),
.B(n_1453),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1534),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1571),
.B(n_1558),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1539),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1581),
.B(n_1573),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1533),
.A2(n_1454),
.B1(n_1502),
.B2(n_1477),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1578),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1548),
.A2(n_1555),
.B1(n_1553),
.B2(n_1556),
.Y(n_1600)
);

INVxp67_ASAP7_75t_SL g1601 ( 
.A(n_1569),
.Y(n_1601)
);

INVxp67_ASAP7_75t_SL g1602 ( 
.A(n_1578),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1531),
.Y(n_1603)
);

BUFx2_ASAP7_75t_L g1604 ( 
.A(n_1531),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1548),
.B(n_1524),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1558),
.B(n_1524),
.Y(n_1606)
);

NOR2x1_ASAP7_75t_SL g1607 ( 
.A(n_1550),
.B(n_1526),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1573),
.B(n_1448),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1579),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1573),
.B(n_1567),
.Y(n_1610)
);

NOR2x1p5_ASAP7_75t_L g1611 ( 
.A(n_1549),
.B(n_1517),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1559),
.B(n_1448),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1585),
.B(n_1461),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1584),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1594),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1612),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1588),
.B(n_1560),
.Y(n_1617)
);

INVxp67_ASAP7_75t_SL g1618 ( 
.A(n_1601),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1610),
.B(n_1587),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1608),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1600),
.A2(n_1555),
.B1(n_1556),
.B2(n_1583),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1588),
.B(n_1568),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1610),
.Y(n_1623)
);

INVx5_ASAP7_75t_L g1624 ( 
.A(n_1597),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1590),
.B(n_1578),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1590),
.B(n_1592),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1610),
.B(n_1552),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1586),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1594),
.Y(n_1629)
);

CKINVDCx16_ASAP7_75t_R g1630 ( 
.A(n_1586),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1596),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1590),
.B(n_1540),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1588),
.B(n_1574),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1592),
.B(n_1540),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1592),
.B(n_1563),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1600),
.A2(n_1582),
.B1(n_1551),
.B2(n_1577),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1596),
.Y(n_1637)
);

NAND4xp25_ASAP7_75t_L g1638 ( 
.A(n_1605),
.B(n_1566),
.C(n_1562),
.D(n_1542),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1587),
.B(n_1540),
.Y(n_1639)
);

NAND3xp33_ASAP7_75t_SL g1640 ( 
.A(n_1598),
.B(n_1557),
.C(n_1535),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1587),
.B(n_1541),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1613),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1597),
.B(n_1541),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1593),
.B(n_1541),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1606),
.B(n_1546),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1593),
.B(n_1572),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1593),
.B(n_1575),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1599),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1613),
.Y(n_1649)
);

NOR2x1_ASAP7_75t_L g1650 ( 
.A(n_1586),
.B(n_1530),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1609),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1620),
.Y(n_1652)
);

INVx4_ASAP7_75t_L g1653 ( 
.A(n_1624),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1624),
.B(n_1607),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1618),
.B(n_1589),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1624),
.B(n_1607),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1615),
.Y(n_1657)
);

NOR2x1p5_ASAP7_75t_L g1658 ( 
.A(n_1618),
.B(n_1601),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1624),
.B(n_1595),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1624),
.B(n_1603),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1624),
.B(n_1603),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1615),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_R g1663 ( 
.A(n_1628),
.B(n_1521),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_R g1664 ( 
.A(n_1630),
.B(n_1464),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1624),
.B(n_1604),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1621),
.A2(n_1557),
.B(n_1564),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1642),
.B(n_1589),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1642),
.B(n_1597),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1626),
.B(n_1604),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1645),
.B(n_1638),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1629),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1629),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1631),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1649),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1649),
.B(n_1614),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1619),
.B(n_1591),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1644),
.B(n_1623),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1651),
.B(n_1631),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1637),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1648),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1637),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1623),
.B(n_1606),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1620),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1623),
.B(n_1635),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1657),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1657),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1669),
.B(n_1630),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1669),
.B(n_1650),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1666),
.A2(n_1640),
.B1(n_1621),
.B2(n_1636),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1657),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1662),
.Y(n_1691)
);

INVxp67_ASAP7_75t_SL g1692 ( 
.A(n_1658),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1676),
.B(n_1619),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1670),
.B(n_1617),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1666),
.A2(n_1636),
.B(n_1640),
.Y(n_1695)
);

NAND2x1p5_ASAP7_75t_L g1696 ( 
.A(n_1653),
.B(n_1650),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1662),
.Y(n_1697)
);

OAI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1668),
.A2(n_1633),
.B1(n_1617),
.B2(n_1622),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1662),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1676),
.B(n_1617),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1669),
.B(n_1656),
.Y(n_1701)
);

NAND4xp25_ASAP7_75t_L g1702 ( 
.A(n_1670),
.B(n_1562),
.C(n_1638),
.D(n_1566),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1663),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1671),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1658),
.A2(n_1627),
.B1(n_1605),
.B2(n_1622),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1676),
.B(n_1622),
.Y(n_1706)
);

INVxp33_ASAP7_75t_SL g1707 ( 
.A(n_1664),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1667),
.B(n_1627),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1674),
.B(n_1633),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1671),
.Y(n_1710)
);

INVxp67_ASAP7_75t_SL g1711 ( 
.A(n_1658),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1674),
.B(n_1633),
.Y(n_1712)
);

NOR2x1_ASAP7_75t_L g1713 ( 
.A(n_1653),
.B(n_1528),
.Y(n_1713)
);

NOR2xp67_ASAP7_75t_R g1714 ( 
.A(n_1653),
.B(n_1674),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1671),
.Y(n_1715)
);

NAND2x1p5_ASAP7_75t_L g1716 ( 
.A(n_1653),
.B(n_1611),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1672),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1655),
.B(n_1625),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1652),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1656),
.B(n_1646),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1652),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1652),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1656),
.B(n_1646),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1654),
.B(n_1646),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1654),
.B(n_1647),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1667),
.B(n_1616),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1654),
.B(n_1647),
.Y(n_1727)
);

OR2x6_ASAP7_75t_L g1728 ( 
.A(n_1695),
.B(n_1653),
.Y(n_1728)
);

NOR4xp25_ASAP7_75t_L g1729 ( 
.A(n_1689),
.B(n_1655),
.C(n_1668),
.D(n_1648),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1687),
.B(n_1654),
.Y(n_1730)
);

AND3x2_ASAP7_75t_L g1731 ( 
.A(n_1692),
.B(n_1535),
.C(n_1547),
.Y(n_1731)
);

NAND3xp33_ASAP7_75t_L g1732 ( 
.A(n_1694),
.B(n_1653),
.C(n_1680),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1700),
.B(n_1682),
.Y(n_1733)
);

OR2x6_ASAP7_75t_L g1734 ( 
.A(n_1713),
.B(n_1716),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1697),
.Y(n_1735)
);

INVxp33_ASAP7_75t_L g1736 ( 
.A(n_1687),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1700),
.B(n_1682),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1719),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1685),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1703),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1706),
.B(n_1675),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1705),
.A2(n_1598),
.B1(n_1711),
.B2(n_1639),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1685),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1707),
.B(n_1545),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1706),
.B(n_1682),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1698),
.B(n_1673),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1719),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1709),
.B(n_1673),
.Y(n_1748)
);

INVxp33_ASAP7_75t_L g1749 ( 
.A(n_1714),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1686),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1721),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1710),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1686),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1712),
.B(n_1679),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1690),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1690),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1721),
.Y(n_1757)
);

OAI21xp33_ASAP7_75t_L g1758 ( 
.A1(n_1702),
.A2(n_1684),
.B(n_1659),
.Y(n_1758)
);

OAI31xp33_ASAP7_75t_L g1759 ( 
.A1(n_1718),
.A2(n_1643),
.A3(n_1639),
.B(n_1634),
.Y(n_1759)
);

OR2x6_ASAP7_75t_L g1760 ( 
.A(n_1716),
.B(n_1580),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1717),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1691),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1693),
.B(n_1679),
.Y(n_1763)
);

INVxp67_ASAP7_75t_L g1764 ( 
.A(n_1691),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1728),
.B(n_1688),
.Y(n_1765)
);

OAI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1729),
.A2(n_1707),
.B(n_1688),
.Y(n_1766)
);

OAI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1760),
.A2(n_1643),
.B1(n_1602),
.B2(n_1693),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1742),
.A2(n_1696),
.B1(n_1660),
.B2(n_1661),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1735),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1733),
.B(n_1708),
.Y(n_1770)
);

INVx1_ASAP7_75t_SL g1771 ( 
.A(n_1740),
.Y(n_1771)
);

OAI22xp5_ASAP7_75t_L g1772 ( 
.A1(n_1736),
.A2(n_1696),
.B1(n_1660),
.B2(n_1661),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1728),
.B(n_1701),
.Y(n_1773)
);

INVx1_ASAP7_75t_SL g1774 ( 
.A(n_1740),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1728),
.B(n_1701),
.Y(n_1775)
);

OAI332xp33_ASAP7_75t_L g1776 ( 
.A1(n_1746),
.A2(n_1708),
.A3(n_1726),
.B1(n_1648),
.B2(n_1722),
.B3(n_1704),
.C1(n_1699),
.C2(n_1715),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1760),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1752),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1761),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1744),
.B(n_1645),
.Y(n_1780)
);

A2O1A1Ixp33_ASAP7_75t_L g1781 ( 
.A1(n_1759),
.A2(n_1602),
.B(n_1564),
.C(n_1625),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1760),
.Y(n_1782)
);

OAI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1760),
.A2(n_1599),
.B1(n_1639),
.B2(n_1632),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1728),
.Y(n_1784)
);

AOI21xp33_ASAP7_75t_L g1785 ( 
.A1(n_1749),
.A2(n_1704),
.B(n_1699),
.Y(n_1785)
);

A2O1A1Ixp33_ASAP7_75t_L g1786 ( 
.A1(n_1758),
.A2(n_1625),
.B(n_1634),
.C(n_1632),
.Y(n_1786)
);

XNOR2x1_ASAP7_75t_L g1787 ( 
.A(n_1731),
.B(n_1543),
.Y(n_1787)
);

AOI32xp33_ASAP7_75t_L g1788 ( 
.A1(n_1737),
.A2(n_1677),
.A3(n_1632),
.B1(n_1634),
.B2(n_1684),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1739),
.Y(n_1789)
);

INVx1_ASAP7_75t_SL g1790 ( 
.A(n_1748),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1771),
.B(n_1730),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1789),
.Y(n_1792)
);

OAI21xp33_ASAP7_75t_L g1793 ( 
.A1(n_1766),
.A2(n_1745),
.B(n_1754),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_1774),
.B(n_1664),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1790),
.B(n_1763),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1770),
.B(n_1741),
.Y(n_1796)
);

AOI221xp5_ASAP7_75t_L g1797 ( 
.A1(n_1776),
.A2(n_1764),
.B1(n_1732),
.B2(n_1762),
.C(n_1756),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1773),
.B(n_1730),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1770),
.B(n_1741),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1773),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1769),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1777),
.A2(n_1738),
.B1(n_1751),
.B2(n_1757),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1778),
.B(n_1739),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1777),
.A2(n_1738),
.B1(n_1747),
.B2(n_1757),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1779),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1784),
.B(n_1743),
.Y(n_1806)
);

AOI211xp5_ASAP7_75t_L g1807 ( 
.A1(n_1767),
.A2(n_1762),
.B(n_1756),
.C(n_1755),
.Y(n_1807)
);

A2O1A1Ixp33_ASAP7_75t_L g1808 ( 
.A1(n_1781),
.A2(n_1751),
.B(n_1747),
.C(n_1635),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1787),
.A2(n_1641),
.B1(n_1734),
.B2(n_1635),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1782),
.Y(n_1810)
);

OAI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1782),
.A2(n_1734),
.B1(n_1755),
.B2(n_1753),
.Y(n_1811)
);

OAI21xp33_ASAP7_75t_L g1812 ( 
.A1(n_1793),
.A2(n_1781),
.B(n_1775),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1796),
.Y(n_1813)
);

INVxp67_ASAP7_75t_L g1814 ( 
.A(n_1794),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1799),
.B(n_1726),
.Y(n_1815)
);

AOI222xp33_ASAP7_75t_L g1816 ( 
.A1(n_1797),
.A2(n_1804),
.B1(n_1802),
.B2(n_1810),
.C1(n_1808),
.C2(n_1795),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1794),
.B(n_1780),
.Y(n_1817)
);

XOR2xp5_ASAP7_75t_L g1818 ( 
.A(n_1791),
.B(n_1787),
.Y(n_1818)
);

OAI21xp5_ASAP7_75t_SL g1819 ( 
.A1(n_1809),
.A2(n_1765),
.B(n_1775),
.Y(n_1819)
);

OA21x2_ASAP7_75t_L g1820 ( 
.A1(n_1802),
.A2(n_1785),
.B(n_1786),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1800),
.A2(n_1786),
.B1(n_1734),
.B2(n_1768),
.Y(n_1821)
);

OAI211xp5_ASAP7_75t_L g1822 ( 
.A1(n_1807),
.A2(n_1765),
.B(n_1788),
.C(n_1772),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1818),
.B(n_1798),
.Y(n_1823)
);

NOR2x1_ASAP7_75t_L g1824 ( 
.A(n_1817),
.B(n_1811),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1815),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1813),
.B(n_1801),
.Y(n_1826)
);

OAI21xp33_ASAP7_75t_L g1827 ( 
.A1(n_1816),
.A2(n_1805),
.B(n_1803),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1814),
.Y(n_1828)
);

BUFx2_ASAP7_75t_L g1829 ( 
.A(n_1820),
.Y(n_1829)
);

NAND3xp33_ASAP7_75t_L g1830 ( 
.A(n_1820),
.B(n_1804),
.C(n_1806),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1812),
.B(n_1811),
.Y(n_1831)
);

NAND3xp33_ASAP7_75t_L g1832 ( 
.A(n_1830),
.B(n_1819),
.C(n_1822),
.Y(n_1832)
);

AOI221xp5_ASAP7_75t_L g1833 ( 
.A1(n_1829),
.A2(n_1827),
.B1(n_1831),
.B2(n_1821),
.C(n_1783),
.Y(n_1833)
);

NAND3xp33_ASAP7_75t_L g1834 ( 
.A(n_1824),
.B(n_1792),
.C(n_1734),
.Y(n_1834)
);

AOI211xp5_ASAP7_75t_SL g1835 ( 
.A1(n_1827),
.A2(n_1753),
.B(n_1750),
.C(n_1743),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1828),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1835),
.B(n_1825),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1832),
.A2(n_1823),
.B1(n_1826),
.B2(n_1750),
.Y(n_1838)
);

O2A1O1Ixp33_ASAP7_75t_L g1839 ( 
.A1(n_1833),
.A2(n_1680),
.B(n_1722),
.C(n_1648),
.Y(n_1839)
);

OAI211xp5_ASAP7_75t_L g1840 ( 
.A1(n_1836),
.A2(n_1834),
.B(n_1663),
.C(n_1715),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_SL g1841 ( 
.A1(n_1832),
.A2(n_1716),
.B1(n_1696),
.B2(n_1547),
.Y(n_1841)
);

AOI211xp5_ASAP7_75t_L g1842 ( 
.A1(n_1832),
.A2(n_1525),
.B(n_1684),
.C(n_1677),
.Y(n_1842)
);

XNOR2xp5_ASAP7_75t_L g1843 ( 
.A(n_1838),
.B(n_1524),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1841),
.B(n_1720),
.Y(n_1844)
);

INVxp67_ASAP7_75t_SL g1845 ( 
.A(n_1837),
.Y(n_1845)
);

INVxp67_ASAP7_75t_SL g1846 ( 
.A(n_1839),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1840),
.B(n_1720),
.Y(n_1847)
);

NAND4xp75_ASAP7_75t_L g1848 ( 
.A(n_1844),
.B(n_1842),
.C(n_1665),
.D(n_1661),
.Y(n_1848)
);

AOI211xp5_ASAP7_75t_L g1849 ( 
.A1(n_1845),
.A2(n_1677),
.B(n_1524),
.C(n_1660),
.Y(n_1849)
);

OAI21xp33_ASAP7_75t_SL g1850 ( 
.A1(n_1845),
.A2(n_1727),
.B(n_1725),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1850),
.B(n_1847),
.Y(n_1851)
);

OAI22x1_ASAP7_75t_L g1852 ( 
.A1(n_1851),
.A2(n_1846),
.B1(n_1843),
.B2(n_1847),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1852),
.Y(n_1853)
);

OA21x2_ASAP7_75t_L g1854 ( 
.A1(n_1852),
.A2(n_1848),
.B(n_1849),
.Y(n_1854)
);

OAI22x1_ASAP7_75t_L g1855 ( 
.A1(n_1853),
.A2(n_1544),
.B1(n_1652),
.B2(n_1683),
.Y(n_1855)
);

INVxp67_ASAP7_75t_L g1856 ( 
.A(n_1854),
.Y(n_1856)
);

OAI21x1_ASAP7_75t_L g1857 ( 
.A1(n_1856),
.A2(n_1854),
.B(n_1723),
.Y(n_1857)
);

OAI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1855),
.A2(n_1683),
.B(n_1675),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1857),
.A2(n_1683),
.B(n_1678),
.Y(n_1859)
);

OAI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1859),
.A2(n_1858),
.B(n_1683),
.Y(n_1860)
);

AOI22x1_ASAP7_75t_L g1861 ( 
.A1(n_1860),
.A2(n_1727),
.B1(n_1725),
.B2(n_1724),
.Y(n_1861)
);

AOI221xp5_ASAP7_75t_L g1862 ( 
.A1(n_1861),
.A2(n_1681),
.B1(n_1672),
.B2(n_1538),
.C(n_1659),
.Y(n_1862)
);

AOI211xp5_ASAP7_75t_L g1863 ( 
.A1(n_1862),
.A2(n_1532),
.B(n_1665),
.C(n_1723),
.Y(n_1863)
);


endmodule