module fake_jpeg_28861_n_102 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_6),
.B(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_10),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_21),
.B(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_18),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_1),
.B(n_4),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_20),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_33),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_27),
.Y(n_40)
);

INVxp33_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_47),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_26),
.C(n_28),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_41),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_36),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_49),
.Y(n_63)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_29),
.B1(n_24),
.B2(n_18),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_35),
.B1(n_23),
.B2(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_34),
.B1(n_36),
.B2(n_35),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_64),
.B1(n_39),
.B2(n_40),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_62),
.C(n_19),
.Y(n_74)
);

AO21x1_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_61),
.B(n_52),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_22),
.B1(n_14),
.B2(n_15),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_11),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_68),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_64),
.B1(n_39),
.B2(n_47),
.Y(n_80)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_72),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_42),
.B(n_40),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_74),
.C(n_19),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_R g71 ( 
.A(n_54),
.B(n_42),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_61),
.B(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_73),
.B(n_59),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_76),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_80),
.B(n_13),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_68),
.C(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_16),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_82),
.A2(n_14),
.B(n_15),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_84),
.C(n_85),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_71),
.B(n_69),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_70),
.C(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_78),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_77),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_91),
.B1(n_92),
.B2(n_67),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_75),
.Y(n_91)
);

OAI21x1_ASAP7_75t_SL g93 ( 
.A1(n_91),
.A2(n_90),
.B(n_81),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_12),
.B1(n_9),
.B2(n_5),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_67),
.A3(n_23),
.B1(n_12),
.B2(n_8),
.C1(n_7),
.C2(n_9),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_8),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_93),
.Y(n_97)
);

AOI322xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_1),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_52),
.C2(n_97),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_97),
.A2(n_98),
.B(n_4),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_101),
.Y(n_102)
);


endmodule