module fake_jpeg_191_n_577 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_577);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_577;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_54),
.B(n_62),
.Y(n_119)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_25),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_63),
.B(n_67),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_70),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_65),
.Y(n_140)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_31),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_68),
.B(n_79),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_21),
.B(n_9),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_91),
.Y(n_131)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_74),
.Y(n_164)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_85),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_86),
.B(n_90),
.Y(n_161)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_89),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_22),
.B(n_0),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_28),
.B(n_38),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_92),
.B(n_105),
.Y(n_169)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

BUFx10_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_98),
.Y(n_168)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_40),
.B(n_1),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_106),
.B(n_35),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_108),
.Y(n_136)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_61),
.A2(n_26),
.B1(n_27),
.B2(n_24),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_109),
.A2(n_110),
.B1(n_129),
.B2(n_130),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_75),
.A2(n_26),
.B1(n_27),
.B2(n_24),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_72),
.A2(n_23),
.B1(n_22),
.B2(n_53),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_122),
.A2(n_141),
.B1(n_146),
.B2(n_95),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_64),
.A2(n_38),
.B1(n_52),
.B2(n_51),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_26),
.B1(n_27),
.B2(n_24),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_89),
.A2(n_52),
.B1(n_51),
.B2(n_28),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_137),
.A2(n_142),
.B1(n_144),
.B2(n_147),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_91),
.A2(n_22),
.B1(n_53),
.B2(n_42),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_71),
.A2(n_26),
.B1(n_22),
.B2(n_34),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_60),
.A2(n_48),
.B1(n_43),
.B2(n_53),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_113),
.B(n_169),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_58),
.A2(n_50),
.B1(n_42),
.B2(n_33),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_55),
.A2(n_48),
.B1(n_43),
.B2(n_35),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_106),
.A2(n_33),
.B1(n_23),
.B2(n_50),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_151),
.A2(n_163),
.B1(n_56),
.B2(n_100),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_SL g157 ( 
.A1(n_66),
.A2(n_35),
.B(n_41),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_150),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_87),
.A2(n_48),
.B1(n_43),
.B2(n_41),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_159),
.A2(n_77),
.B1(n_83),
.B2(n_82),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_73),
.A2(n_48),
.B1(n_43),
.B2(n_41),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_74),
.B(n_48),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_167),
.B(n_172),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_85),
.B(n_1),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_173),
.B(n_194),
.Y(n_239)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_138),
.B(n_93),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_174),
.A2(n_195),
.B(n_221),
.Y(n_263)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_175),
.Y(n_240)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_176),
.Y(n_271)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_178),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_131),
.B(n_99),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_179),
.B(n_185),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_180),
.B(n_190),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_L g182 ( 
.A1(n_142),
.A2(n_84),
.B1(n_78),
.B2(n_107),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_182),
.A2(n_184),
.B1(n_196),
.B2(n_222),
.Y(n_242)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_115),
.Y(n_183)
);

INVx4_ASAP7_75t_SL g238 ( 
.A(n_183),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_144),
.A2(n_136),
.B1(n_81),
.B2(n_147),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_102),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_186),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_108),
.B(n_96),
.C(n_94),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_188),
.B(n_202),
.Y(n_253)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_119),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_104),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_191),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_112),
.B(n_101),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_192),
.B(n_193),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_114),
.B(n_103),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_98),
.B1(n_97),
.B2(n_57),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_88),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_197),
.B(n_209),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g274 ( 
.A1(n_198),
.A2(n_194),
.B1(n_182),
.B2(n_123),
.Y(n_274)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_199),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_154),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_204),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_116),
.B(n_80),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_232),
.Y(n_245)
);

A2O1A1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_96),
.B(n_2),
.C(n_3),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_139),
.Y(n_203)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_203),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_127),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_205),
.Y(n_283)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_206),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_153),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_160),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_208),
.B(n_212),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_76),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_132),
.Y(n_210)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_210),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_126),
.B(n_69),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_211),
.B(n_223),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_117),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_117),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_213),
.B(n_217),
.Y(n_275)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_121),
.Y(n_214)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_150),
.Y(n_215)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_126),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_216),
.Y(n_278)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_133),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_124),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_226),
.Y(n_257)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_219),
.B(n_229),
.Y(n_256)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_111),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_220),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_124),
.A2(n_65),
.B1(n_59),
.B2(n_96),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_133),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_132),
.B(n_3),
.Y(n_223)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_128),
.B(n_18),
.Y(n_224)
);

AND2x2_ASAP7_75t_SL g267 ( 
.A(n_224),
.B(n_7),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_159),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_225),
.A2(n_231),
.B1(n_11),
.B2(n_12),
.Y(n_287)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_155),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_162),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_228),
.Y(n_264)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_118),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_162),
.Y(n_229)
);

INVx11_ASAP7_75t_L g230 ( 
.A(n_118),
.Y(n_230)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_165),
.A2(n_168),
.B1(n_158),
.B2(n_152),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_128),
.B(n_5),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_233),
.B(n_174),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_165),
.B(n_5),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_8),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_120),
.B(n_6),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_235),
.B(n_8),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_185),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_255),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_173),
.A2(n_158),
.B1(n_152),
.B2(n_120),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_254),
.A2(n_220),
.B1(n_210),
.B2(n_199),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_207),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_187),
.A2(n_130),
.B1(n_109),
.B2(n_110),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_259),
.A2(n_265),
.B1(n_280),
.B2(n_290),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_179),
.B(n_134),
.C(n_111),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_261),
.B(n_288),
.C(n_213),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_181),
.A2(n_140),
.B1(n_123),
.B2(n_121),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_267),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_272),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_190),
.B(n_134),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_270),
.B(n_285),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_177),
.B(n_140),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_274),
.A2(n_287),
.B1(n_13),
.B2(n_14),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_200),
.B(n_9),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_195),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_281),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_224),
.B(n_9),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_289),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_212),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_189),
.B(n_11),
.C(n_12),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_224),
.B(n_12),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_195),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_291),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_244),
.B(n_232),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_292),
.B(n_315),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_253),
.A2(n_224),
.B(n_192),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_294),
.A2(n_283),
.B(n_248),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_239),
.A2(n_184),
.B1(n_225),
.B2(n_224),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_296),
.A2(n_267),
.B1(n_274),
.B2(n_268),
.Y(n_345)
);

BUFx24_ASAP7_75t_L g297 ( 
.A(n_238),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_297),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_271),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_298),
.B(n_301),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_239),
.A2(n_201),
.B1(n_193),
.B2(n_234),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_299),
.A2(n_308),
.B1(n_310),
.B2(n_312),
.Y(n_343)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_250),
.Y(n_300)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_300),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_271),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_252),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_304),
.B(n_314),
.Y(n_358)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_256),
.Y(n_306)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_306),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_239),
.A2(n_202),
.B1(n_188),
.B2(n_203),
.Y(n_308)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_309),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_251),
.A2(n_175),
.B1(n_204),
.B2(n_229),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_253),
.A2(n_176),
.B1(n_214),
.B2(n_208),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_252),
.B(n_205),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_244),
.B(n_183),
.Y(n_315)
);

OAI32xp33_ASAP7_75t_L g316 ( 
.A1(n_237),
.A2(n_233),
.A3(n_227),
.B1(n_226),
.B2(n_178),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_316),
.B(n_328),
.Y(n_374)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_256),
.Y(n_317)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_317),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_242),
.A2(n_243),
.B1(n_265),
.B2(n_237),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_318),
.A2(n_323),
.B1(n_333),
.B2(n_337),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_236),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_319),
.B(n_324),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_245),
.B(n_243),
.Y(n_320)
);

XNOR2x1_ASAP7_75t_L g362 ( 
.A(n_320),
.B(n_329),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_263),
.A2(n_210),
.B(n_218),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_321),
.A2(n_263),
.B(n_284),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_242),
.A2(n_219),
.B1(n_217),
.B2(n_206),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_236),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_246),
.B(n_216),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_325),
.B(n_330),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_326),
.A2(n_282),
.B1(n_271),
.B2(n_266),
.Y(n_369)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_238),
.Y(n_327)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_327),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_255),
.B(n_241),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_246),
.B(n_215),
.Y(n_330)
);

AO22x1_ASAP7_75t_L g331 ( 
.A1(n_259),
.A2(n_230),
.B1(n_228),
.B2(n_186),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_331),
.B(n_335),
.Y(n_383)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_279),
.Y(n_332)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_332),
.Y(n_378)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_334),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_245),
.B(n_15),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_272),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_336),
.A2(n_338),
.B1(n_340),
.B2(n_282),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_281),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_274),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_240),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_339),
.B(n_316),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_274),
.A2(n_17),
.B1(n_267),
.B2(n_289),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_341),
.A2(n_337),
.B(n_322),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_302),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_342),
.B(n_371),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_320),
.B(n_329),
.C(n_305),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_344),
.B(n_352),
.C(n_376),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_345),
.A2(n_348),
.B1(n_357),
.B2(n_305),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_296),
.A2(n_274),
.B1(n_267),
.B2(n_261),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_320),
.B(n_290),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_350),
.B(n_372),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_240),
.C(n_285),
.Y(n_352)
);

XOR2x2_ASAP7_75t_L g353 ( 
.A(n_294),
.B(n_280),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_318),
.A2(n_270),
.B1(n_287),
.B2(n_248),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_311),
.A2(n_273),
.B(n_275),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_359),
.A2(n_361),
.B(n_365),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_311),
.A2(n_273),
.B(n_275),
.Y(n_361)
);

OAI32xp33_ASAP7_75t_L g363 ( 
.A1(n_302),
.A2(n_264),
.A3(n_257),
.B1(n_283),
.B2(n_249),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_368),
.Y(n_389)
);

OAI21xp33_ASAP7_75t_L g419 ( 
.A1(n_364),
.A2(n_334),
.B(n_332),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_321),
.A2(n_262),
.B(n_258),
.Y(n_365)
);

FAx1_ASAP7_75t_SL g367 ( 
.A(n_299),
.B(n_288),
.CI(n_238),
.CON(n_367),
.SN(n_367)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_367),
.B(n_292),
.Y(n_397)
);

OAI32xp33_ASAP7_75t_L g368 ( 
.A1(n_306),
.A2(n_266),
.A3(n_249),
.B1(n_260),
.B2(n_276),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_369),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_328),
.Y(n_371)
);

XNOR2x1_ASAP7_75t_L g372 ( 
.A(n_295),
.B(n_276),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_295),
.B(n_260),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_317),
.B(n_258),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_379),
.C(n_291),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_335),
.B(n_278),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_310),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_325),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_338),
.Y(n_396)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_384),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_375),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_385),
.B(n_400),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_387),
.A2(n_388),
.B1(n_396),
.B2(n_399),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_384),
.A2(n_296),
.B1(n_307),
.B2(n_333),
.Y(n_388)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_347),
.Y(n_393)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_393),
.Y(n_424)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_394),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_370),
.Y(n_395)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_395),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_397),
.B(n_410),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_398),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_380),
.A2(n_307),
.B1(n_323),
.B2(n_293),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_354),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_355),
.A2(n_340),
.B1(n_308),
.B2(n_312),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_403),
.A2(n_413),
.B1(n_420),
.B2(n_352),
.Y(n_438)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_349),
.Y(n_404)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_343),
.A2(n_304),
.B1(n_314),
.B2(n_303),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_405),
.A2(n_374),
.B1(n_348),
.B2(n_343),
.Y(n_423)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_406),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_342),
.B(n_303),
.Y(n_407)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_407),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_358),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_408),
.B(n_411),
.Y(n_436)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_349),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_409),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_346),
.B(n_315),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_351),
.B(n_330),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_378),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_412),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_374),
.A2(n_300),
.B1(n_331),
.B2(n_326),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_358),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_417),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_415),
.A2(n_367),
.B(n_378),
.Y(n_456)
);

NAND3xp33_ASAP7_75t_L g417 ( 
.A(n_371),
.B(n_313),
.C(n_322),
.Y(n_417)
);

BUFx5_ASAP7_75t_L g418 ( 
.A(n_366),
.Y(n_418)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_418),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_363),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_345),
.A2(n_331),
.B1(n_339),
.B2(n_336),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_351),
.B(n_301),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_422),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_360),
.B(n_298),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_423),
.A2(n_428),
.B1(n_429),
.B2(n_431),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_388),
.A2(n_360),
.B1(n_383),
.B2(n_364),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_392),
.A2(n_383),
.B1(n_341),
.B2(n_382),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_392),
.A2(n_361),
.B1(n_359),
.B2(n_377),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_391),
.B(n_362),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_437),
.B(n_440),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_438),
.A2(n_445),
.B1(n_389),
.B2(n_399),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_391),
.B(n_362),
.C(n_344),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_443),
.C(n_407),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_390),
.B(n_376),
.Y(n_440)
);

OAI21xp33_ASAP7_75t_L g484 ( 
.A1(n_441),
.A2(n_456),
.B(n_400),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_368),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_442),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_398),
.B(n_350),
.C(n_372),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_405),
.A2(n_331),
.B1(n_367),
.B2(n_381),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_402),
.A2(n_365),
.B(n_353),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_447),
.A2(n_389),
.B(n_406),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_421),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_454),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_390),
.B(n_379),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_452),
.B(n_403),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_422),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_386),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_455),
.B(n_408),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_401),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_457),
.B(n_465),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_458),
.B(n_477),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_440),
.B(n_387),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_459),
.B(n_475),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_460),
.B(n_430),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_402),
.C(n_415),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_462),
.B(n_463),
.C(n_478),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_386),
.C(n_414),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_397),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_466),
.A2(n_467),
.B1(n_471),
.B2(n_444),
.Y(n_489)
);

CKINVDCx14_ASAP7_75t_R g467 ( 
.A(n_436),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_469),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_432),
.Y(n_470)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_470),
.Y(n_500)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_436),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_425),
.Y(n_473)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_473),
.Y(n_509)
);

XNOR2x1_ASAP7_75t_L g504 ( 
.A(n_474),
.B(n_428),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_452),
.B(n_411),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_425),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_476),
.B(n_480),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_456),
.B(n_410),
.Y(n_477)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_446),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_481),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_431),
.B(n_395),
.C(n_385),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_429),
.B(n_420),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_423),
.B(n_393),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_482),
.B(n_485),
.Y(n_492)
);

INVx13_ASAP7_75t_L g483 ( 
.A(n_432),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_483),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_484),
.A2(n_441),
.B(n_447),
.Y(n_503)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_446),
.Y(n_485)
);

FAx1_ASAP7_75t_SL g487 ( 
.A(n_474),
.B(n_463),
.CI(n_462),
.CON(n_487),
.SN(n_487)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_487),
.B(n_495),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_489),
.A2(n_493),
.B1(n_502),
.B2(n_424),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_461),
.A2(n_449),
.B1(n_433),
.B2(n_444),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_430),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_472),
.A2(n_435),
.B1(n_442),
.B2(n_448),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_496),
.A2(n_506),
.B1(n_507),
.B2(n_451),
.Y(n_511)
);

A2O1A1Ixp33_ASAP7_75t_L g497 ( 
.A1(n_464),
.A2(n_448),
.B(n_441),
.C(n_442),
.Y(n_497)
);

XNOR2x1_ASAP7_75t_L g517 ( 
.A(n_497),
.B(n_504),
.Y(n_517)
);

BUFx12f_ASAP7_75t_SL g499 ( 
.A(n_484),
.Y(n_499)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_499),
.Y(n_522)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_501),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_483),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_503),
.B(n_426),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_464),
.A2(n_445),
.B1(n_396),
.B2(n_416),
.Y(n_506)
);

NOR3xp33_ASAP7_75t_SL g507 ( 
.A(n_477),
.B(n_451),
.C(n_434),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_509),
.A2(n_482),
.B1(n_481),
.B2(n_478),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_510),
.A2(n_528),
.B1(n_500),
.B2(n_505),
.Y(n_540)
);

OAI21xp33_ASAP7_75t_L g531 ( 
.A1(n_511),
.A2(n_506),
.B(n_509),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_494),
.B(n_457),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_512),
.B(n_513),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_494),
.B(n_465),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_508),
.B(n_458),
.C(n_468),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_514),
.B(n_516),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_488),
.B(n_475),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_515),
.B(n_523),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_500),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_505),
.B(n_459),
.Y(n_518)
);

NOR2xp67_ASAP7_75t_SL g543 ( 
.A(n_518),
.B(n_520),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_488),
.C(n_498),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_498),
.B(n_468),
.C(n_373),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_521),
.B(n_525),
.C(n_497),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_496),
.A2(n_434),
.B1(n_426),
.B2(n_424),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_524),
.B(n_527),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_486),
.B(n_373),
.C(n_356),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_503),
.B(n_356),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_529),
.B(n_540),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_522),
.B(n_492),
.Y(n_530)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_530),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_531),
.B(n_539),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_523),
.A2(n_499),
.B(n_490),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_534),
.A2(n_535),
.B(n_366),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_519),
.A2(n_487),
.B(n_501),
.Y(n_535)
);

NOR2x1_ASAP7_75t_L g537 ( 
.A(n_526),
.B(n_504),
.Y(n_537)
);

AOI21x1_ASAP7_75t_L g556 ( 
.A1(n_537),
.A2(n_297),
.B(n_247),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_510),
.A2(n_507),
.B1(n_487),
.B2(n_491),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_525),
.A2(n_394),
.B1(n_412),
.B2(n_409),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_541),
.B(n_521),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_520),
.B(n_309),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_542),
.B(n_309),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_514),
.B(n_404),
.C(n_381),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_544),
.B(n_518),
.C(n_366),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_531),
.A2(n_517),
.B1(n_524),
.B2(n_527),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_546),
.B(n_552),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_537),
.A2(n_517),
.B(n_515),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_547),
.A2(n_530),
.B(n_532),
.Y(n_563)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_548),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_549),
.B(n_536),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_550),
.B(n_534),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_544),
.B(n_327),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_553),
.B(n_555),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_533),
.B(n_418),
.C(n_278),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_556),
.B(n_539),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_559),
.A2(n_563),
.B(n_564),
.Y(n_567)
);

CKINVDCx14_ASAP7_75t_R g568 ( 
.A(n_560),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_562),
.B(n_536),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g564 ( 
.A(n_554),
.B(n_530),
.Y(n_564)
);

A2O1A1O1Ixp25_ASAP7_75t_L g565 ( 
.A1(n_557),
.A2(n_545),
.B(n_551),
.C(n_529),
.D(n_547),
.Y(n_565)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_565),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_561),
.A2(n_554),
.B(n_543),
.Y(n_566)
);

AOI321xp33_ASAP7_75t_L g571 ( 
.A1(n_566),
.A2(n_559),
.A3(n_546),
.B1(n_538),
.B2(n_297),
.C(n_247),
.Y(n_571)
);

A2O1A1O1Ixp25_ASAP7_75t_L g570 ( 
.A1(n_569),
.A2(n_558),
.B(n_549),
.C(n_555),
.D(n_563),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_SL g574 ( 
.A(n_570),
.B(n_571),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_572),
.B(n_567),
.C(n_568),
.Y(n_573)
);

AOI31xp33_ASAP7_75t_L g575 ( 
.A1(n_573),
.A2(n_538),
.A3(n_297),
.B(n_247),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_575),
.B(n_574),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_576),
.B(n_297),
.Y(n_577)
);


endmodule