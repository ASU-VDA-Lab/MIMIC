module real_jpeg_28936_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_1),
.B(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_2),
.B(n_14),
.Y(n_28)
);

HAxp5_ASAP7_75t_SL g16 ( 
.A(n_3),
.B(n_17),
.CON(n_16),
.SN(n_16)
);

AOI21xp5_ASAP7_75t_SL g9 ( 
.A1(n_4),
.A2(n_10),
.B(n_11),
.Y(n_9)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_12),
.Y(n_11)
);

OR2x2_ASAP7_75t_SL g32 ( 
.A(n_5),
.B(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g6 ( 
.A(n_7),
.B(n_20),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_13),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_9),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_18),
.B(n_19),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_14),
.B(n_18),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx24_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_18),
.B(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_19),
.B(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_28),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);


endmodule