module fake_jpeg_28250_n_248 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_16),
.Y(n_40)
);

NAND2x1_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_28),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_43),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_44),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_16),
.B1(n_18),
.B2(n_22),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_52),
.B1(n_56),
.B2(n_60),
.Y(n_84)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

HAxp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_28),
.CON(n_48),
.SN(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_63),
.B(n_33),
.C(n_23),
.Y(n_68)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx6p67_ASAP7_75t_R g80 ( 
.A(n_49),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_42),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_16),
.B1(n_18),
.B2(n_22),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_39),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_18),
.B1(n_22),
.B2(n_19),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_33),
.B1(n_20),
.B2(n_24),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_19),
.B1(n_36),
.B2(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_26),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_19),
.B1(n_29),
.B2(n_30),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

NOR4xp25_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_30),
.C(n_29),
.D(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_66),
.B(n_73),
.Y(n_106)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_68),
.B(n_63),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

NOR2x1_ASAP7_75t_R g99 ( 
.A(n_71),
.B(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_28),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_86),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_20),
.B1(n_24),
.B2(n_32),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_85),
.B1(n_62),
.B2(n_54),
.Y(n_101)
);

BUFx4f_ASAP7_75t_SL g78 ( 
.A(n_58),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_83),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_88),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_20),
.B1(n_24),
.B2(n_32),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_42),
.B(n_38),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_47),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_94),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_50),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_107),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_101),
.A2(n_110),
.B1(n_111),
.B2(n_86),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_54),
.B1(n_50),
.B2(n_61),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_80),
.B1(n_72),
.B2(n_61),
.Y(n_119)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_105),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_53),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_73),
.B(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_66),
.B(n_26),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_28),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_112),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_69),
.A2(n_76),
.B1(n_84),
.B2(n_85),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_54),
.B1(n_61),
.B2(n_46),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_84),
.B(n_23),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_15),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_124),
.B1(n_125),
.B2(n_128),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_116),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_68),
.B(n_75),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_106),
.B(n_97),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_93),
.B1(n_98),
.B2(n_95),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_42),
.C(n_38),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_132),
.C(n_31),
.Y(n_161)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_126),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_127),
.Y(n_148)
);

AO21x2_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_77),
.B(n_80),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_46),
.B1(n_49),
.B2(n_80),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_64),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_80),
.B1(n_49),
.B2(n_44),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_110),
.A2(n_44),
.B1(n_72),
.B2(n_83),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_131),
.B1(n_100),
.B2(n_99),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_38),
.B1(n_20),
.B2(n_24),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_78),
.C(n_58),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_78),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_106),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_90),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_134),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_90),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_137),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_102),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_121),
.A2(n_99),
.B(n_109),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_135),
.B(n_122),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_147),
.B(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_145),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_107),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_101),
.B(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_154),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_153),
.B1(n_70),
.B2(n_25),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_129),
.A2(n_100),
.B1(n_94),
.B2(n_108),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_98),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_31),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_161),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_120),
.C(n_114),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_159),
.C(n_139),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_123),
.B1(n_124),
.B2(n_119),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_163),
.A2(n_165),
.B1(n_176),
.B2(n_178),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_15),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_124),
.B1(n_116),
.B2(n_137),
.Y(n_165)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_175),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_148),
.B(n_152),
.C(n_25),
.Y(n_196)
);

OAI22x1_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_122),
.B1(n_131),
.B2(n_134),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_180),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_127),
.B1(n_130),
.B2(n_82),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_31),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_145),
.B1(n_151),
.B2(n_142),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_156),
.A2(n_25),
.B1(n_2),
.B2(n_4),
.Y(n_180)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_181),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_186),
.C(n_199),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_140),
.C(n_143),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_141),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_189),
.Y(n_211)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_193),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_192),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_141),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_175),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_195),
.B1(n_181),
.B2(n_168),
.Y(n_204)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_197),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_0),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_179),
.C(n_170),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_208),
.C(n_199),
.Y(n_213)
);

A2O1A1O1Ixp25_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_172),
.B(n_170),
.C(n_171),
.D(n_164),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_204),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_178),
.B1(n_165),
.B2(n_163),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_206),
.A2(n_212),
.B1(n_185),
.B2(n_198),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_174),
.C(n_173),
.Y(n_208)
);

BUFx12f_ASAP7_75t_SL g210 ( 
.A(n_187),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_210),
.Y(n_220)
);

OAI321xp33_ASAP7_75t_L g212 ( 
.A1(n_194),
.A2(n_0),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_222),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_215),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g215 ( 
.A(n_210),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_205),
.A2(n_198),
.B1(n_197),
.B2(n_188),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_221),
.B1(n_203),
.B2(n_202),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_211),
.A2(n_184),
.B1(n_193),
.B2(n_5),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_219),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_209),
.A2(n_0),
.B(n_2),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_208),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_14),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_225),
.Y(n_233)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_216),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_229),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_200),
.C(n_201),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_207),
.B1(n_8),
.B2(n_10),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_236)
);

OAI21x1_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_217),
.B(n_222),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_231),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_224),
.A2(n_207),
.B(n_8),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_228),
.C(n_229),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_7),
.B(n_10),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_236),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_235),
.B(n_226),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_237),
.Y(n_242)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_239),
.A2(n_233),
.B(n_228),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_241),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_245),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

OAI321xp33_ASAP7_75t_L g247 ( 
.A1(n_246),
.A2(n_240),
.A3(n_242),
.B1(n_14),
.B2(n_12),
.C(n_13),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_13),
.Y(n_248)
);


endmodule