module fake_jpeg_8618_n_47 (n_3, n_2, n_1, n_0, n_4, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx12_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

FAx1_ASAP7_75t_SL g22 ( 
.A(n_16),
.B(n_19),
.CI(n_21),
.CON(n_22),
.SN(n_22)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_10),
.B1(n_8),
.B2(n_5),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_6),
.A2(n_2),
.B(n_3),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_17),
.B(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_5),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_2),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_4),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_26),
.B1(n_18),
.B2(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_4),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_30),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_8),
.B1(n_16),
.B2(n_7),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_14),
.C(n_15),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_32),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_7),
.C(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_22),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_31),
.B1(n_22),
.B2(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_38),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_23),
.C(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_40),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_4),
.Y(n_40)
);

NOR2x1_ASAP7_75t_SL g41 ( 
.A(n_40),
.B(n_36),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_12),
.B(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_7),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_45),
.B(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_12),
.Y(n_47)
);


endmodule