module fake_netlist_5_950_n_50 (n_8, n_10, n_4, n_5, n_7, n_0, n_12, n_9, n_2, n_13, n_3, n_11, n_6, n_1, n_50);

input n_8;
input n_10;
input n_4;
input n_5;
input n_7;
input n_0;
input n_12;
input n_9;
input n_2;
input n_13;
input n_3;
input n_11;
input n_6;
input n_1;

output n_50;

wire n_29;
wire n_16;
wire n_43;
wire n_47;
wire n_36;
wire n_25;
wire n_18;
wire n_27;
wire n_42;
wire n_22;
wire n_45;
wire n_24;
wire n_28;
wire n_46;
wire n_21;
wire n_44;
wire n_40;
wire n_34;
wire n_38;
wire n_35;
wire n_32;
wire n_41;
wire n_17;
wire n_19;
wire n_37;
wire n_15;
wire n_26;
wire n_30;
wire n_33;
wire n_14;
wire n_48;
wire n_31;
wire n_23;
wire n_49;
wire n_20;
wire n_39;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

OA21x2_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_9),
.B(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_8),
.B(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_20),
.B1(n_15),
.B2(n_16),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_26),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2x1_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_18),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_19),
.Y(n_38)
);

INVxp67_ASAP7_75t_SL g39 ( 
.A(n_35),
.Y(n_39)
);

INVxp67_ASAP7_75t_SL g40 ( 
.A(n_39),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_32),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_42),
.B1(n_44),
.B2(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_46),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_48),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_11),
.B1(n_4),
.B2(n_10),
.Y(n_50)
);


endmodule