module fake_jpeg_32107_n_441 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_441);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_8),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_47),
.B(n_48),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_9),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_50),
.B(n_56),
.Y(n_134)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_54),
.Y(n_139)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_9),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_58),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_7),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_59),
.B(n_65),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_7),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_60),
.B(n_91),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_66),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_29),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_73),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_7),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_74),
.B(n_84),
.Y(n_97)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_76),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_7),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_85),
.B(n_90),
.Y(n_132)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_86),
.B(n_87),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_38),
.A2(n_10),
.B(n_1),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_88),
.A2(n_27),
.B(n_35),
.C(n_33),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_16),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_89),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_38),
.B1(n_28),
.B2(n_37),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_92),
.A2(n_111),
.B1(n_127),
.B2(n_23),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_51),
.A2(n_37),
.B1(n_28),
.B2(n_32),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_101),
.A2(n_119),
.B1(n_124),
.B2(n_138),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_52),
.A2(n_39),
.B1(n_37),
.B2(n_28),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_102),
.A2(n_24),
.B1(n_44),
.B2(n_49),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_53),
.A2(n_37),
.B1(n_18),
.B2(n_45),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_63),
.A2(n_21),
.B1(n_42),
.B2(n_29),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_113),
.A2(n_123),
.B1(n_126),
.B2(n_135),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_47),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_105),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_82),
.A2(n_32),
.B1(n_21),
.B2(n_45),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_68),
.A2(n_42),
.B1(n_29),
.B2(n_32),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_54),
.A2(n_32),
.B1(n_35),
.B2(n_33),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_62),
.A2(n_42),
.B1(n_29),
.B2(n_45),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_48),
.A2(n_39),
.B1(n_42),
.B2(n_30),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_59),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_64),
.A2(n_42),
.B1(n_30),
.B2(n_27),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_89),
.A2(n_91),
.B1(n_69),
.B2(n_79),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_86),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_61),
.A2(n_27),
.B1(n_25),
.B2(n_35),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_71),
.A2(n_42),
.B1(n_25),
.B2(n_33),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_143),
.A2(n_57),
.B1(n_67),
.B2(n_23),
.Y(n_174)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_144),
.Y(n_198)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_146),
.B(n_178),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_147),
.A2(n_96),
.B(n_122),
.Y(n_210)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_148),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_156),
.Y(n_194)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_150),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_60),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_151),
.B(n_154),
.Y(n_218)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_131),
.A2(n_80),
.B1(n_66),
.B2(n_85),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_153),
.A2(n_155),
.B1(n_159),
.B2(n_170),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_25),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_76),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_98),
.B(n_30),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_157),
.B(n_163),
.Y(n_222)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_158),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_92),
.A2(n_90),
.B1(n_83),
.B2(n_81),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_161),
.Y(n_200)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_162),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_114),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_164),
.B(n_187),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_167),
.Y(n_197)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_18),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_172),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_111),
.A2(n_87),
.B1(n_78),
.B2(n_75),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_171),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_127),
.B(n_23),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_174),
.A2(n_175),
.B1(n_184),
.B2(n_188),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_117),
.A2(n_77),
.B1(n_58),
.B2(n_67),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_97),
.B(n_76),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_176),
.Y(n_223)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_177),
.Y(n_233)
);

NAND2x1p5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_57),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_99),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_180),
.Y(n_193)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_186),
.A2(n_93),
.B1(n_125),
.B2(n_110),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_141),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_141),
.A2(n_24),
.B1(n_44),
.B2(n_2),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_136),
.B(n_11),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_189),
.B(n_192),
.Y(n_214)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_95),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_190),
.A2(n_191),
.B1(n_93),
.B2(n_118),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_122),
.A2(n_24),
.B1(n_44),
.B2(n_2),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_94),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_183),
.A2(n_132),
.B1(n_129),
.B2(n_115),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_196),
.A2(n_208),
.B1(n_187),
.B2(n_148),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_146),
.A2(n_130),
.B1(n_118),
.B2(n_96),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_205),
.B(n_95),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_155),
.A2(n_115),
.B1(n_121),
.B2(n_100),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_209),
.Y(n_264)
);

A2O1A1O1Ixp25_ASAP7_75t_L g265 ( 
.A1(n_210),
.A2(n_44),
.B(n_163),
.C(n_167),
.D(n_168),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_151),
.B(n_154),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_227),
.C(n_229),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_169),
.B(n_110),
.C(n_125),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_231),
.B1(n_232),
.B2(n_170),
.Y(n_242)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_189),
.B(n_107),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_178),
.A2(n_146),
.B1(n_166),
.B2(n_147),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_166),
.A2(n_121),
.B1(n_100),
.B2(n_139),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g234 ( 
.A(n_152),
.B(n_142),
.C(n_107),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_158),
.C(n_180),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_195),
.A2(n_173),
.B1(n_178),
.B2(n_172),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_235),
.A2(n_252),
.B1(n_260),
.B2(n_228),
.Y(n_276)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_237),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_164),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_238),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_144),
.Y(n_239)
);

A2O1A1O1Ixp25_ASAP7_75t_L g292 ( 
.A1(n_239),
.A2(n_240),
.B(n_246),
.C(n_255),
.D(n_257),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_145),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_198),
.Y(n_241)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_242),
.A2(n_243),
.B1(n_256),
.B2(n_200),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_214),
.A2(n_159),
.B1(n_171),
.B2(n_160),
.Y(n_243)
);

NOR2x1_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_157),
.Y(n_244)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_244),
.A2(n_211),
.B(n_212),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_192),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_245),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_220),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_199),
.Y(n_247)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_258),
.Y(n_281)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_249),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_177),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_250),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_181),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_251),
.B(n_263),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_253),
.A2(n_265),
.B(n_197),
.Y(n_279)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_254),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_220),
.B(n_179),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_214),
.A2(n_139),
.B1(n_142),
.B2(n_165),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_221),
.B(n_162),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_161),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_202),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_259),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_195),
.A2(n_165),
.B1(n_185),
.B2(n_190),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_207),
.Y(n_261)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_203),
.Y(n_262)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_262),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_202),
.Y(n_263)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_203),
.Y(n_266)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_266),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_222),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_267),
.B(n_233),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_227),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_269),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_184),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_217),
.B(n_0),
.Y(n_270)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_270),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_150),
.C(n_182),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_234),
.C(n_201),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_264),
.A2(n_232),
.B1(n_206),
.B2(n_210),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

OAI32xp33_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_196),
.A3(n_208),
.B1(n_205),
.B2(n_234),
.Y(n_273)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_273),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_276),
.A2(n_293),
.B1(n_242),
.B2(n_257),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_286),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_193),
.C(n_230),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_271),
.C(n_246),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_279),
.B(n_294),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_253),
.A2(n_230),
.B(n_207),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_283),
.A2(n_290),
.B(n_303),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_253),
.A2(n_235),
.B(n_269),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_260),
.A2(n_211),
.B1(n_212),
.B2(n_233),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_295),
.A2(n_237),
.B1(n_247),
.B2(n_254),
.Y(n_315)
);

OAI32xp33_ASAP7_75t_L g297 ( 
.A1(n_263),
.A2(n_200),
.A3(n_226),
.B1(n_204),
.B2(n_225),
.Y(n_297)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_264),
.A2(n_226),
.B1(n_204),
.B2(n_197),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_299),
.A2(n_286),
.B(n_303),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g302 ( 
.A(n_236),
.B(n_215),
.C(n_197),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_248),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_268),
.A2(n_219),
.B(n_216),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_305),
.A2(n_323),
.B1(n_332),
.B2(n_333),
.Y(n_336)
);

BUFx4f_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_307),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_308),
.B(n_328),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_240),
.Y(n_310)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_310),
.Y(n_335)
);

AO22x1_ASAP7_75t_L g311 ( 
.A1(n_286),
.A2(n_271),
.B1(n_252),
.B2(n_265),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_315),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_312),
.B(n_322),
.C(n_279),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_251),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_313),
.B(n_314),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_288),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_321),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_285),
.A2(n_266),
.B1(n_262),
.B2(n_261),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_318),
.A2(n_320),
.B(n_330),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_277),
.A2(n_288),
.B(n_272),
.Y(n_320)
);

OA21x2_ASAP7_75t_L g321 ( 
.A1(n_292),
.A2(n_244),
.B(n_258),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_239),
.C(n_255),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_276),
.A2(n_241),
.B1(n_270),
.B2(n_244),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_284),
.B(n_215),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_325),
.B(n_331),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_249),
.Y(n_326)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_326),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_216),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_328),
.Y(n_337)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_274),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_329),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_290),
.A2(n_216),
.B(n_224),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_284),
.B(n_5),
.Y(n_331)
);

OAI32xp33_ASAP7_75t_L g332 ( 
.A1(n_273),
.A2(n_15),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_293),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_308),
.B(n_281),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_339),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_281),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_306),
.B(n_278),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_344),
.C(n_347),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_305),
.A2(n_298),
.B1(n_304),
.B2(n_280),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_341),
.B(n_342),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_316),
.A2(n_304),
.B1(n_280),
.B2(n_297),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_316),
.A2(n_292),
.B1(n_275),
.B2(n_291),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_346),
.B(n_350),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_283),
.C(n_289),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_322),
.B(n_299),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_348),
.B(n_309),
.C(n_323),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_326),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_319),
.A2(n_274),
.B1(n_275),
.B2(n_291),
.Y(n_350)
);

BUFx24_ASAP7_75t_SL g355 ( 
.A(n_314),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_282),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_307),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_356),
.B(n_307),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_319),
.A2(n_289),
.B1(n_282),
.B2(n_301),
.Y(n_358)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_358),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_359),
.B(n_363),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_339),
.B(n_320),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_361),
.B(n_365),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_340),
.B(n_324),
.C(n_330),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_371),
.C(n_373),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_324),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_352),
.A2(n_327),
.B1(n_333),
.B2(n_311),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_366),
.A2(n_367),
.B1(n_336),
.B2(n_342),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_317),
.Y(n_367)
);

XNOR2x2_ASAP7_75t_SL g368 ( 
.A(n_357),
.B(n_310),
.Y(n_368)
);

AOI31xp33_ASAP7_75t_L g395 ( 
.A1(n_368),
.A2(n_354),
.A3(n_3),
.B(n_4),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_370),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_338),
.B(n_321),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_344),
.C(n_349),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_335),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_376),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_357),
.A2(n_327),
.B(n_311),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_375),
.B(n_379),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_341),
.A2(n_321),
.B(n_315),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_343),
.B(n_329),
.C(n_287),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_378),
.B(n_343),
.C(n_337),
.Y(n_386)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_372),
.Y(n_381)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_381),
.Y(n_396)
);

A2O1A1Ixp33_ASAP7_75t_SL g382 ( 
.A1(n_368),
.A2(n_334),
.B(n_345),
.C(n_332),
.Y(n_382)
);

A2O1A1Ixp33_ASAP7_75t_SL g403 ( 
.A1(n_382),
.A2(n_377),
.B(n_363),
.C(n_371),
.Y(n_403)
);

MAJx2_ASAP7_75t_L g383 ( 
.A(n_364),
.B(n_345),
.C(n_334),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_361),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_386),
.B(n_390),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_369),
.Y(n_398)
);

AOI322xp5_ASAP7_75t_L g390 ( 
.A1(n_367),
.A2(n_336),
.A3(n_346),
.B1(n_351),
.B2(n_358),
.C1(n_353),
.C2(n_350),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_334),
.C(n_351),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_392),
.B(n_393),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_360),
.B(n_362),
.C(n_373),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_365),
.A2(n_301),
.B1(n_296),
.B2(n_287),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_394),
.B(n_12),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_395),
.B(n_15),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_402),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_400),
.B(n_388),
.Y(n_412)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_380),
.Y(n_401)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_401),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_403),
.A2(n_408),
.B1(n_382),
.B2(n_383),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_378),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_386),
.Y(n_414)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_384),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_406),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_359),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_382),
.A2(n_362),
.B1(n_5),
.B2(n_10),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_407),
.B(n_12),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_399),
.A2(n_382),
.B1(n_392),
.B2(n_394),
.Y(n_409)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_409),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_410),
.B(n_408),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_412),
.A2(n_418),
.B(n_419),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_414),
.B(n_417),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_393),
.C(n_385),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_0),
.C(n_13),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_385),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_396),
.B(n_391),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_421),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_415),
.A2(n_403),
.B(n_391),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_423),
.B(n_426),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_409),
.B(n_398),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_424),
.B(n_410),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_413),
.B(n_403),
.C(n_12),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_425),
.B(n_13),
.Y(n_429)
);

NOR2x1_ASAP7_75t_L g428 ( 
.A(n_421),
.B(n_414),
.Y(n_428)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_428),
.Y(n_435)
);

O2A1O1Ixp33_ASAP7_75t_L g433 ( 
.A1(n_429),
.A2(n_411),
.B(n_422),
.C(n_416),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_430),
.A2(n_420),
.B(n_427),
.Y(n_434)
);

AOI21xp33_ASAP7_75t_L g436 ( 
.A1(n_433),
.A2(n_432),
.B(n_431),
.Y(n_436)
);

A2O1A1Ixp33_ASAP7_75t_L g437 ( 
.A1(n_434),
.A2(n_424),
.B(n_426),
.C(n_14),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_436),
.B(n_437),
.C(n_435),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_438),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_439),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_14),
.Y(n_441)
);


endmodule