module fake_jpeg_15963_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx8_ASAP7_75t_SL g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_9),
.Y(n_40)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_58),
.C(n_66),
.Y(n_77)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_41),
.B(n_54),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_9),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_42),
.A2(n_11),
.B(n_12),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_17),
.A2(n_9),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_43),
.B(n_49),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_19),
.B(n_8),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_56),
.B(n_57),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_64),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_63),
.Y(n_103)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_33),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_10),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_67),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_42),
.B(n_21),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_70),
.B(n_84),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_27),
.B1(n_22),
.B2(n_34),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_72),
.A2(n_76),
.B1(n_79),
.B2(n_81),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_22),
.B1(n_34),
.B2(n_32),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_22),
.B1(n_34),
.B2(n_32),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_38),
.B1(n_24),
.B2(n_31),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_26),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_105),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_47),
.A2(n_38),
.B1(n_24),
.B2(n_31),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_88),
.A2(n_89),
.B1(n_100),
.B2(n_102),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_50),
.A2(n_55),
.B1(n_53),
.B2(n_33),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_92),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_59),
.A2(n_33),
.B1(n_0),
.B2(n_2),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_104),
.B1(n_95),
.B2(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_28),
.Y(n_92)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_25),
.B1(n_21),
.B2(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_52),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_99),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_26),
.B1(n_25),
.B2(n_20),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_48),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_48),
.A2(n_4),
.B1(n_6),
.B2(n_10),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_49),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_107),
.B(n_68),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_42),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_108),
.A2(n_99),
.B1(n_73),
.B2(n_101),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_11),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_111),
.B(n_127),
.Y(n_149)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_13),
.B1(n_14),
.B2(n_80),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_103),
.B1(n_106),
.B2(n_71),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_78),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_13),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_123),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_86),
.A2(n_97),
.B1(n_74),
.B2(n_91),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_98),
.B(n_103),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_131),
.B1(n_109),
.B2(n_112),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_128),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_81),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_125),
.B(n_126),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_83),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_133),
.Y(n_153)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_86),
.A2(n_93),
.B1(n_82),
.B2(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_75),
.B(n_72),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_134),
.B(n_137),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_140),
.B(n_112),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_75),
.B(n_93),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_136),
.A2(n_113),
.B(n_110),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_94),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_71),
.C(n_106),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_136),
.C(n_114),
.Y(n_167)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

AOI21x1_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_74),
.B(n_98),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_147),
.B(n_155),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_140),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_144),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_159),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_129),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_156),
.C(n_158),
.Y(n_175)
);

OA21x2_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_123),
.B(n_126),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_109),
.A2(n_115),
.B(n_121),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_167),
.B1(n_149),
.B2(n_162),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_116),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_124),
.B1(n_117),
.B2(n_139),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_160),
.A2(n_161),
.B1(n_163),
.B2(n_146),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_124),
.A2(n_131),
.B1(n_132),
.B2(n_137),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_155),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_125),
.A2(n_128),
.B1(n_133),
.B2(n_118),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_113),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_168),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_114),
.B(n_119),
.C(n_130),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_164),
.B(n_152),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_171),
.B(n_173),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_153),
.Y(n_173)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_164),
.Y(n_179)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_179),
.B(n_186),
.CI(n_173),
.CON(n_192),
.SN(n_192)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_154),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_143),
.A2(n_147),
.B1(n_156),
.B2(n_155),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_183),
.A2(n_145),
.B1(n_150),
.B2(n_168),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_188),
.B1(n_186),
.B2(n_177),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_185),
.A2(n_188),
.B1(n_187),
.B2(n_172),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

A2O1A1O1Ixp25_ASAP7_75t_L g190 ( 
.A1(n_187),
.A2(n_159),
.B(n_144),
.C(n_150),
.D(n_165),
.Y(n_190)
);

AOI221xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_193),
.B1(n_174),
.B2(n_169),
.C(n_184),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_202),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_145),
.C(n_154),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_196),
.C(n_197),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_170),
.C(n_182),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_199),
.A2(n_201),
.B1(n_183),
.B2(n_172),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_170),
.C(n_182),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_171),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_203),
.B(n_174),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_207),
.C(n_193),
.Y(n_215)
);

AO221x1_ASAP7_75t_L g205 ( 
.A1(n_198),
.A2(n_176),
.B1(n_181),
.B2(n_180),
.C(n_178),
.Y(n_205)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_209),
.Y(n_218)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_183),
.B(n_200),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_211),
.A2(n_195),
.B(n_189),
.Y(n_214)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

NOR3xp33_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_211),
.C(n_210),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_212),
.Y(n_219)
);

NAND4xp25_ASAP7_75t_SL g217 ( 
.A(n_205),
.B(n_191),
.C(n_190),
.D(n_194),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_209),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_219),
.B(n_222),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_216),
.B(n_213),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_218),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_223),
.A2(n_225),
.B(n_206),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_215),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_226),
.Y(n_229)
);


endmodule