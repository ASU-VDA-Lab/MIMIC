module fake_ariane_1160_n_110 (n_8, n_3, n_2, n_11, n_7, n_16, n_5, n_14, n_1, n_0, n_12, n_15, n_6, n_13, n_9, n_17, n_4, n_10, n_110);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_16;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_15;
input n_6;
input n_13;
input n_9;
input n_17;
input n_4;
input n_10;

output n_110;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_18;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_19;
wire n_40;
wire n_106;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_109;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_108;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx5p33_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

OA21x2_ASAP7_75t_L g34 ( 
.A1(n_20),
.A2(n_0),
.B(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

AND2x6_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_21),
.B(n_2),
.Y(n_42)
);

OAI21x1_ASAP7_75t_L g43 ( 
.A1(n_23),
.A2(n_10),
.B(n_11),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_30),
.Y(n_48)
);

OAI221xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_27),
.B1(n_19),
.B2(n_28),
.C(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_3),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_40),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_37),
.Y(n_56)
);

AND2x4_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_53),
.Y(n_60)
);

CKINVDCx6p67_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_54),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_52),
.B1(n_49),
.B2(n_54),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_52),
.B(n_46),
.C(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

O2A1O1Ixp5_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_35),
.B(n_39),
.C(n_36),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_57),
.Y(n_68)
);

AO32x2_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_34),
.A3(n_43),
.B1(n_57),
.B2(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_63),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_71),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

OAI21x1_ASAP7_75t_L g79 ( 
.A1(n_75),
.A2(n_67),
.B(n_65),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_73),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_34),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_35),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_R g91 ( 
.A(n_87),
.B(n_89),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_SL g94 ( 
.A1(n_92),
.A2(n_88),
.B(n_79),
.Y(n_94)
);

NAND2x1_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_39),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_95),
.B(n_91),
.Y(n_96)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_79),
.Y(n_99)
);

NAND4xp75_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_34),
.C(n_69),
.D(n_38),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

NAND3xp33_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_101),
.C(n_100),
.Y(n_106)
);

NAND3x1_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_69),
.C(n_57),
.Y(n_107)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_105),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

OAI221xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_38),
.B1(n_106),
.B2(n_105),
.C(n_104),
.Y(n_110)
);


endmodule