module real_jpeg_25532_n_11 (n_8, n_0, n_84, n_93, n_2, n_91, n_10, n_9, n_92, n_6, n_88, n_90, n_7, n_3, n_87, n_5, n_4, n_86, n_85, n_1, n_89, n_11);

input n_8;
input n_0;
input n_84;
input n_93;
input n_2;
input n_91;
input n_10;
input n_9;
input n_92;
input n_6;
input n_88;
input n_90;
input n_7;
input n_3;
input n_87;
input n_5;
input n_4;
input n_86;
input n_85;
input n_1;
input n_89;

output n_11;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_68;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_61;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_16;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_1),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_1),
.B(n_53),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_2),
.B(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_3),
.B(n_31),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_4),
.B(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_7),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_8),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_8),
.B(n_70),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_10),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_20),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_19),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_18),
.Y(n_15)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_17),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_17),
.B(n_54),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B(n_82),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_25),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_73),
.B(n_81),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_69),
.B(n_72),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_63),
.B(n_68),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_36),
.B(n_62),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_56),
.B(n_61),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_52),
.B(n_55),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B(n_51),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_57),
.B(n_58),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_65),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_74),
.B(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_84),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_85),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_86),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_87),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_88),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_89),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_90),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_91),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_92),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_93),
.Y(n_80)
);


endmodule