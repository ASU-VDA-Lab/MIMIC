module fake_netlist_6_4732_n_39 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_9, n_8, n_39);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_9;
input n_8;

output n_39;

wire n_16;
wire n_34;
wire n_24;
wire n_18;
wire n_10;
wire n_21;
wire n_37;
wire n_15;
wire n_33;
wire n_27;
wire n_14;
wire n_38;
wire n_32;
wire n_36;
wire n_22;
wire n_26;
wire n_13;
wire n_35;
wire n_11;
wire n_28;
wire n_17;
wire n_23;
wire n_12;
wire n_20;
wire n_30;
wire n_19;
wire n_29;
wire n_31;
wire n_25;

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g12 ( 
.A(n_6),
.B(n_9),
.Y(n_12)
);

AND2x4_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_2),
.Y(n_13)
);

NOR2xp67_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx5p33_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

AND2x6_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_1),
.Y(n_23)
);

NAND2xp33_ASAP7_75t_SL g24 ( 
.A(n_17),
.B(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_23),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

AOI221xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_18),
.B1(n_10),
.B2(n_11),
.C(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2x1_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_12),
.Y(n_30)
);

AOI221xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_27),
.B1(n_18),
.B2(n_13),
.C(n_16),
.Y(n_31)
);

NOR4xp25_ASAP7_75t_SL g32 ( 
.A(n_30),
.B(n_27),
.C(n_20),
.D(n_15),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OAI211xp5_ASAP7_75t_SL g34 ( 
.A1(n_33),
.A2(n_29),
.B(n_28),
.C(n_19),
.Y(n_34)
);

AOI222xp33_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_13),
.B1(n_20),
.B2(n_14),
.C1(n_26),
.C2(n_30),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

OAI211xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_32),
.B(n_21),
.C(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_36),
.B1(n_13),
.B2(n_3),
.Y(n_39)
);


endmodule