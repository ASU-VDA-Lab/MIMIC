module real_jpeg_26457_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_1),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_1),
.A2(n_66),
.B1(n_67),
.B2(n_149),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_1),
.A2(n_51),
.B1(n_52),
.B2(n_149),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_1),
.A2(n_31),
.B1(n_40),
.B2(n_149),
.Y(n_284)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_5),
.A2(n_32),
.B1(n_51),
.B2(n_52),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_5),
.A2(n_32),
.B1(n_66),
.B2(n_67),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_6),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_6),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_6),
.A2(n_30),
.B1(n_41),
.B2(n_70),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_70),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_7),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_7),
.B(n_104),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_7),
.B(n_62),
.C(n_66),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_7),
.A2(n_51),
.B1(n_52),
.B2(n_152),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_7),
.B(n_58),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_7),
.A2(n_89),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_10),
.A2(n_40),
.B1(n_118),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_10),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_156),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_156),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_10),
.A2(n_66),
.B1(n_67),
.B2(n_156),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_11),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_147),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_11),
.A2(n_51),
.B1(n_52),
.B2(n_147),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_11),
.A2(n_66),
.B1(n_67),
.B2(n_147),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g34 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_13),
.A2(n_35),
.B1(n_51),
.B2(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_13),
.A2(n_35),
.B1(n_66),
.B2(n_67),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_14),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_14),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_14),
.A2(n_46),
.B1(n_118),
.B2(n_121),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_14),
.A2(n_46),
.B1(n_66),
.B2(n_67),
.Y(n_135)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_15),
.Y(n_90)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_15),
.Y(n_169)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_15),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_125),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_123),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_105),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_19),
.B(n_105),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.C(n_85),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_20),
.A2(n_73),
.B1(n_74),
.B2(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_20),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_42),
.B2(n_72),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_21),
.A2(n_22),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_22),
.B(n_43),
.C(n_71),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B(n_33),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_23),
.A2(n_100),
.B1(n_155),
.B2(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_24),
.A2(n_27),
.B(n_153),
.C(n_171),
.Y(n_170)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_25),
.B(n_26),
.C(n_31),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_26),
.A2(n_27),
.B1(n_50),
.B2(n_54),
.Y(n_55)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

HAxp5_ASAP7_75t_SL g243 ( 
.A(n_27),
.B(n_152),
.CON(n_243),
.SN(n_243)
);

NAND3xp33_ASAP7_75t_L g244 ( 
.A(n_27),
.B(n_51),
.C(n_54),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_29),
.Y(n_116)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_30),
.Y(n_120)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_34),
.B(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_38),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_38),
.A2(n_104),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_38),
.A2(n_104),
.B1(n_151),
.B2(n_154),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_38),
.A2(n_104),
.B1(n_162),
.B2(n_284),
.Y(n_283)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_41),
.B(n_152),
.Y(n_153)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_59),
.B2(n_71),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_56),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_45),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_47),
.A2(n_112),
.B(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_47),
.A2(n_49),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g286 ( 
.A1(n_47),
.A2(n_56),
.B(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_58),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_48),
.B(n_57),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_48),
.A2(n_58),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_48),
.A2(n_58),
.B1(n_181),
.B2(n_243),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_49),
.A2(n_77),
.B(n_114),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_49)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_50),
.A2(n_52),
.B(n_243),
.C(n_244),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_52),
.B1(n_62),
.B2(n_64),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_52),
.B(n_197),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_58),
.B(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_59),
.A2(n_71),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_65),
.B(n_68),
.Y(n_59)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_60),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_60),
.A2(n_68),
.B(n_97),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_60),
.A2(n_65),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_60),
.A2(n_65),
.B1(n_201),
.B2(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_60),
.A2(n_80),
.B(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_60),
.A2(n_65),
.B1(n_96),
.B2(n_140),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_65),
.A2(n_82),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_65),
.B(n_152),
.Y(n_234)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_67),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_74),
.A2(n_75),
.B(n_79),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_83),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_81),
.A2(n_84),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_85),
.B(n_331),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_98),
.B(n_99),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_86),
.A2(n_87),
.B1(n_321),
.B2(n_323),
.Y(n_320)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_95),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_88),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_88),
.A2(n_95),
.B1(n_98),
.B2(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_88),
.A2(n_98),
.B1(n_99),
.B2(n_322),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B(n_93),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_89),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_89),
.A2(n_135),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_89),
.B(n_138),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_89),
.A2(n_210),
.B(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_89),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_89),
.A2(n_218),
.B1(n_225),
.B2(n_231),
.Y(n_235)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_90),
.Y(n_187)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_90),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_91),
.Y(n_212)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_94),
.B(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_94),
.A2(n_137),
.B(n_216),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_95),
.Y(n_303)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_99),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B(n_103),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_100),
.A2(n_308),
.B(n_309),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_102),
.B(n_104),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_122),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_115),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_113),
.Y(n_287)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_328),
.B(n_333),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_315),
.B(n_327),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_298),
.B(n_314),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_189),
.B(n_275),
.C(n_297),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_173),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_130),
.B(n_173),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_157),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_141),
.B2(n_142),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_132),
.B(n_142),
.C(n_157),
.Y(n_276)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_139),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_134),
.B(n_139),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_150),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_146),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_152),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_165),
.B2(n_172),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_160),
.B(n_163),
.C(n_172),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_165),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_170),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_187),
.B(n_188),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.C(n_178),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_174),
.B(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_177),
.B(n_178),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.C(n_185),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_179),
.B(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_260)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_216),
.B1(n_217),
.B2(n_219),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_188),
.B(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_274),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_269),
.B(n_273),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_255),
.B(n_268),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_239),
.B(n_254),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_213),
.B(n_238),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_202),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_202),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_198),
.B1(n_199),
.B2(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_209),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_204),
.B(n_207),
.C(n_209),
.Y(n_253)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_210),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_211),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_222),
.B(n_237),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_220),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_220),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_233),
.B(n_236),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_234),
.B(n_235),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_253),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_253),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_249),
.C(n_252),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_242),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_247),
.Y(n_263)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_245),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_251),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_256),
.B(n_257),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_264),
.C(n_266),
.Y(n_272)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_263),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_264),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_272),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_277),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_296),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_288),
.B1(n_294),
.B2(n_295),
.Y(n_278)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_283),
.C(n_285),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_285),
.B2(n_286),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_284),
.Y(n_308)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_288),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_294),
.C(n_296),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_293),
.Y(n_311)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_299),
.B(n_300),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_313),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_304),
.C(n_313),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_311),
.B2(n_312),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_310),
.C(n_312),
.Y(n_326)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_311),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_316),
.B(n_317),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_326),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_324),
.B2(n_325),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_324),
.C(n_326),
.Y(n_329)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_321),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);


endmodule