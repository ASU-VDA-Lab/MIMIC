module fake_jpeg_29014_n_287 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_287);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_287;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_35),
.Y(n_38)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_14),
.B1(n_18),
.B2(n_25),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_24),
.B1(n_25),
.B2(n_17),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_18),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_40),
.B1(n_32),
.B2(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_30),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_26),
.B1(n_34),
.B2(n_36),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_62),
.B1(n_64),
.B2(n_41),
.Y(n_71)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_55),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_27),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_41),
.C(n_43),
.Y(n_67)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_60),
.Y(n_75)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_34),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_SL g61 ( 
.A1(n_46),
.A2(n_30),
.B(n_32),
.C(n_31),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_62),
.B(n_58),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_40),
.B1(n_31),
.B2(n_29),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_26),
.B1(n_25),
.B2(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_43),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_72),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_80),
.B1(n_61),
.B2(n_62),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_42),
.C(n_45),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_42),
.C(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_76),
.Y(n_90)
);

BUFx24_ASAP7_75t_SL g76 ( 
.A(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_79),
.Y(n_106)
);

OA21x2_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_53),
.B(n_48),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_15),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_42),
.C(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_40),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_42),
.B1(n_33),
.B2(n_27),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_103),
.B1(n_107),
.B2(n_67),
.Y(n_117)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_58),
.B1(n_60),
.B2(n_62),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_82),
.B1(n_73),
.B2(n_72),
.Y(n_119)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_61),
.B(n_60),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_99),
.B(n_40),
.Y(n_137)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_20),
.Y(n_130)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

OR2x2_ASAP7_75t_SL g98 ( 
.A(n_68),
.B(n_56),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_72),
.C(n_69),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_56),
.B(n_63),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_109),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_64),
.B1(n_50),
.B2(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_21),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_71),
.A2(n_26),
.B1(n_49),
.B2(n_37),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_57),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_105),
.B(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_111),
.Y(n_153)
);

NOR2x1_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_80),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_112),
.B(n_113),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

OA21x2_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_79),
.B(n_67),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_132),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_116),
.B(n_130),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_125),
.B1(n_135),
.B2(n_102),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_127),
.B1(n_33),
.B2(n_29),
.Y(n_151)
);

CKINVDCx11_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_121),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_32),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_88),
.A2(n_37),
.B1(n_49),
.B2(n_86),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_87),
.A2(n_81),
.B1(n_37),
.B2(n_59),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_95),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_17),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_137),
.B(n_138),
.C(n_101),
.D(n_13),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_90),
.B(n_20),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_37),
.B1(n_81),
.B2(n_59),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_102),
.A2(n_28),
.B1(n_54),
.B2(n_21),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_103),
.B1(n_107),
.B2(n_97),
.Y(n_143)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_30),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_91),
.C(n_119),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_145),
.C(n_150),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_141),
.A2(n_167),
.B1(n_31),
.B2(n_29),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g142 ( 
.A(n_126),
.B(n_91),
.CI(n_106),
.CON(n_142),
.SN(n_142)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_164),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_98),
.C(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_108),
.B1(n_54),
.B2(n_57),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_54),
.C(n_47),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_136),
.A2(n_14),
.B1(n_18),
.B2(n_32),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_159),
.B(n_163),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_47),
.C(n_40),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_19),
.B1(n_18),
.B2(n_14),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_131),
.B1(n_130),
.B2(n_132),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_13),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_115),
.C(n_112),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_113),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_111),
.A2(n_22),
.B1(n_19),
.B2(n_0),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_115),
.B(n_40),
.C(n_32),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_135),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_121),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_169),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_191),
.Y(n_200)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_174),
.Y(n_198)
);

AND2x6_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_138),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_176),
.A2(n_40),
.B(n_31),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_139),
.B(n_133),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_188),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_154),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_180),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_153),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_187),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_111),
.B1(n_125),
.B2(n_129),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_185),
.A2(n_189),
.B1(n_173),
.B2(n_141),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_147),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_129),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_151),
.A2(n_127),
.B1(n_123),
.B2(n_22),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_163),
.B(n_123),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_167),
.Y(n_192)
);

NOR3xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_168),
.C(n_160),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_194),
.A2(n_182),
.B1(n_172),
.B2(n_175),
.Y(n_207)
);

OAI21x1_ASAP7_75t_L g195 ( 
.A1(n_184),
.A2(n_146),
.B(n_142),
.Y(n_195)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_201),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_185),
.A2(n_150),
.B(n_140),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_158),
.C(n_142),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_214),
.C(n_190),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_173),
.A2(n_140),
.B1(n_146),
.B2(n_152),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_212),
.B1(n_213),
.B2(n_1),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_162),
.B(n_2),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_208),
.Y(n_223)
);

XOR2x2_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_191),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_211),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_207),
.A2(n_182),
.B1(n_183),
.B2(n_193),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_174),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_29),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_186),
.A2(n_29),
.B1(n_2),
.B2(n_3),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_189),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_23),
.C(n_4),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_207),
.B1(n_214),
.B2(n_5),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_218),
.B(n_205),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_190),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_226),
.C(n_228),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_209),
.A2(n_181),
.B1(n_176),
.B2(n_194),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_23),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_227),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_23),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_23),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_23),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_204),
.B1(n_213),
.B2(n_199),
.Y(n_241)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_231),
.Y(n_236)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_203),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_229),
.A2(n_211),
.B(n_198),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_235),
.A2(n_219),
.B(n_227),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_201),
.C(n_206),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_244),
.C(n_226),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_212),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_242),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_241),
.A2(n_243),
.B1(n_1),
.B2(n_4),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_1),
.C(n_4),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_245),
.B(n_246),
.Y(n_255)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_249),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_224),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_253),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_217),
.B(n_243),
.Y(n_249)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_252),
.B1(n_7),
.B2(n_8),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_241),
.A2(n_219),
.B1(n_228),
.B2(n_7),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_11),
.C(n_6),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_234),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_11),
.Y(n_264)
);

OA21x2_ASAP7_75t_L g257 ( 
.A1(n_238),
.A2(n_5),
.B(n_6),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_5),
.Y(n_258)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_245),
.C(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_264),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_237),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_265),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_6),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_251),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_7),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_257),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_249),
.B(n_253),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_275),
.B(n_258),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_273),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_247),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_274),
.A2(n_261),
.B(n_8),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_252),
.Y(n_275)
);

AOI21xp33_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_275),
.B(n_271),
.Y(n_277)
);

OAI21x1_ASAP7_75t_SL g281 ( 
.A1(n_277),
.A2(n_280),
.B(n_9),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_278),
.B(n_279),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_272),
.A2(n_7),
.B(n_8),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_282),
.B(n_9),
.Y(n_285)
);

A2O1A1O1Ixp25_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_9),
.B(n_10),
.C(n_11),
.D(n_222),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_283),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_285),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_9),
.Y(n_287)
);


endmodule