module fake_ariane_2314_n_614 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_614);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_614;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_133;
wire n_610;
wire n_205;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_139;
wire n_524;
wire n_391;
wire n_349;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_566;
wire n_578;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_427;
wire n_587;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_588;
wire n_136;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_601;
wire n_565;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_613;
wire n_475;
wire n_135;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_540;
wire n_216;
wire n_544;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_509;
wire n_583;
wire n_306;
wire n_313;
wire n_430;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_337;
wire n_437;
wire n_274;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_132;
wire n_147;
wire n_204;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_508;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_155;
wire n_573;
wire n_531;

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_52),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_72),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_36),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_15),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_0),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_85),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_1),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_50),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_71),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_28),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_7),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_35),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_49),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_11),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_39),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_107),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_59),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_27),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_75),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_93),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_16),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_70),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_24),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_120),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_51),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_76),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_116),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_77),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_86),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_129),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_119),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_48),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_41),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_42),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_97),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_20),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_29),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_60),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_17),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_100),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_106),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_68),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_78),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_44),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_126),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_110),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_79),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_63),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_13),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_98),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_117),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_127),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_83),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_10),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_132),
.B(n_0),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_163),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_176),
.Y(n_201)
);

BUFx2_ASAP7_75t_SL g202 ( 
.A(n_174),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_177),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_183),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_148),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_189),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_192),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

NOR2xp67_ASAP7_75t_L g210 ( 
.A(n_133),
.B(n_1),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_135),
.Y(n_211)
);

BUFx6f_ASAP7_75t_SL g212 ( 
.A(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_140),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_134),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_178),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_136),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_137),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_139),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_143),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_146),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_141),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_147),
.Y(n_223)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_144),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_149),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_168),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_151),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_153),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_156),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_180),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_164),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_168),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_165),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_150),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_152),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_154),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_169),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_173),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_179),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

BUFx2_ASAP7_75t_SL g245 ( 
.A(n_237),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_158),
.B1(n_145),
.B2(n_195),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_219),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_178),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_220),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

OAI22x1_ASAP7_75t_L g258 ( 
.A1(n_200),
.A2(n_181),
.B1(n_190),
.B2(n_191),
.Y(n_258)
);

AND2x4_ASAP7_75t_L g259 ( 
.A(n_209),
.B(n_162),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_210),
.B(n_157),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_159),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_231),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_233),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g273 ( 
.A(n_213),
.B(n_160),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_242),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_201),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_243),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_198),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_197),
.Y(n_279)
);

OA21x2_ASAP7_75t_L g280 ( 
.A1(n_198),
.A2(n_196),
.B(n_194),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_215),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_214),
.B(n_161),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_222),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_202),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_225),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_232),
.A2(n_238),
.B1(n_208),
.B2(n_205),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_212),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_212),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_238),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_203),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_204),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_207),
.B(n_166),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_227),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_232),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_167),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_2),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_288),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_276),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_267),
.B(n_170),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_264),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_251),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_254),
.B(n_2),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_171),
.Y(n_305)
);

AND2x4_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_3),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_251),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_172),
.Y(n_308)
);

AND2x6_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_168),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_245),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_264),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_288),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_289),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g314 ( 
.A(n_248),
.B(n_3),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_249),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_255),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_255),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

NAND3x1_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_4),
.C(n_5),
.Y(n_320)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_289),
.Y(n_321)
);

AND2x4_ASAP7_75t_L g322 ( 
.A(n_281),
.B(n_4),
.Y(n_322)
);

AND2x6_ASAP7_75t_L g323 ( 
.A(n_283),
.B(n_168),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_282),
.B(n_182),
.Y(n_324)
);

AND2x6_ASAP7_75t_L g325 ( 
.A(n_285),
.B(n_184),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_263),
.Y(n_326)
);

OR2x2_ASAP7_75t_SL g327 ( 
.A(n_257),
.B(n_5),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_276),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_291),
.Y(n_329)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_264),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_247),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_264),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_247),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_257),
.Y(n_334)
);

INVx4_ASAP7_75t_SL g335 ( 
.A(n_291),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_291),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_268),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_279),
.B(n_187),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_250),
.Y(n_339)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_271),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_295),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_290),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_250),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_261),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_273),
.B(n_188),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_278),
.B(n_193),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_294),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_286),
.B(n_184),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_278),
.B(n_184),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_292),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_268),
.Y(n_352)
);

INVx5_ASAP7_75t_L g353 ( 
.A(n_259),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_292),
.B(n_184),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_269),
.Y(n_355)
);

BUFx4f_ASAP7_75t_L g356 ( 
.A(n_292),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_356),
.B(n_292),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_299),
.B(n_277),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_355),
.Y(n_359)
);

A2O1A1Ixp33_ASAP7_75t_L g360 ( 
.A1(n_322),
.A2(n_262),
.B(n_252),
.C(n_256),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_259),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_328),
.B(n_290),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_355),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_329),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_348),
.Y(n_366)
);

NAND2x1p5_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_265),
.Y(n_367)
);

OAI221xp5_ASAP7_75t_L g368 ( 
.A1(n_297),
.A2(n_253),
.B1(n_270),
.B2(n_275),
.C(n_272),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_348),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_326),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_315),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_324),
.B(n_266),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_337),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_351),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_352),
.Y(n_375)
);

OAI221xp5_ASAP7_75t_L g376 ( 
.A1(n_356),
.A2(n_253),
.B1(n_269),
.B2(n_246),
.C(n_244),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_331),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_305),
.B(n_342),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_333),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

NAND2x1p5_ASAP7_75t_L g381 ( 
.A(n_345),
.B(n_260),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_343),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_344),
.Y(n_384)
);

OAI221xp5_ASAP7_75t_L g385 ( 
.A1(n_346),
.A2(n_280),
.B1(n_287),
.B2(n_258),
.C(n_9),
.Y(n_385)
);

BUFx8_ASAP7_75t_L g386 ( 
.A(n_303),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_310),
.Y(n_387)
);

NAND2x1p5_ASAP7_75t_L g388 ( 
.A(n_312),
.B(n_280),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_313),
.B(n_184),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_317),
.Y(n_390)
);

AO22x2_ASAP7_75t_L g391 ( 
.A1(n_314),
.A2(n_322),
.B1(n_306),
.B2(n_304),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_318),
.Y(n_392)
);

AND2x6_ASAP7_75t_L g393 ( 
.A(n_304),
.B(n_12),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_334),
.B(n_308),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

OAI221xp5_ASAP7_75t_L g396 ( 
.A1(n_349),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_396)
);

AO22x2_ASAP7_75t_L g397 ( 
.A1(n_306),
.A2(n_8),
.B1(n_14),
.B2(n_18),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_301),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_335),
.B(n_19),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_301),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_353),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_311),
.Y(n_402)
);

NAND2x1p5_ASAP7_75t_L g403 ( 
.A(n_312),
.B(n_21),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_298),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_330),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_296),
.B(n_22),
.Y(n_406)
);

AO22x2_ASAP7_75t_L g407 ( 
.A1(n_320),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_330),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_332),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_347),
.B(n_30),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_332),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_302),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_353),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_307),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_374),
.B(n_321),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_372),
.B(n_338),
.Y(n_416)
);

NAND2xp33_ASAP7_75t_SL g417 ( 
.A(n_404),
.B(n_321),
.Y(n_417)
);

NAND2xp33_ASAP7_75t_SL g418 ( 
.A(n_394),
.B(n_298),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_378),
.B(n_340),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_364),
.B(n_340),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_387),
.B(n_340),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_361),
.B(n_353),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_361),
.B(n_300),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_362),
.B(n_354),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_358),
.B(n_325),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_382),
.B(n_408),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_408),
.B(n_316),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_399),
.B(n_350),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_399),
.B(n_360),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_SL g430 ( 
.A(n_371),
.B(n_327),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_357),
.B(n_325),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_381),
.B(n_323),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_405),
.B(n_323),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_409),
.B(n_323),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_411),
.B(n_323),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_367),
.B(n_309),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_401),
.B(n_413),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_366),
.B(n_309),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_SL g439 ( 
.A(n_398),
.B(n_31),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_369),
.B(n_32),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_359),
.B(n_33),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_391),
.B(n_34),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_391),
.B(n_37),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_363),
.B(n_38),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_377),
.B(n_40),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_373),
.B(n_386),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_386),
.B(n_43),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_400),
.B(n_45),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_365),
.B(n_46),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_402),
.B(n_47),
.Y(n_450)
);

NAND2x1p5_ASAP7_75t_L g451 ( 
.A(n_446),
.B(n_379),
.Y(n_451)
);

NAND2x1p5_ASAP7_75t_L g452 ( 
.A(n_422),
.B(n_383),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_430),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_442),
.A2(n_396),
.B(n_385),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_416),
.B(n_393),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_425),
.B(n_370),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_447),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_445),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_426),
.B(n_393),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_445),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_419),
.Y(n_461)
);

NAND3xp33_ASAP7_75t_L g462 ( 
.A(n_418),
.B(n_368),
.C(n_417),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_449),
.A2(n_410),
.B(n_406),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_393),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_429),
.B(n_423),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_436),
.Y(n_466)
);

AOI21xp33_ASAP7_75t_L g467 ( 
.A1(n_428),
.A2(n_376),
.B(n_397),
.Y(n_467)
);

AO31x2_ASAP7_75t_L g468 ( 
.A1(n_438),
.A2(n_412),
.A3(n_414),
.B(n_375),
.Y(n_468)
);

AO21x2_ASAP7_75t_L g469 ( 
.A1(n_433),
.A2(n_412),
.B(n_389),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_424),
.B(n_380),
.Y(n_470)
);

AOI21x1_ASAP7_75t_L g471 ( 
.A1(n_434),
.A2(n_390),
.B(n_395),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_435),
.A2(n_388),
.B(n_403),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_415),
.A2(n_397),
.B1(n_407),
.B2(n_384),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_437),
.Y(n_474)
);

OAI21x1_ASAP7_75t_SL g475 ( 
.A1(n_439),
.A2(n_392),
.B(n_407),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_431),
.A2(n_53),
.B(n_54),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_432),
.B(n_55),
.Y(n_477)
);

OA21x2_ASAP7_75t_L g478 ( 
.A1(n_463),
.A2(n_441),
.B(n_444),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_470),
.Y(n_479)
);

O2A1O1Ixp33_ASAP7_75t_SL g480 ( 
.A1(n_455),
.A2(n_440),
.B(n_448),
.C(n_450),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_472),
.A2(n_427),
.B(n_420),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_471),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_421),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_456),
.A2(n_56),
.B(n_57),
.Y(n_484)
);

OAI21x1_ASAP7_75t_L g485 ( 
.A1(n_476),
.A2(n_58),
.B(n_61),
.Y(n_485)
);

OAI21x1_ASAP7_75t_L g486 ( 
.A1(n_466),
.A2(n_62),
.B(n_64),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_460),
.B(n_130),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_465),
.B(n_65),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_461),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_128),
.Y(n_490)
);

OA21x2_ASAP7_75t_L g491 ( 
.A1(n_467),
.A2(n_66),
.B(n_67),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_466),
.A2(n_73),
.B(n_74),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_458),
.Y(n_493)
);

AO31x2_ASAP7_75t_L g494 ( 
.A1(n_473),
.A2(n_80),
.A3(n_81),
.B(n_82),
.Y(n_494)
);

OR2x6_ASAP7_75t_L g495 ( 
.A(n_451),
.B(n_88),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_477),
.A2(n_89),
.B(n_91),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_474),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_452),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_468),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_464),
.B(n_95),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_475),
.A2(n_459),
.B(n_462),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_454),
.B(n_96),
.Y(n_502)
);

BUFx4f_ASAP7_75t_SL g503 ( 
.A(n_487),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_487),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_499),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_497),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_489),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_479),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_493),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_482),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_502),
.A2(n_469),
.B(n_457),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_493),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_490),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_498),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_501),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_488),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_488),
.Y(n_517)
);

HB1xp67_ASAP7_75t_SL g518 ( 
.A(n_490),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_495),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_481),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_500),
.Y(n_521)
);

INVx4_ASAP7_75t_SL g522 ( 
.A(n_494),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_500),
.Y(n_523)
);

NAND2x1p5_ASAP7_75t_L g524 ( 
.A(n_483),
.B(n_99),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_494),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_494),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_502),
.B(n_102),
.Y(n_527)
);

OR2x6_ASAP7_75t_L g528 ( 
.A(n_495),
.B(n_104),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_495),
.B(n_105),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_494),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_503),
.B(n_491),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_503),
.B(n_108),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_R g533 ( 
.A(n_518),
.B(n_109),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_R g534 ( 
.A(n_528),
.B(n_491),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_514),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_R g536 ( 
.A(n_528),
.B(n_491),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_506),
.B(n_478),
.Y(n_537)
);

NAND2xp33_ASAP7_75t_R g538 ( 
.A(n_528),
.B(n_478),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_507),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_508),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g541 ( 
.A(n_518),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_512),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_504),
.B(n_513),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_R g544 ( 
.A(n_504),
.B(n_111),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_513),
.B(n_478),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_509),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_R g547 ( 
.A(n_519),
.B(n_112),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_505),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_505),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_510),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_519),
.B(n_492),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_527),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_521),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_539),
.B(n_516),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_540),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_537),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_552),
.B(n_519),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_543),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_531),
.A2(n_522),
.B1(n_519),
.B2(n_526),
.Y(n_559)
);

NOR2x1_ASAP7_75t_SL g560 ( 
.A(n_541),
.B(n_517),
.Y(n_560)
);

INVxp67_ASAP7_75t_SL g561 ( 
.A(n_538),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_548),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_533),
.A2(n_530),
.B1(n_526),
.B2(n_525),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_549),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_535),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_546),
.B(n_542),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_544),
.A2(n_525),
.B1(n_522),
.B2(n_529),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_550),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_558),
.B(n_545),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_565),
.B(n_543),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_560),
.B(n_515),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_566),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_555),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_556),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_564),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_556),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_574),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_576),
.B(n_554),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_572),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_575),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_572),
.B(n_557),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_573),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_572),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_578),
.B(n_570),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_577),
.B(n_571),
.Y(n_585)
);

NOR4xp25_ASAP7_75t_SL g586 ( 
.A(n_581),
.B(n_534),
.C(n_536),
.D(n_561),
.Y(n_586)
);

OAI22xp33_ASAP7_75t_L g587 ( 
.A1(n_579),
.A2(n_561),
.B1(n_583),
.B2(n_582),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_580),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_588),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_585),
.B(n_569),
.Y(n_590)
);

NAND2xp33_ASAP7_75t_SL g591 ( 
.A(n_586),
.B(n_547),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_584),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_587),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_589),
.A2(n_522),
.B1(n_567),
.B2(n_563),
.Y(n_594)
);

INVx1_ASAP7_75t_SL g595 ( 
.A(n_593),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_591),
.A2(n_567),
.B1(n_563),
.B2(n_559),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_595),
.B(n_592),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_596),
.B(n_590),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_597),
.Y(n_599)
);

NOR2x1_ASAP7_75t_L g600 ( 
.A(n_599),
.B(n_598),
.Y(n_600)
);

NOR3xp33_ASAP7_75t_L g601 ( 
.A(n_600),
.B(n_591),
.C(n_532),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_601),
.B(n_594),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_R g603 ( 
.A(n_602),
.B(n_113),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_603),
.Y(n_604)
);

OAI21x1_ASAP7_75t_SL g605 ( 
.A1(n_604),
.A2(n_524),
.B(n_523),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_605),
.A2(n_524),
.B(n_551),
.Y(n_606)
);

AOI31xp33_ASAP7_75t_L g607 ( 
.A1(n_606),
.A2(n_551),
.A3(n_480),
.B(n_553),
.Y(n_607)
);

NOR4xp25_ASAP7_75t_L g608 ( 
.A(n_607),
.B(n_480),
.C(n_520),
.D(n_121),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_608),
.A2(n_568),
.B1(n_486),
.B2(n_562),
.Y(n_609)
);

AOI211xp5_ASAP7_75t_L g610 ( 
.A1(n_608),
.A2(n_511),
.B(n_496),
.C(n_485),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_610),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_609),
.Y(n_612)
);

OAI221xp5_ASAP7_75t_R g613 ( 
.A1(n_611),
.A2(n_114),
.B1(n_115),
.B2(n_122),
.C(n_123),
.Y(n_613)
);

AOI211xp5_ASAP7_75t_L g614 ( 
.A1(n_613),
.A2(n_612),
.B(n_484),
.C(n_125),
.Y(n_614)
);


endmodule