module fake_jpeg_13353_n_49 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_49);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_49;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_1),
.B(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_24),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_20),
.B(n_18),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_26),
.B(n_20),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_20),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_22),
.B1(n_3),
.B2(n_5),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_29),
.B(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_19),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_19),
.C(n_22),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_9),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_38),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_12),
.C(n_13),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_10),
.B(n_11),
.Y(n_40)
);

AO21x1_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_27),
.B(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_39),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_34),
.B1(n_14),
.B2(n_16),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_44),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_46),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_48),
.B(n_45),
.Y(n_49)
);


endmodule