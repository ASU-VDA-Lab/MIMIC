module fake_jpeg_13289_n_476 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_476);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_476;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_56),
.Y(n_154)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_57),
.Y(n_145)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_61),
.B(n_76),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_63),
.Y(n_183)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_66),
.Y(n_141)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_69),
.Y(n_176)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_71),
.Y(n_161)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_73),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_42),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_35),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_77),
.B(n_102),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_78),
.B(n_81),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_79),
.Y(n_151)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_80),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_42),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

BUFx4f_ASAP7_75t_SL g160 ( 
.A(n_83),
.Y(n_160)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_84),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_85),
.B(n_105),
.Y(n_143)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_91),
.Y(n_187)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_92),
.Y(n_173)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_94),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx5_ASAP7_75t_SL g120 ( 
.A(n_95),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g178 ( 
.A(n_96),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_97),
.B(n_101),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_99),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_33),
.B(n_17),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_103),
.B(n_110),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_106),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_44),
.Y(n_105)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_107),
.B(n_108),
.Y(n_155)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_18),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_113),
.Y(n_153)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_111),
.B(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_45),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_19),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_114),
.B(n_115),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_31),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_33),
.B(n_17),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_116),
.B(n_117),
.Y(n_180)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_18),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_77),
.A2(n_109),
.B1(n_106),
.B2(n_99),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_121),
.A2(n_125),
.B1(n_136),
.B2(n_146),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_23),
.B1(n_36),
.B2(n_19),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_56),
.A2(n_40),
.B1(n_36),
.B2(n_23),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_135),
.A2(n_147),
.B1(n_156),
.B2(n_167),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_31),
.B1(n_52),
.B2(n_40),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_60),
.A2(n_31),
.B1(n_54),
.B2(n_53),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_73),
.A2(n_51),
.B1(n_37),
.B2(n_53),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_93),
.A2(n_55),
.B1(n_54),
.B2(n_48),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_148),
.A2(n_152),
.B1(n_157),
.B2(n_165),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_113),
.B(n_55),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_168),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_74),
.A2(n_48),
.B1(n_38),
.B2(n_51),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_87),
.A2(n_37),
.B1(n_38),
.B2(n_6),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_79),
.A2(n_44),
.B1(n_4),
.B2(n_6),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_90),
.A2(n_44),
.B1(n_15),
.B2(n_14),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_95),
.B(n_0),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_171),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_91),
.A2(n_0),
.B1(n_4),
.B2(n_6),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_94),
.Y(n_168)
);

AND2x4_ASAP7_75t_SL g171 ( 
.A(n_59),
.B(n_0),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_96),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_172),
.A2(n_181),
.B1(n_131),
.B2(n_165),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_103),
.A2(n_12),
.B1(n_14),
.B2(n_13),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_179),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_62),
.A2(n_12),
.B1(n_14),
.B2(n_13),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_100),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_66),
.A2(n_11),
.B1(n_15),
.B2(n_68),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_188),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_94),
.A2(n_11),
.B(n_69),
.C(n_83),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_185),
.B(n_157),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_115),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_186),
.B(n_160),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_77),
.A2(n_102),
.B1(n_106),
.B2(n_109),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_102),
.B(n_77),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_193),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_102),
.B(n_77),
.Y(n_193)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

INVx5_ASAP7_75t_SL g281 ( 
.A(n_194),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_197),
.Y(n_282)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_198),
.Y(n_264)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_202),
.Y(n_262)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_118),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_180),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_205),
.B(n_207),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_206),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_143),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_209),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g296 ( 
.A(n_210),
.Y(n_296)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_141),
.Y(n_212)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_212),
.Y(n_265)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_213),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_124),
.B(n_166),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_214),
.Y(n_287)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_141),
.Y(n_215)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_215),
.Y(n_269)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_123),
.Y(n_216)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_216),
.Y(n_270)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_217),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_153),
.B(n_122),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_221),
.B(n_225),
.Y(n_284)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_222),
.Y(n_275)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_223),
.Y(n_278)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_138),
.Y(n_224)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_224),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_166),
.B(n_134),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_177),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_228),
.Y(n_257)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_227),
.Y(n_292)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_145),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_229),
.A2(n_239),
.B1(n_245),
.B2(n_246),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_171),
.B(n_189),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_233),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_171),
.B(n_144),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_231),
.B(n_232),
.Y(n_293)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_142),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_177),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_137),
.B(n_161),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_235),
.Y(n_267)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_175),
.B(n_155),
.C(n_183),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_236),
.B(n_251),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_126),
.B(n_161),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_238),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_147),
.Y(n_238)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_159),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_240),
.A2(n_254),
.B(n_256),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_182),
.B(n_126),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_241),
.B(n_242),
.Y(n_291)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_138),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_145),
.B(n_182),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_243),
.B(n_247),
.Y(n_288)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_139),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_244),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_149),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_151),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_164),
.B(n_154),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_133),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_249),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_133),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_139),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_154),
.B(n_164),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_185),
.B(n_131),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_128),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_191),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_130),
.B(n_191),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_159),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_218),
.A2(n_135),
.B1(n_125),
.B2(n_156),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_263),
.A2(n_271),
.B1(n_285),
.B2(n_289),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_195),
.A2(n_200),
.B1(n_203),
.B2(n_208),
.Y(n_271)
);

AO21x2_ASAP7_75t_L g273 ( 
.A1(n_208),
.A2(n_181),
.B(n_172),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_273),
.A2(n_283),
.B1(n_286),
.B2(n_297),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_279),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_231),
.A2(n_187),
.B1(n_162),
.B2(n_151),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_195),
.A2(n_162),
.B1(n_187),
.B2(n_130),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_231),
.A2(n_128),
.B1(n_129),
.B2(n_176),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_203),
.A2(n_129),
.B1(n_160),
.B2(n_176),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_211),
.A2(n_160),
.B1(n_214),
.B2(n_229),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_219),
.A2(n_236),
.B1(n_211),
.B2(n_196),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_299),
.A2(n_206),
.B1(n_202),
.B2(n_250),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_224),
.A2(n_242),
.B1(n_213),
.B2(n_209),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_300),
.A2(n_244),
.B1(n_246),
.B2(n_245),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_281),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_301),
.B(n_305),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_302),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_299),
.Y(n_303)
);

XNOR2x1_ASAP7_75t_L g343 ( 
.A(n_303),
.B(n_304),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_251),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_281),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_SL g306 ( 
.A(n_297),
.B(n_194),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_306),
.A2(n_315),
.B(n_323),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_204),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_307),
.B(n_319),
.Y(n_355)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_298),
.Y(n_310)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_310),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_220),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_311),
.B(n_318),
.Y(n_349)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_324),
.Y(n_339)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_314),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_272),
.A2(n_255),
.B(n_210),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_210),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_320),
.Y(n_348)
);

INVx13_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_261),
.B(n_270),
.Y(n_318)
);

XNOR2x1_ASAP7_75t_SL g319 ( 
.A(n_293),
.B(n_287),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_288),
.B(n_212),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_271),
.A2(n_199),
.B1(n_201),
.B2(n_215),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_321),
.A2(n_333),
.B1(n_334),
.B2(n_275),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_222),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_328),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_257),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_259),
.B(n_239),
.C(n_232),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_284),
.B(n_197),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_326),
.Y(n_364)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_291),
.Y(n_327)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_295),
.B(n_294),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_273),
.A2(n_283),
.B1(n_279),
.B2(n_290),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_329),
.A2(n_336),
.B1(n_280),
.B2(n_258),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_295),
.B(n_284),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_330),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_294),
.B(n_267),
.C(n_278),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_331),
.B(n_335),
.Y(n_358)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_262),
.Y(n_332)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_332),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_285),
.A2(n_263),
.B1(n_273),
.B2(n_264),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_273),
.A2(n_264),
.B1(n_294),
.B2(n_266),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_266),
.B(n_260),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_273),
.A2(n_300),
.B1(n_269),
.B2(n_292),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_276),
.B(n_292),
.Y(n_337)
);

BUFx24_ASAP7_75t_SL g350 ( 
.A(n_337),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_335),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_344),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_316),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_353),
.A2(n_333),
.B1(n_309),
.B2(n_321),
.Y(n_378)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_310),
.Y(n_354)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_354),
.Y(n_372)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_312),
.Y(n_356)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_356),
.Y(n_390)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_332),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_359),
.Y(n_379)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_320),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_363),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_362),
.A2(n_323),
.B1(n_315),
.B2(n_324),
.Y(n_384)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_313),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_303),
.B(n_278),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_365),
.B(n_307),
.C(n_323),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_352),
.A2(n_334),
.B(n_325),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_367),
.A2(n_381),
.B(n_385),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_387),
.C(n_343),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_366),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_369),
.B(n_374),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_352),
.A2(n_325),
.B(n_328),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_371),
.A2(n_375),
.B(n_367),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_327),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_362),
.A2(n_329),
.B1(n_336),
.B2(n_363),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_349),
.Y(n_376)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_376),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_348),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_384),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_378),
.A2(n_382),
.B1(n_383),
.B2(n_388),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_331),
.Y(n_380)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_380),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_353),
.A2(n_309),
.B(n_304),
.Y(n_381)
);

AOI22x1_ASAP7_75t_L g382 ( 
.A1(n_346),
.A2(n_308),
.B1(n_304),
.B2(n_314),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_361),
.A2(n_330),
.B1(n_322),
.B2(n_319),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_361),
.A2(n_276),
.B(n_317),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_357),
.B(n_258),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_386),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_365),
.B(n_260),
.C(n_268),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_357),
.A2(n_282),
.B1(n_302),
.B2(n_269),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_268),
.Y(n_389)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_389),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_368),
.B(n_343),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_394),
.B(n_401),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_396),
.B(n_398),
.C(n_400),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_368),
.B(n_358),
.C(n_355),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_378),
.A2(n_339),
.B1(n_346),
.B2(n_364),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_407),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_358),
.C(n_355),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_339),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_347),
.C(n_354),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_404),
.C(n_406),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_383),
.B(n_350),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_371),
.B(n_356),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_370),
.A2(n_345),
.B1(n_341),
.B2(n_340),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_408),
.A2(n_375),
.B(n_371),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_370),
.A2(n_345),
.B1(n_341),
.B2(n_340),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_410),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_386),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_392),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_406),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_413),
.A2(n_392),
.B(n_402),
.Y(n_428)
);

MAJx2_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_374),
.C(n_373),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_416),
.C(n_417),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_400),
.B(n_401),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_396),
.B(n_384),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_393),
.B(n_369),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_424),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_408),
.A2(n_377),
.B1(n_386),
.B2(n_388),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_420),
.A2(n_397),
.B1(n_407),
.B2(n_409),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_386),
.C(n_381),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_405),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_425),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_395),
.B(n_373),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_426),
.B(n_427),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_389),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_433),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_413),
.A2(n_402),
.B1(n_391),
.B2(n_397),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_429),
.A2(n_415),
.B1(n_382),
.B2(n_379),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_399),
.Y(n_430)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_430),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_423),
.B(n_404),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_434),
.B(n_416),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_437),
.A2(n_382),
.B1(n_379),
.B2(n_421),
.Y(n_447)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_419),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_438),
.B(n_439),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_412),
.A2(n_420),
.B(n_424),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_445),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_443),
.B(n_429),
.Y(n_450)
);

BUFx24_ASAP7_75t_SL g445 ( 
.A(n_431),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_SL g446 ( 
.A1(n_428),
.A2(n_382),
.B(n_385),
.C(n_372),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_446),
.A2(n_439),
.B(n_438),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_447),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_422),
.C(n_417),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_448),
.B(n_449),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_422),
.C(n_414),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_444),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_451),
.A2(n_457),
.B(n_446),
.Y(n_461)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_441),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_455),
.B(n_456),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_436),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_444),
.A2(n_433),
.B(n_432),
.Y(n_457)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_458),
.Y(n_465)
);

AO21x1_ASAP7_75t_SL g459 ( 
.A1(n_452),
.A2(n_446),
.B(n_437),
.Y(n_459)
);

AOI21xp33_ASAP7_75t_L g464 ( 
.A1(n_459),
.A2(n_462),
.B(n_451),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_461),
.A2(n_450),
.B(n_342),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_454),
.A2(n_446),
.B(n_372),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_390),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_463),
.B(n_379),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_464),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_466),
.B(n_467),
.C(n_460),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_469),
.A2(n_470),
.B(n_467),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_465),
.B(n_421),
.C(n_394),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_471),
.A2(n_472),
.B(n_351),
.Y(n_473)
);

OAI311xp33_ASAP7_75t_L g472 ( 
.A1(n_468),
.A2(n_390),
.A3(n_342),
.B1(n_351),
.C1(n_359),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_473),
.A2(n_274),
.B1(n_262),
.B2(n_265),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_474),
.B(n_265),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_475),
.B(n_296),
.Y(n_476)
);


endmodule