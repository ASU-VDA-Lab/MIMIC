module real_jpeg_27445_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_298, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;
input n_298;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_292;
wire n_288;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_202;
wire n_213;
wire n_128;
wire n_179;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

INVx5_ASAP7_75t_L g85 ( 
.A(n_0),
.Y(n_85)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_1),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_1),
.A2(n_32),
.B1(n_35),
.B2(n_147),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_1),
.A2(n_44),
.B1(n_45),
.B2(n_147),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_1),
.A2(n_73),
.B1(n_74),
.B2(n_147),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_2),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_2),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_76),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_2),
.A2(n_32),
.B1(n_35),
.B2(n_76),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_76),
.Y(n_239)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_4),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_4),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_7),
.A2(n_73),
.B1(n_74),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_7),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_99),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_7),
.A2(n_32),
.B1(n_35),
.B2(n_99),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_99),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_8),
.A2(n_32),
.B1(n_35),
.B2(n_40),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_9),
.A2(n_32),
.B1(n_35),
.B2(n_54),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_10),
.B(n_26),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_10),
.A2(n_25),
.B(n_26),
.C(n_135),
.D(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_10),
.B(n_48),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_10),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_10),
.A2(n_84),
.B(n_152),
.Y(n_172)
);

A2O1A1O1Ixp25_ASAP7_75t_L g182 ( 
.A1(n_10),
.A2(n_44),
.B(n_47),
.C(n_183),
.D(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_10),
.B(n_44),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_10),
.A2(n_45),
.B(n_71),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_10),
.A2(n_73),
.B1(n_74),
.B2(n_167),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_11),
.A2(n_26),
.B(n_28),
.C(n_31),
.Y(n_25)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_12),
.A2(n_46),
.B1(n_73),
.B2(n_74),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_46),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_12),
.A2(n_32),
.B1(n_35),
.B2(n_46),
.Y(n_208)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_15),
.A2(n_73),
.B1(n_74),
.B2(n_122),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_15),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_15),
.A2(n_32),
.B1(n_35),
.B2(n_122),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_122),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_122),
.Y(n_236)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_100),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_20),
.B(n_100),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_81),
.B2(n_82),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_55),
.B1(n_56),
.B2(n_80),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_23),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_23),
.A2(n_24),
.B(n_41),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_36),
.B2(n_38),
.Y(n_24)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_25),
.A2(n_31),
.B1(n_36),
.B2(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_25),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_25),
.A2(n_31),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_26),
.B(n_29),
.Y(n_28)
);

AOI32xp33_ASAP7_75t_L g193 ( 
.A1(n_26),
.A2(n_45),
.A3(n_183),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI32xp33_ASAP7_75t_L g134 ( 
.A1(n_27),
.A2(n_30),
.A3(n_35),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g195 ( 
.A(n_27),
.B(n_52),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_29),
.B(n_32),
.Y(n_136)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_32),
.B(n_85),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_35),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_62),
.B(n_63),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_43),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_45),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_45),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_48),
.B1(n_53),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_47),
.B(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_47),
.A2(n_48),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_52),
.Y(n_194)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_66),
.B2(n_79),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_59),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_62),
.A2(n_63),
.B1(n_94),
.B2(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_62),
.A2(n_212),
.B(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_62),
.A2(n_63),
.B1(n_114),
.B2(n_239),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_63),
.B(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_63),
.A2(n_146),
.B(n_148),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_63),
.B(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_63),
.A2(n_148),
.B(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_67),
.A2(n_120),
.B(n_123),
.Y(n_119)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_68),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_68),
.A2(n_69),
.B1(n_121),
.B2(n_253),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_69),
.B(n_98),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_70),
.A2(n_73),
.B(n_167),
.C(n_226),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_73),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_77),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_77),
.B(n_167),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_77),
.A2(n_97),
.B(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_90),
.B(n_95),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_95),
.B1(n_96),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_83),
.A2(n_91),
.B1(n_92),
.B2(n_104),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B(n_89),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_89),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_84),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_84),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_84),
.B(n_154),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_84),
.A2(n_88),
.B1(n_192),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_84),
.A2(n_88),
.B1(n_111),
.B2(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_86),
.A2(n_159),
.B(n_169),
.Y(n_168)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_SL g112 ( 
.A(n_87),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_87),
.B(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_87),
.A2(n_160),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_88),
.B(n_167),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_103),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.C(n_107),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_101),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_285)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_107),
.B(n_285),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_115),
.C(n_119),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_108),
.A2(n_109),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_110),
.B(n_113),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_115),
.B(n_119),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_116),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_117),
.A2(n_118),
.B(n_203),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_118),
.B(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_118),
.A2(n_202),
.B(n_203),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_123),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI321xp33_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_277),
.A3(n_286),
.B1(n_291),
.B2(n_296),
.C(n_298),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_241),
.C(n_273),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_215),
.B(n_240),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_197),
.B(n_214),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_178),
.B(n_196),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_155),
.B(n_177),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_133),
.B(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_137),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_138),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_150),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_145),
.C(n_150),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_146),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_151),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_164),
.B(n_176),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_163),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_170),
.B(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_171),
.B(n_175),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_166),
.B(n_168),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_179),
.B(n_180),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_189),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_186),
.C(n_189),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_184),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_188),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_198),
.B(n_199),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_209),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_210),
.C(n_211),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_206),
.C(n_207),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_202),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_208),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_216),
.B(n_217),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_228),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_219),
.B(n_220),
.C(n_228),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_220)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_221),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_223),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_227),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_234),
.C(n_237),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_238),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_236),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_242),
.A2(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_260),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_243),
.B(n_260),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_255),
.C(n_259),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_247),
.C(n_254),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_251),
.B2(n_254),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_251),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_259),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_258),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_260)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_269),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_269),
.C(n_272),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_266),
.C(n_267),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_270),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_275),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_284),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_284),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_282),
.C(n_283),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_282),
.Y(n_290)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_287),
.A2(n_292),
.B(n_295),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_288),
.B(n_289),
.Y(n_295)
);


endmodule