module real_jpeg_4491_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_1),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_1),
.Y(n_109)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_1),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_2),
.A2(n_161),
.B1(n_165),
.B2(n_168),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_2),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_2),
.A2(n_168),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_3),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_3),
.Y(n_111)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_3),
.Y(n_131)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_5),
.A2(n_84),
.B1(n_86),
.B2(n_89),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_5),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_5),
.A2(n_48),
.B1(n_89),
.B2(n_226),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_5),
.A2(n_89),
.B1(n_278),
.B2(n_280),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_5),
.A2(n_89),
.B1(n_189),
.B2(n_294),
.Y(n_293)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_6),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_6),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_6),
.Y(n_194)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_6),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_6),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_7),
.A2(n_46),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_7),
.B(n_111),
.C(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_7),
.B(n_74),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_7),
.B(n_154),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_7),
.B(n_250),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_7),
.B(n_183),
.Y(n_329)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_8),
.Y(n_146)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_10),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_10),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_11),
.A2(n_113),
.B1(n_116),
.B2(n_118),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_11),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_11),
.A2(n_118),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_12),
.A2(n_190),
.B1(n_210),
.B2(n_214),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_12),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_13),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_13),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_13),
.A2(n_95),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_13),
.A2(n_95),
.B1(n_319),
.B2(n_321),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_14),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_14),
.A2(n_52),
.B1(n_79),
.B2(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_14),
.A2(n_52),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_14),
.A2(n_52),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_15),
.A2(n_105),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_15),
.Y(n_174)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_236),
.B1(n_237),
.B2(n_360),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_18),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_235),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_197),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_20),
.B(n_197),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_134),
.C(n_176),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_21),
.B(n_357),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_59),
.B2(n_133),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_22),
.B(n_60),
.C(n_100),
.Y(n_217)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_43),
.B(n_49),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_24),
.B(n_51),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_27),
.Y(n_143)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_40),
.B2(n_42),
.Y(n_34)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_37),
.Y(n_140)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_39),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_41),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_46),
.B(n_47),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_46),
.B(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_46),
.A2(n_152),
.B(n_264),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_SL g324 ( 
.A1(n_46),
.A2(n_325),
.B(n_328),
.Y(n_324)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_47),
.A2(n_138),
.A3(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_137)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.Y(n_50)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_58),
.Y(n_196)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_100),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_83),
.B1(n_90),
.B2(n_91),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_61),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_74),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_67),
.B1(n_69),
.B2(n_72),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_65),
.Y(n_336)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_71),
.Y(n_341)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_74),
.Y(n_90)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_79),
.B2(n_81),
.Y(n_74)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_76),
.Y(n_253)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_76),
.Y(n_279)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_77),
.Y(n_320)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_78),
.Y(n_205)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_78),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_80),
.Y(n_282)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_83),
.A2(n_90),
.B(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_90),
.B(n_180),
.Y(n_234)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_91),
.Y(n_233)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

AOI32xp33_ASAP7_75t_L g333 ( 
.A1(n_96),
.A2(n_319),
.A3(n_329),
.B1(n_334),
.B2(n_337),
.Y(n_333)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_99),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_112),
.B(n_119),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_101),
.A2(n_112),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_101),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_101),
.A2(n_119),
.B(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_101),
.A2(n_201),
.B1(n_277),
.B2(n_318),
.Y(n_317)
);

AOI22x1_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_105),
.B1(n_108),
.B2(n_110),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx8_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_107),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_109),
.Y(n_256)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_109),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_126),
.B1(n_129),
.B2(n_132),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_115),
.Y(n_246)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_120),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_128),
.Y(n_321)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_134),
.A2(n_135),
.B1(n_176),
.B2(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_150),
.B2(n_151),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_137),
.B(n_150),
.Y(n_221)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_159),
.B1(n_169),
.B2(n_172),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_152),
.A2(n_259),
.B(n_264),
.Y(n_258)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_153),
.A2(n_160),
.B1(n_186),
.B2(n_193),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_153),
.A2(n_173),
.B1(n_208),
.B2(n_215),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_153),
.B(n_268),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_153),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_162),
.Y(n_269)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_164),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_165),
.B(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_176),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_185),
.C(n_195),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_177),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_184),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_233),
.B(n_234),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_184),
.A2(n_234),
.B(n_324),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_185),
.B(n_195),
.Y(n_351)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_186),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_187),
.Y(n_260)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_225),
.B(n_230),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_220),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_198)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_207),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_201),
.A2(n_244),
.B(n_249),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_201),
.A2(n_249),
.B(n_318),
.Y(n_348)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp33_ASAP7_75t_SL g337 ( 
.A(n_204),
.B(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_216),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_216),
.A2(n_299),
.B(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_217),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_231),
.B2(n_232),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

AOI21x1_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_354),
.B(n_359),
.Y(n_237)
);

AO21x1_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_343),
.B(n_353),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_312),
.B(n_342),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_285),
.B(n_311),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_257),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_242),
.B(n_257),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_251),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_243),
.A2(n_251),
.B1(n_252),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_243),
.Y(n_309)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_274),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_258),
.B(n_275),
.C(n_284),
.Y(n_313)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_259),
.Y(n_305)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_283),
.B2(n_284),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_302),
.B(n_310),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_291),
.B(n_301),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_300),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_300),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_296),
.B(n_299),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_308),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_308),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_313),
.B(n_314),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_330),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_322),
.B2(n_323),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_322),
.C(n_330),
.Y(n_344)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_333),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_333),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx8_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_344),
.B(n_345),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_350),
.B2(n_352),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_348),
.B(n_349),
.C(n_352),
.Y(n_355)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_350),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_355),
.B(n_356),
.Y(n_359)
);


endmodule