module fake_jpeg_14523_n_154 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_154);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_25),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_27),
.Y(n_56)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_16),
.Y(n_45)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_49),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_16),
.B1(n_15),
.B2(n_19),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_19),
.B(n_29),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_53),
.Y(n_73)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_54),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_16),
.B1(n_19),
.B2(n_24),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_55),
.A2(n_29),
.B(n_23),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_56),
.B(n_11),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_39),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_58),
.C(n_68),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_46),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_39),
.B1(n_33),
.B2(n_30),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_60),
.A2(n_49),
.B1(n_42),
.B2(n_50),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_23),
.B(n_22),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_33),
.B1(n_24),
.B2(n_25),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_71),
.B1(n_42),
.B2(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_14),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_49),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_28),
.C(n_27),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_70),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_28),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_22),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_78),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_41),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_53),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_48),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_49),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_86),
.B1(n_71),
.B2(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_87),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_90),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_42),
.Y(n_90)
);

NOR2xp67_ASAP7_75t_R g91 ( 
.A(n_75),
.B(n_73),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_57),
.C(n_67),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_95),
.C(n_100),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_83),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_61),
.C(n_60),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_59),
.B1(n_1),
.B2(n_2),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_54),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_54),
.C(n_18),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_10),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_103),
.B(n_11),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_94),
.B(n_78),
.C(n_95),
.D(n_104),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_114),
.C(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_108),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_105),
.A2(n_88),
.B(n_90),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_18),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_88),
.Y(n_112)
);

XNOR2x2_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_98),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_9),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_18),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_17),
.C(n_21),
.Y(n_128)
);

OAI321xp33_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_106),
.A3(n_117),
.B1(n_109),
.B2(n_107),
.C(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_119),
.B(n_125),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_128),
.Y(n_134)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_127),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_113),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_136),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_123),
.A2(n_109),
.B1(n_113),
.B2(n_116),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_118),
.B(n_17),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_21),
.C(n_3),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_3),
.B(n_4),
.C(n_6),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_135),
.A2(n_124),
.B1(n_121),
.B2(n_122),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_18),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_134),
.C(n_131),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_139),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_141),
.B(n_136),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_142),
.A2(n_135),
.B1(n_138),
.B2(n_13),
.Y(n_146)
);

NAND2x1_ASAP7_75t_SL g143 ( 
.A(n_137),
.B(n_131),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_143),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_140),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_147),
.Y(n_148)
);

OAI31xp33_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_13),
.A3(n_3),
.B(n_21),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_143),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_149),
.A2(n_145),
.B(n_146),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_152),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_148),
.Y(n_154)
);


endmodule