module fake_aes_7668_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_40;
wire n_29;
wire n_39;
INVx1_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_2), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_1), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_14), .B(n_0), .Y(n_20) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_13), .B(n_3), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_12), .Y(n_22) );
CKINVDCx6p67_ASAP7_75t_R g23 ( .A(n_21), .Y(n_23) );
AOI221xp5_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_12), .B1(n_16), .B2(n_11), .C(n_17), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_20), .Y(n_25) );
INVx1_ASAP7_75t_SL g26 ( .A(n_25), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_23), .B(n_19), .Y(n_28) );
NAND2xp5_ASAP7_75t_SL g29 ( .A(n_26), .B(n_24), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
NOR2x1_ASAP7_75t_L g31 ( .A(n_29), .B(n_27), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_32), .B(n_28), .Y(n_33) );
OAI21xp5_ASAP7_75t_L g34 ( .A1(n_31), .A2(n_27), .B(n_21), .Y(n_34) );
AOI221x1_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_13), .B1(n_15), .B2(n_18), .C(n_19), .Y(n_35) );
OAI221xp5_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_18), .B1(n_15), .B2(n_5), .C(n_6), .Y(n_36) );
CKINVDCx5p33_ASAP7_75t_R g37 ( .A(n_34), .Y(n_37) );
OAI211xp5_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_15), .B(n_4), .C(n_5), .Y(n_38) );
AND2x4_ASAP7_75t_L g39 ( .A(n_37), .B(n_15), .Y(n_39) );
AOI322xp5_ASAP7_75t_SL g40 ( .A1(n_36), .A2(n_3), .A3(n_4), .B1(n_15), .B2(n_8), .C1(n_10), .C2(n_7), .Y(n_40) );
AOI22xp5_ASAP7_75t_L g41 ( .A1(n_39), .A2(n_36), .B1(n_38), .B2(n_40), .Y(n_41) );
endmodule