module fake_jpeg_27141_n_295 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_18),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_0),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_44),
.C(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_17),
.B1(n_27),
.B2(n_33),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_19),
.B1(n_34),
.B2(n_41),
.Y(n_82)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_55),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_20),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_63),
.B(n_22),
.Y(n_98)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_33),
.B1(n_31),
.B2(n_23),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_21),
.B1(n_31),
.B2(n_23),
.Y(n_68)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_74),
.B1(n_82),
.B2(n_86),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_71),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_62),
.B1(n_47),
.B2(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_75),
.B(n_91),
.Y(n_113)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_43),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_80),
.A2(n_98),
.B(n_103),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_28),
.B1(n_41),
.B2(n_40),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_36),
.B1(n_39),
.B2(n_18),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_94),
.C(n_29),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_54),
.A2(n_19),
.B1(n_30),
.B2(n_34),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_22),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_90),
.Y(n_133)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_52),
.A2(n_43),
.B1(n_21),
.B2(n_24),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_22),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_50),
.A2(n_43),
.B1(n_28),
.B2(n_30),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_29),
.B1(n_25),
.B2(n_24),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_37),
.Y(n_94)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_22),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

NAND2x1_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_37),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_64),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_104),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_37),
.B(n_24),
.C(n_25),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_88),
.B(n_77),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_103),
.A2(n_67),
.B1(n_45),
.B2(n_65),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_80),
.A2(n_39),
.B1(n_28),
.B2(n_30),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_119),
.B1(n_120),
.B2(n_85),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_80),
.A2(n_39),
.B1(n_36),
.B2(n_18),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_78),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_102),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_29),
.B1(n_25),
.B2(n_24),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_128),
.A2(n_130),
.B1(n_95),
.B2(n_84),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_89),
.A2(n_29),
.B(n_1),
.C(n_3),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_0),
.B(n_1),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_73),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_131),
.B(n_132),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_72),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_69),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_148),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_SL g190 ( 
.A(n_136),
.B(n_137),
.C(n_150),
.Y(n_190)
);

OAI21x1_ASAP7_75t_SL g137 ( 
.A1(n_108),
.A2(n_71),
.B(n_83),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_138),
.B(n_141),
.Y(n_182)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_147),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_116),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_144),
.B(n_158),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_93),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_145),
.B(n_152),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_149),
.B1(n_115),
.B2(n_107),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_82),
.B1(n_77),
.B2(n_84),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_151),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_113),
.B(n_99),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_70),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_153),
.B(n_161),
.Y(n_166)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_126),
.A2(n_105),
.B(n_86),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_157),
.B(n_0),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_125),
.B(n_127),
.C(n_126),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_111),
.A2(n_70),
.B(n_25),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_72),
.Y(n_191)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_96),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_90),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_101),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_107),
.B(n_13),
.Y(n_163)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_163),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_130),
.C(n_123),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_164),
.B(n_177),
.C(n_142),
.Y(n_208)
);

AO22x1_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_129),
.B1(n_128),
.B2(n_95),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_187),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_140),
.B1(n_138),
.B2(n_151),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_162),
.A2(n_129),
.B1(n_115),
.B2(n_123),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_172),
.A2(n_141),
.B1(n_147),
.B2(n_136),
.Y(n_203)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_181),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_129),
.B(n_132),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_174),
.A2(n_176),
.B(n_186),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_121),
.C(n_118),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_143),
.B1(n_135),
.B2(n_146),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_180),
.A2(n_183),
.B1(n_160),
.B2(n_101),
.Y(n_213)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_121),
.B1(n_76),
.B2(n_79),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_72),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_184),
.B(n_191),
.Y(n_210)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_189),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_106),
.Y(n_186)
);

XOR2x2_ASAP7_75t_L g188 ( 
.A(n_137),
.B(n_11),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_188),
.A2(n_12),
.B(n_16),
.Y(n_206)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_157),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_200),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_179),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_194),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_197),
.Y(n_217)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

AOI22x1_ASAP7_75t_SL g198 ( 
.A1(n_188),
.A2(n_135),
.B1(n_157),
.B2(n_156),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_168),
.B1(n_182),
.B2(n_171),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_186),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_199),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_158),
.Y(n_200)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_209),
.B1(n_211),
.B2(n_215),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_213),
.B1(n_175),
.B2(n_198),
.Y(n_222)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_214),
.B(n_186),
.C(n_187),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_142),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_208),
.C(n_210),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_216),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_190),
.B1(n_180),
.B2(n_177),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_190),
.A2(n_169),
.B1(n_176),
.B2(n_192),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_167),
.A2(n_3),
.B(n_4),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_168),
.A2(n_10),
.B1(n_15),
.B2(n_6),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_11),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_215),
.C(n_206),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_221),
.A2(n_229),
.B(n_230),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_222),
.A2(n_235),
.B1(n_202),
.B2(n_11),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_174),
.C(n_183),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_232),
.C(n_234),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_227),
.A2(n_8),
.B1(n_15),
.B2(n_6),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_175),
.C(n_170),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_165),
.C(n_178),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_216),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_239),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_209),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_245),
.Y(n_260)
);

AO21x1_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_201),
.B(n_214),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_203),
.C(n_200),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_241),
.C(n_246),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_211),
.C(n_201),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_249),
.Y(n_254)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_244),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_8),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_223),
.C(n_232),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_235),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_7),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_7),
.C(n_12),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_222),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_255),
.B(n_257),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_256),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_224),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_259),
.B(n_3),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_226),
.B(n_219),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_262),
.C(n_236),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_229),
.B(n_230),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_246),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_239),
.C(n_251),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_267),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_R g266 ( 
.A(n_259),
.B(n_250),
.C(n_245),
.Y(n_266)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_252),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_252),
.C(n_260),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_269),
.B(n_16),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_228),
.B1(n_240),
.B2(n_7),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_255),
.B1(n_254),
.B2(n_257),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g278 ( 
.A(n_272),
.B(n_257),
.CI(n_14),
.CON(n_278),
.SN(n_278)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_258),
.A2(n_14),
.B(n_15),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_16),
.B(n_4),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_268),
.C(n_277),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_279),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_265),
.B(n_270),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_272),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_280),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_284),
.C(n_281),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_266),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_286),
.B(n_276),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_289),
.A2(n_264),
.B(n_285),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_291),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_288),
.B(n_290),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_278),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_278),
.Y(n_295)
);


endmodule