module fake_netlist_6_2488_n_134 (n_41, n_52, n_16, n_45, n_1, n_46, n_34, n_42, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_54, n_27, n_3, n_14, n_38, n_0, n_61, n_39, n_63, n_60, n_59, n_32, n_4, n_36, n_22, n_26, n_55, n_13, n_35, n_11, n_28, n_17, n_23, n_58, n_12, n_20, n_50, n_49, n_7, n_30, n_64, n_2, n_43, n_5, n_19, n_47, n_48, n_29, n_62, n_31, n_25, n_40, n_57, n_53, n_51, n_44, n_56, n_134);

input n_41;
input n_52;
input n_16;
input n_45;
input n_1;
input n_46;
input n_34;
input n_42;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_54;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_61;
input n_39;
input n_63;
input n_60;
input n_59;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_55;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_58;
input n_12;
input n_20;
input n_50;
input n_49;
input n_7;
input n_30;
input n_64;
input n_2;
input n_43;
input n_5;
input n_19;
input n_47;
input n_48;
input n_29;
input n_62;
input n_31;
input n_25;
input n_40;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_134;

wire n_91;
wire n_119;
wire n_88;
wire n_98;
wire n_113;
wire n_73;
wire n_68;
wire n_83;
wire n_101;
wire n_127;
wire n_125;
wire n_77;
wire n_106;
wire n_92;
wire n_133;
wire n_96;
wire n_90;
wire n_105;
wire n_131;
wire n_132;
wire n_102;
wire n_87;
wire n_66;
wire n_99;
wire n_85;
wire n_78;
wire n_84;
wire n_130;
wire n_100;
wire n_129;
wire n_121;
wire n_75;
wire n_109;
wire n_122;
wire n_70;
wire n_120;
wire n_67;
wire n_82;
wire n_110;
wire n_112;
wire n_81;
wire n_76;
wire n_124;
wire n_126;
wire n_94;
wire n_108;
wire n_97;
wire n_116;
wire n_117;
wire n_118;
wire n_65;
wire n_93;
wire n_80;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_115;
wire n_69;
wire n_128;
wire n_79;

AND2x2_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_0),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_4),
.B(n_36),
.Y(n_68)
);

AND2x4_ASAP7_75t_L g69 ( 
.A(n_6),
.B(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_20),
.B(n_44),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

AND2x4_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_10),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_9),
.B(n_50),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_8),
.B(n_15),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_1),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_39),
.B(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_61),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_13),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_12),
.Y(n_86)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_22),
.B(n_21),
.Y(n_87)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_30),
.B(n_19),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_57),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_40),
.B(n_28),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_47),
.A2(n_63),
.B1(n_11),
.B2(n_2),
.Y(n_96)
);

AO22x1_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_14),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_23),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

NOR2x2_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_24),
.Y(n_101)
);

AND2x4_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_25),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_27),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_73),
.B1(n_72),
.B2(n_65),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_79),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

NAND2x1p5_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_29),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

OAI21x1_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_77),
.B(n_95),
.Y(n_111)
);

AO21x2_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_86),
.B(n_75),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_90),
.C(n_84),
.Y(n_113)
);

OAI21x1_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_80),
.B(n_103),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_102),
.A2(n_105),
.B(n_107),
.Y(n_115)
);

OAI21x1_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_85),
.B(n_82),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_74),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_91),
.C(n_93),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

AO21x2_ASAP7_75t_L g123 ( 
.A1(n_119),
.A2(n_111),
.B(n_112),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_120),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

AOI32xp33_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_96),
.A3(n_87),
.B1(n_83),
.B2(n_101),
.Y(n_128)
);

OAI221xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_113),
.B1(n_68),
.B2(n_78),
.C(n_76),
.Y(n_129)
);

OAI31xp33_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_97),
.A3(n_88),
.B(n_123),
.Y(n_130)
);

NAND4xp75_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_128),
.C(n_127),
.D(n_34),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_131),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_59),
.Y(n_133)
);

OA331x2_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_31),
.A3(n_32),
.B1(n_37),
.B2(n_38),
.B3(n_42),
.C1(n_45),
.Y(n_134)
);


endmodule