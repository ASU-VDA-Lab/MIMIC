module fake_jpeg_22912_n_37 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_37);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_37;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_32;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_19),
.A2(n_0),
.B(n_1),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_4),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_24),
.B(n_3),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_2),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_27),
.C(n_28),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_17),
.B1(n_4),
.B2(n_5),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_29),
.B(n_5),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_3),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.B(n_6),
.C(n_7),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_26),
.C(n_17),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_31),
.C(n_10),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_35),
.A2(n_9),
.B(n_11),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_13),
.B(n_14),
.Y(n_37)
);


endmodule