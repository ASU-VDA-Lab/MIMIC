module fake_netlist_5_2480_n_1494 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_451, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_483, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_507, n_119, n_497, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_492, n_171, n_153, n_399, n_341, n_204, n_394, n_250, n_260, n_298, n_320, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_470, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_457, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_145, n_48, n_50, n_337, n_430, n_313, n_88, n_479, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_309, n_30, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_441, n_450, n_312, n_476, n_429, n_345, n_210, n_494, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_407, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_409, n_500, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_391, n_434, n_175, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_52, n_278, n_110, n_1494);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_451;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_483;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_507;
input n_119;
input n_497;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_171;
input n_153;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_260;
input n_298;
input n_320;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_407;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_409;
input n_500;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_391;
input n_434;
input n_175;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1494;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_516;
wire n_933;
wire n_1152;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_1483;
wire n_1314;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_976;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1097;
wire n_1036;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_777;
wire n_1070;
wire n_1030;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_845;
wire n_663;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_901;
wire n_553;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_889;
wire n_973;
wire n_571;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_868;
wire n_639;
wire n_914;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_1194;
wire n_851;
wire n_615;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1233;
wire n_526;
wire n_677;
wire n_1333;
wire n_1121;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_999;
wire n_758;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_1163;
wire n_906;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_1033;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_1383;
wire n_1073;
wire n_662;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_860;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_824;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_950;
wire n_1346;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_912;
wire n_968;
wire n_619;
wire n_1386;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_1432;
wire n_1357;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_1048;
wire n_1288;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1149;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_917;
wire n_601;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_665;
wire n_1440;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1125;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_1067;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_827;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_1235;
wire n_980;
wire n_698;
wire n_703;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_1227;
wire n_840;
wire n_1334;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1330;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_751;
wire n_1083;
wire n_786;
wire n_1142;
wire n_1129;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_517;
wire n_1086;
wire n_796;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_542;
wire n_595;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_379),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_238),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_373),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_100),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_268),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_404),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_283),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_96),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_376),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_270),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_315),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_148),
.Y(n_520)
);

BUFx8_ASAP7_75t_SL g521 ( 
.A(n_318),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_464),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_26),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_497),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_349),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_314),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_201),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_458),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_389),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_230),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_93),
.Y(n_531)
);

BUFx5_ASAP7_75t_L g532 ( 
.A(n_489),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_507),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_282),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_417),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_486),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_350),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_144),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_494),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_36),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_181),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_311),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_22),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_226),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_359),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_324),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_179),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_218),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_83),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_431),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_207),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_84),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_251),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_2),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_465),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_176),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_276),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_396),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_410),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_394),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_135),
.Y(n_561)
);

BUFx10_ASAP7_75t_L g562 ( 
.A(n_203),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_386),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_257),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_194),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_124),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_158),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_504),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_366),
.Y(n_569)
);

CKINVDCx14_ASAP7_75t_R g570 ( 
.A(n_150),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_134),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_498),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_488),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_310),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_362),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_473),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_403),
.Y(n_577)
);

CKINVDCx16_ASAP7_75t_R g578 ( 
.A(n_493),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_500),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_130),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_364),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_472),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_490),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_219),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_197),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_416),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_6),
.Y(n_587)
);

BUFx10_ASAP7_75t_L g588 ( 
.A(n_193),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_405),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_508),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_2),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_351),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_178),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_409),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_61),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_181),
.Y(n_596)
);

BUFx8_ASAP7_75t_SL g597 ( 
.A(n_477),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_167),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_408),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_103),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_375),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_72),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_108),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_407),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_503),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_401),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_481),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_255),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_139),
.Y(n_609)
);

BUFx8_ASAP7_75t_SL g610 ( 
.A(n_470),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_385),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_471),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_421),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_328),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_442),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_111),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_195),
.Y(n_617)
);

BUFx5_ASAP7_75t_L g618 ( 
.A(n_299),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_7),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_154),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_260),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_496),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_190),
.Y(n_623)
);

BUFx10_ASAP7_75t_L g624 ( 
.A(n_86),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_420),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_265),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_312),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_146),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_482),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_96),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_415),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_361),
.Y(n_632)
);

BUFx8_ASAP7_75t_SL g633 ( 
.A(n_412),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_485),
.Y(n_634)
);

BUFx10_ASAP7_75t_L g635 ( 
.A(n_287),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_378),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_25),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_501),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_426),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_445),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_373),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_387),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_225),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_117),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_299),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_502),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_367),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_337),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_381),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_62),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_491),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_47),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_171),
.Y(n_653)
);

INVxp33_ASAP7_75t_SL g654 ( 
.A(n_102),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_157),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_123),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_169),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_236),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_322),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_388),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_346),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_484),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_432),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_61),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_186),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_286),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_145),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_147),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_264),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_288),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_369),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_137),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_53),
.Y(n_673)
);

INVx1_ASAP7_75t_SL g674 ( 
.A(n_69),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_384),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_232),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_62),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_348),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_296),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_391),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_74),
.Y(n_681)
);

BUFx10_ASAP7_75t_L g682 ( 
.A(n_341),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_257),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_191),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_479),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_221),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_11),
.Y(n_687)
);

CKINVDCx14_ASAP7_75t_R g688 ( 
.A(n_433),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_135),
.Y(n_689)
);

BUFx2_ASAP7_75t_L g690 ( 
.A(n_371),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_180),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_220),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_262),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_397),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_255),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_261),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_242),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_60),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_374),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_217),
.Y(n_700)
);

BUFx2_ASAP7_75t_SL g701 ( 
.A(n_303),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_186),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_224),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_237),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_368),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_383),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_406),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_185),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_377),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_304),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_19),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_370),
.Y(n_712)
);

INVxp67_ASAP7_75t_SL g713 ( 
.A(n_43),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_258),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_156),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_244),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_487),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_402),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_345),
.Y(n_719)
);

BUFx10_ASAP7_75t_L g720 ( 
.A(n_183),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_97),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_253),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_308),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_297),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_159),
.Y(n_725)
);

BUFx8_ASAP7_75t_SL g726 ( 
.A(n_363),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_281),
.Y(n_727)
);

INVxp33_ASAP7_75t_SL g728 ( 
.A(n_505),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_495),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_149),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_454),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_317),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_371),
.Y(n_733)
);

BUFx10_ASAP7_75t_L g734 ( 
.A(n_342),
.Y(n_734)
);

CKINVDCx14_ASAP7_75t_R g735 ( 
.A(n_499),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_103),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_438),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_372),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_263),
.Y(n_739)
);

BUFx10_ASAP7_75t_L g740 ( 
.A(n_285),
.Y(n_740)
);

BUFx10_ASAP7_75t_L g741 ( 
.A(n_476),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_365),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_434),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_400),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_172),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_411),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_24),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_229),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_122),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_178),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_196),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_313),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_492),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_474),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_436),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_192),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_456),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_113),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_166),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_116),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_228),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_118),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_395),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_154),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_380),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_235),
.Y(n_766)
);

CKINVDCx16_ASAP7_75t_R g767 ( 
.A(n_128),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_289),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_266),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_392),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_245),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_243),
.Y(n_772)
);

BUFx10_ASAP7_75t_L g773 ( 
.A(n_424),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_478),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_441),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_266),
.Y(n_776)
);

BUFx5_ASAP7_75t_L g777 ( 
.A(n_256),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_382),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_279),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_114),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_85),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_161),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_170),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_227),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_75),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_30),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_129),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_341),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_302),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_483),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_216),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_290),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_393),
.Y(n_793)
);

INVxp33_ASAP7_75t_SL g794 ( 
.A(n_480),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_115),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_338),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_94),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_162),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_339),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_390),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_213),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_243),
.Y(n_802)
);

CKINVDCx14_ASAP7_75t_R g803 ( 
.A(n_297),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_422),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_23),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_475),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_168),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_184),
.Y(n_808)
);

BUFx10_ASAP7_75t_L g809 ( 
.A(n_335),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_100),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_506),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_618),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_514),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_622),
.B(n_1),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_524),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_R g816 ( 
.A(n_688),
.B(n_735),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_651),
.B(n_1),
.Y(n_817)
);

INVxp67_ASAP7_75t_SL g818 ( 
.A(n_535),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_597),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_618),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_522),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_610),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_633),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_777),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_605),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_777),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_777),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_606),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_643),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_521),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_777),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_726),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_636),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_589),
.Y(n_834)
);

INVxp67_ASAP7_75t_SL g835 ( 
.A(n_737),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_767),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_730),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_570),
.B(n_3),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_803),
.B(n_3),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_730),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_528),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_538),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_752),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_752),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_639),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_752),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_533),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_662),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_769),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_728),
.B(n_4),
.Y(n_850)
);

CKINVDCx14_ASAP7_75t_R g851 ( 
.A(n_690),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_794),
.B(n_4),
.Y(n_852)
);

CKINVDCx16_ASAP7_75t_R g853 ( 
.A(n_578),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_718),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_691),
.B(n_0),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_798),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_536),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_654),
.B(n_5),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_539),
.Y(n_859)
);

INVxp67_ASAP7_75t_SL g860 ( 
.A(n_743),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_550),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_559),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_754),
.B(n_5),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_800),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_SL g865 ( 
.A1(n_858),
.A2(n_526),
.B1(n_560),
.B2(n_513),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_836),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_849),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_815),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_833),
.Y(n_869)
);

BUFx12f_ASAP7_75t_L g870 ( 
.A(n_819),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_838),
.A2(n_768),
.B1(n_731),
.B2(n_757),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_837),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_840),
.Y(n_873)
);

OAI21x1_ASAP7_75t_L g874 ( 
.A1(n_812),
.A2(n_573),
.B(n_568),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_853),
.B(n_741),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_843),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_844),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_846),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_856),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_839),
.A2(n_804),
.B1(n_713),
.B2(n_509),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_842),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_864),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_841),
.B(n_646),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_820),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_818),
.B(n_511),
.Y(n_885)
);

NAND2xp33_ASAP7_75t_L g886 ( 
.A(n_855),
.B(n_800),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_814),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_824),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_826),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_847),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_827),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_831),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_851),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_817),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_834),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_835),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_860),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_857),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_859),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_863),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_861),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_862),
.Y(n_902)
);

INVxp67_ASAP7_75t_L g903 ( 
.A(n_829),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_850),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_852),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_816),
.B(n_515),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_906),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_868),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_876),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_894),
.B(n_822),
.Y(n_910)
);

BUFx10_ASAP7_75t_L g911 ( 
.A(n_898),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_887),
.B(n_823),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_893),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_901),
.Y(n_914)
);

OR2x6_ASAP7_75t_L g915 ( 
.A(n_870),
.B(n_701),
.Y(n_915)
);

AO22x2_ASAP7_75t_L g916 ( 
.A1(n_905),
.A2(n_619),
.B1(n_666),
.B2(n_545),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_888),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_889),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_882),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_891),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_882),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_892),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_905),
.B(n_830),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_869),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_890),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_885),
.B(n_632),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_866),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_874),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_893),
.Y(n_929)
);

INVx4_ASAP7_75t_L g930 ( 
.A(n_904),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_883),
.B(n_832),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_878),
.Y(n_932)
);

AND2x2_ASAP7_75t_SL g933 ( 
.A(n_871),
.B(n_541),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_872),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_896),
.B(n_813),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_897),
.B(n_895),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_899),
.B(n_902),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_894),
.B(n_773),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_884),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_873),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_877),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_904),
.Y(n_942)
);

AO22x2_ASAP7_75t_L g943 ( 
.A1(n_900),
.A2(n_714),
.B1(n_751),
.B2(n_674),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_903),
.B(n_821),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_881),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_880),
.B(n_657),
.Y(n_946)
);

INVx8_ASAP7_75t_L g947 ( 
.A(n_886),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_879),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_865),
.Y(n_949)
);

INVx4_ASAP7_75t_L g950 ( 
.A(n_867),
.Y(n_950)
);

INVx4_ASAP7_75t_L g951 ( 
.A(n_875),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_905),
.A2(n_510),
.B1(n_552),
.B2(n_525),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_876),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_887),
.B(n_562),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_898),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_885),
.B(n_642),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_924),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_919),
.B(n_825),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_942),
.B(n_828),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_955),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_935),
.A2(n_848),
.B1(n_854),
.B2(n_845),
.Y(n_961)
);

AO22x2_ASAP7_75t_L g962 ( 
.A1(n_951),
.A2(n_780),
.B1(n_531),
.B2(n_540),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_907),
.A2(n_577),
.B1(n_586),
.B2(n_572),
.Y(n_963)
);

AO22x2_ASAP7_75t_L g964 ( 
.A1(n_933),
.A2(n_543),
.B1(n_547),
.B2(n_523),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_917),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_940),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_954),
.B(n_658),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_927),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_923),
.A2(n_594),
.B1(n_599),
.B2(n_590),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_918),
.B(n_576),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_938),
.B(n_512),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_932),
.B(n_687),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_920),
.Y(n_973)
);

OAI221xp5_ASAP7_75t_L g974 ( 
.A1(n_922),
.A2(n_553),
.B1(n_554),
.B2(n_551),
.C(n_549),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_925),
.A2(n_638),
.B1(n_685),
.B2(n_613),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_936),
.B(n_579),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_908),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_939),
.B(n_604),
.Y(n_978)
);

AO22x2_ASAP7_75t_L g979 ( 
.A1(n_912),
.A2(n_561),
.B1(n_563),
.B2(n_558),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_929),
.B(n_700),
.Y(n_980)
);

NAND2x1p5_ASAP7_75t_L g981 ( 
.A(n_909),
.B(n_582),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_926),
.B(n_562),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_931),
.B(n_583),
.Y(n_983)
);

AO22x2_ASAP7_75t_L g984 ( 
.A1(n_910),
.A2(n_592),
.B1(n_601),
.B2(n_571),
.Y(n_984)
);

OAI221xp5_ASAP7_75t_L g985 ( 
.A1(n_950),
.A2(n_575),
.B1(n_581),
.B2(n_567),
.C(n_564),
.Y(n_985)
);

INVxp33_ASAP7_75t_L g986 ( 
.A(n_944),
.Y(n_986)
);

AO22x2_ASAP7_75t_L g987 ( 
.A1(n_916),
.A2(n_716),
.B1(n_727),
.B2(n_603),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_941),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_956),
.B(n_588),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_948),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_913),
.B(n_947),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_947),
.B(n_516),
.Y(n_992)
);

AO22x2_ASAP7_75t_L g993 ( 
.A1(n_943),
.A2(n_595),
.B1(n_596),
.B2(n_593),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_911),
.B(n_806),
.Y(n_994)
);

AO22x2_ASAP7_75t_L g995 ( 
.A1(n_914),
.A2(n_616),
.B1(n_617),
.B2(n_602),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_915),
.B(n_621),
.Y(n_996)
);

INVxp67_ASAP7_75t_L g997 ( 
.A(n_921),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_953),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_928),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_928),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_924),
.Y(n_1001)
);

AO22x2_ASAP7_75t_L g1002 ( 
.A1(n_949),
.A2(n_679),
.B1(n_683),
.B2(n_664),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_942),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_930),
.B(n_517),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_924),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_930),
.B(n_518),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_934),
.Y(n_1007)
);

AO22x2_ASAP7_75t_L g1008 ( 
.A1(n_949),
.A2(n_697),
.B1(n_712),
.B2(n_678),
.Y(n_1008)
);

AO22x2_ASAP7_75t_L g1009 ( 
.A1(n_949),
.A2(n_648),
.B1(n_649),
.B2(n_647),
.Y(n_1009)
);

AO22x2_ASAP7_75t_L g1010 ( 
.A1(n_949),
.A2(n_656),
.B1(n_661),
.B2(n_650),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_924),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_942),
.B(n_624),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_946),
.A2(n_811),
.B1(n_631),
.B2(n_634),
.Y(n_1013)
);

OAI221xp5_ASAP7_75t_L g1014 ( 
.A1(n_952),
.A2(n_795),
.B1(n_698),
.B2(n_702),
.C(n_689),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_924),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_924),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_924),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_937),
.B(n_629),
.Y(n_1018)
);

AO22x2_ASAP7_75t_L g1019 ( 
.A1(n_949),
.A2(n_704),
.B1(n_705),
.B2(n_684),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_930),
.B(n_607),
.Y(n_1020)
);

AO22x2_ASAP7_75t_L g1021 ( 
.A1(n_949),
.A2(n_788),
.B1(n_715),
.B2(n_711),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_937),
.B(n_707),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_945),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_924),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_983),
.B(n_612),
.Y(n_1025)
);

NAND2xp33_ASAP7_75t_SL g1026 ( 
.A(n_960),
.B(n_585),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_999),
.B(n_717),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_SL g1028 ( 
.A(n_1013),
.B(n_623),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_1023),
.B(n_1004),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_1006),
.B(n_625),
.Y(n_1030)
);

NAND2xp33_ASAP7_75t_SL g1031 ( 
.A(n_967),
.B(n_1003),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1012),
.B(n_624),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1018),
.B(n_729),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_SL g1034 ( 
.A(n_994),
.B(n_628),
.Y(n_1034)
);

NAND2xp33_ASAP7_75t_SL g1035 ( 
.A(n_959),
.B(n_659),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_1022),
.B(n_640),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_957),
.B(n_663),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_966),
.B(n_753),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1001),
.B(n_775),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1005),
.B(n_790),
.Y(n_1040)
);

NAND2xp33_ASAP7_75t_SL g1041 ( 
.A(n_982),
.B(n_667),
.Y(n_1041)
);

NAND2xp33_ASAP7_75t_SL g1042 ( 
.A(n_989),
.B(n_680),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_1011),
.B(n_744),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1015),
.B(n_746),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_992),
.B(n_635),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1016),
.B(n_755),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_1017),
.B(n_1024),
.Y(n_1047)
);

NAND2xp33_ASAP7_75t_SL g1048 ( 
.A(n_990),
.B(n_693),
.Y(n_1048)
);

NAND2xp33_ASAP7_75t_SL g1049 ( 
.A(n_968),
.B(n_710),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_971),
.B(n_963),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1000),
.B(n_774),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_991),
.B(n_635),
.Y(n_1052)
);

NAND2xp33_ASAP7_75t_SL g1053 ( 
.A(n_978),
.B(n_738),
.Y(n_1053)
);

NAND2xp33_ASAP7_75t_SL g1054 ( 
.A(n_976),
.B(n_747),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_969),
.B(n_965),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_973),
.B(n_961),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_988),
.B(n_1007),
.Y(n_1057)
);

NAND2xp33_ASAP7_75t_SL g1058 ( 
.A(n_1020),
.B(n_771),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_977),
.B(n_615),
.Y(n_1059)
);

NAND2xp33_ASAP7_75t_SL g1060 ( 
.A(n_998),
.B(n_807),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_972),
.B(n_970),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_958),
.B(n_615),
.Y(n_1062)
);

NAND2xp33_ASAP7_75t_SL g1063 ( 
.A(n_975),
.B(n_519),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_984),
.B(n_532),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_997),
.B(n_555),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_981),
.B(n_520),
.Y(n_1066)
);

NAND2xp33_ASAP7_75t_SL g1067 ( 
.A(n_979),
.B(n_527),
.Y(n_1067)
);

NAND2xp33_ASAP7_75t_SL g1068 ( 
.A(n_979),
.B(n_529),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_962),
.B(n_665),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_964),
.B(n_530),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1002),
.B(n_534),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_964),
.B(n_537),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1008),
.B(n_542),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1021),
.B(n_544),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_987),
.B(n_546),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_993),
.B(n_548),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_996),
.B(n_723),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_993),
.B(n_556),
.Y(n_1078)
);

NAND2xp33_ASAP7_75t_SL g1079 ( 
.A(n_1009),
.B(n_557),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_1014),
.B(n_565),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_1010),
.B(n_566),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_1019),
.B(n_569),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_1019),
.B(n_574),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_985),
.B(n_584),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_995),
.B(n_587),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_974),
.B(n_591),
.Y(n_1086)
);

NAND2xp33_ASAP7_75t_SL g1087 ( 
.A(n_986),
.B(n_598),
.Y(n_1087)
);

NAND2xp33_ASAP7_75t_SL g1088 ( 
.A(n_986),
.B(n_600),
.Y(n_1088)
);

AND2x2_ASAP7_75t_SL g1089 ( 
.A(n_959),
.B(n_580),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_983),
.B(n_608),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_983),
.B(n_609),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_983),
.B(n_611),
.Y(n_1092)
);

NAND2xp33_ASAP7_75t_SL g1093 ( 
.A(n_986),
.B(n_614),
.Y(n_1093)
);

NAND2xp33_ASAP7_75t_SL g1094 ( 
.A(n_986),
.B(n_620),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_983),
.B(n_626),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_980),
.B(n_792),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_983),
.B(n_637),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_983),
.B(n_641),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_983),
.B(n_644),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_983),
.B(n_645),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_983),
.B(n_653),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_983),
.B(n_655),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_983),
.B(n_660),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_983),
.B(n_668),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_983),
.B(n_669),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_983),
.B(n_670),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_983),
.B(n_671),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_983),
.B(n_672),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_983),
.B(n_675),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_983),
.B(n_677),
.Y(n_1110)
);

NAND2xp33_ASAP7_75t_SL g1111 ( 
.A(n_986),
.B(n_681),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_983),
.B(n_686),
.Y(n_1112)
);

INVx5_ASAP7_75t_L g1113 ( 
.A(n_1077),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_1035),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1055),
.A2(n_1050),
.B(n_1061),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_1049),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1097),
.A2(n_745),
.B(n_739),
.Y(n_1117)
);

AOI211x1_ASAP7_75t_L g1118 ( 
.A1(n_1081),
.A2(n_1082),
.B(n_1083),
.C(n_1056),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1028),
.A2(n_758),
.B(n_759),
.C(n_756),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_1089),
.B(n_692),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1047),
.A2(n_695),
.B1(n_696),
.B2(n_694),
.Y(n_1121)
);

AO31x2_ASAP7_75t_L g1122 ( 
.A1(n_1064),
.A2(n_762),
.A3(n_765),
.B(n_760),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1045),
.B(n_699),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_1029),
.B(n_703),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1051),
.A2(n_708),
.B1(n_709),
.B2(n_706),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1057),
.A2(n_791),
.B(n_786),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1038),
.A2(n_1040),
.B(n_1039),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1027),
.A2(n_793),
.B(n_630),
.Y(n_1128)
);

O2A1O1Ixp5_ASAP7_75t_SL g1129 ( 
.A1(n_1076),
.A2(n_720),
.B(n_734),
.C(n_682),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1033),
.A2(n_652),
.B(n_627),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1112),
.A2(n_676),
.B(n_673),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_1077),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1037),
.A2(n_399),
.B(n_398),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1026),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_1034),
.A2(n_721),
.B(n_722),
.C(n_719),
.Y(n_1135)
);

BUFx4f_ASAP7_75t_L g1136 ( 
.A(n_1032),
.Y(n_1136)
);

BUFx12f_ASAP7_75t_L g1137 ( 
.A(n_1096),
.Y(n_1137)
);

AOI221x1_ASAP7_75t_L g1138 ( 
.A1(n_1067),
.A2(n_7),
.B1(n_0),
.B2(n_6),
.C(n_8),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_L g1139 ( 
.A(n_1087),
.B(n_725),
.C(n_724),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1054),
.A2(n_1058),
.B1(n_1053),
.B2(n_1041),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_1088),
.B(n_733),
.C(n_732),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1044),
.B(n_736),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_1052),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1046),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1042),
.A2(n_748),
.B1(n_749),
.B2(n_742),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1031),
.B(n_750),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1090),
.A2(n_763),
.B1(n_764),
.B2(n_761),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1078),
.A2(n_734),
.B(n_740),
.C(n_720),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1075),
.A2(n_809),
.B(n_740),
.C(n_766),
.Y(n_1149)
);

AO22x2_ASAP7_75t_L g1150 ( 
.A1(n_1085),
.A2(n_809),
.B1(n_13),
.B2(n_20),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1059),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1091),
.B(n_1092),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1062),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_1071),
.Y(n_1154)
);

NAND3x1_ASAP7_75t_L g1155 ( 
.A(n_1069),
.B(n_772),
.C(n_770),
.Y(n_1155)
);

INVx5_ASAP7_75t_L g1156 ( 
.A(n_1060),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1065),
.Y(n_1157)
);

OAI22x1_ASAP7_75t_L g1158 ( 
.A1(n_1070),
.A2(n_778),
.B1(n_779),
.B2(n_776),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1025),
.A2(n_782),
.B1(n_783),
.B2(n_781),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1073),
.Y(n_1160)
);

AO21x1_ASAP7_75t_L g1161 ( 
.A1(n_1068),
.A2(n_9),
.B(n_10),
.Y(n_1161)
);

OA21x2_ASAP7_75t_L g1162 ( 
.A1(n_1043),
.A2(n_785),
.B(n_784),
.Y(n_1162)
);

NAND3xp33_ASAP7_75t_L g1163 ( 
.A(n_1093),
.B(n_789),
.C(n_787),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1074),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1095),
.B(n_796),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1048),
.B(n_797),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1098),
.A2(n_801),
.B1(n_802),
.B2(n_799),
.Y(n_1167)
);

AO21x1_ASAP7_75t_L g1168 ( 
.A1(n_1079),
.A2(n_11),
.B(n_12),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_1094),
.Y(n_1169)
);

OAI22x1_ASAP7_75t_L g1170 ( 
.A1(n_1072),
.A2(n_808),
.B1(n_810),
.B2(n_805),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1030),
.A2(n_414),
.B(n_413),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1080),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1036),
.A2(n_419),
.B(n_418),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1099),
.A2(n_425),
.B(n_423),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1100),
.B(n_14),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1086),
.Y(n_1176)
);

AOI31xp33_ASAP7_75t_L g1177 ( 
.A1(n_1111),
.A2(n_17),
.A3(n_15),
.B(n_16),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1113),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1132),
.Y(n_1179)
);

OAI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1140),
.A2(n_1084),
.B1(n_1102),
.B2(n_1101),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_L g1181 ( 
.A(n_1117),
.B(n_1063),
.C(n_1103),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1137),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_1154),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_1164),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_1175),
.B(n_1105),
.C(n_1104),
.Y(n_1185)
);

OA21x2_ASAP7_75t_L g1186 ( 
.A1(n_1127),
.A2(n_1107),
.B(n_1106),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1176),
.A2(n_1108),
.B(n_1110),
.C(n_1109),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1164),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1144),
.A2(n_1066),
.B(n_427),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_1136),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1122),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1143),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1122),
.Y(n_1193)
);

NAND2x1p5_ASAP7_75t_L g1194 ( 
.A(n_1156),
.B(n_428),
.Y(n_1194)
);

INVx2_ASAP7_75t_SL g1195 ( 
.A(n_1156),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1172),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1114),
.A2(n_21),
.B1(n_18),
.B2(n_19),
.Y(n_1197)
);

AO31x2_ASAP7_75t_L g1198 ( 
.A1(n_1168),
.A2(n_1161),
.A3(n_1138),
.B(n_1158),
.Y(n_1198)
);

AOI21xp33_ASAP7_75t_L g1199 ( 
.A1(n_1123),
.A2(n_21),
.B(n_22),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1152),
.A2(n_430),
.B(n_429),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1116),
.B(n_24),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_1134),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_SL g1203 ( 
.A1(n_1150),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1153),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1160),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1118),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1206)
);

OA21x2_ASAP7_75t_L g1207 ( 
.A1(n_1128),
.A2(n_437),
.B(n_435),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1142),
.B(n_34),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1151),
.Y(n_1209)
);

BUFx12f_ASAP7_75t_L g1210 ( 
.A(n_1155),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1157),
.Y(n_1211)
);

O2A1O1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1177),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_1212)
);

INVxp67_ASAP7_75t_L g1213 ( 
.A(n_1124),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1130),
.Y(n_1214)
);

OAI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1145),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_SL g1216 ( 
.A1(n_1171),
.A2(n_440),
.B(n_439),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1119),
.A2(n_1149),
.B(n_1148),
.C(n_1169),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1131),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1120),
.B(n_40),
.Y(n_1219)
);

AOI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1170),
.A2(n_444),
.B(n_443),
.Y(n_1220)
);

INVx8_ASAP7_75t_L g1221 ( 
.A(n_1129),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1162),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1173),
.A2(n_447),
.B(n_446),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1166),
.B(n_40),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1133),
.A2(n_449),
.B(n_448),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1165),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1146),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1139),
.A2(n_1163),
.B1(n_1141),
.B2(n_1125),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1174),
.A2(n_451),
.B(n_450),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1121),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1135),
.B(n_41),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1159),
.Y(n_1232)
);

BUFx8_ASAP7_75t_L g1233 ( 
.A(n_1147),
.Y(n_1233)
);

OA21x2_ASAP7_75t_L g1234 ( 
.A1(n_1167),
.A2(n_453),
.B(n_452),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1113),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1136),
.B(n_41),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1126),
.A2(n_457),
.B(n_455),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1115),
.A2(n_460),
.B(n_459),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1219),
.A2(n_49),
.B1(n_57),
.B2(n_42),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1192),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1204),
.Y(n_1241)
);

BUFx8_ASAP7_75t_L g1242 ( 
.A(n_1190),
.Y(n_1242)
);

BUFx2_ASAP7_75t_SL g1243 ( 
.A(n_1202),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_1188),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1209),
.Y(n_1245)
);

NAND2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1235),
.B(n_461),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1211),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1201),
.B(n_44),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1196),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1184),
.B(n_462),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1191),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1179),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1224),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1253)
);

OA21x2_ASAP7_75t_L g1254 ( 
.A1(n_1193),
.A2(n_466),
.B(n_463),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1222),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1227),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1226),
.B(n_48),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1231),
.B(n_50),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1218),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1230),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1183),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1186),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1181),
.A2(n_51),
.B(n_52),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1203),
.B(n_51),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1236),
.B(n_53),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1208),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_SL g1267 ( 
.A1(n_1233),
.A2(n_63),
.B1(n_71),
.B2(n_54),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1213),
.B(n_54),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1232),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1198),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1198),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1197),
.B(n_55),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1206),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_1178),
.B(n_467),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1214),
.Y(n_1275)
);

INVx6_ASAP7_75t_L g1276 ( 
.A(n_1205),
.Y(n_1276)
);

AO21x2_ASAP7_75t_L g1277 ( 
.A1(n_1238),
.A2(n_469),
.B(n_468),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1187),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1220),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1185),
.A2(n_59),
.B1(n_56),
.B2(n_58),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1195),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1251),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1244),
.B(n_1182),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_1240),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1266),
.B(n_1221),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_R g1286 ( 
.A(n_1242),
.B(n_1210),
.Y(n_1286)
);

BUFx10_ASAP7_75t_L g1287 ( 
.A(n_1276),
.Y(n_1287)
);

NAND2xp33_ASAP7_75t_R g1288 ( 
.A(n_1250),
.B(n_1234),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_1241),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1278),
.B(n_1256),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1263),
.B(n_1180),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1252),
.B(n_1217),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1258),
.B(n_1199),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1261),
.B(n_1228),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1260),
.B(n_1212),
.Y(n_1295)
);

OR2x6_ASAP7_75t_L g1296 ( 
.A(n_1243),
.B(n_1194),
.Y(n_1296)
);

NAND2xp33_ASAP7_75t_R g1297 ( 
.A(n_1281),
.B(n_1207),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1245),
.Y(n_1298)
);

OR2x4_ASAP7_75t_L g1299 ( 
.A(n_1257),
.B(n_1215),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1264),
.B(n_1189),
.Y(n_1300)
);

XNOR2xp5_ASAP7_75t_L g1301 ( 
.A(n_1265),
.B(n_1200),
.Y(n_1301)
);

NAND2xp33_ASAP7_75t_R g1302 ( 
.A(n_1268),
.B(n_1274),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1287),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1282),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1294),
.B(n_1248),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1298),
.B(n_1255),
.Y(n_1306)
);

AOI222xp33_ASAP7_75t_L g1307 ( 
.A1(n_1291),
.A2(n_1253),
.B1(n_1293),
.B2(n_1272),
.C1(n_1280),
.C2(n_1300),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1301),
.A2(n_1239),
.B1(n_1267),
.B2(n_1277),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1299),
.A2(n_1273),
.B1(n_1249),
.B2(n_1269),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1290),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1283),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1284),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1292),
.B(n_1275),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1289),
.B(n_1247),
.Y(n_1314)
);

OAI22xp33_ASAP7_75t_SL g1315 ( 
.A1(n_1295),
.A2(n_1279),
.B1(n_1271),
.B2(n_1270),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1296),
.B(n_1259),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1286),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1302),
.B(n_1262),
.Y(n_1318)
);

INVx5_ASAP7_75t_L g1319 ( 
.A(n_1297),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1288),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1285),
.B(n_1254),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1303),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1304),
.Y(n_1323)
);

NAND3xp33_ASAP7_75t_L g1324 ( 
.A(n_1307),
.B(n_1216),
.C(n_1246),
.Y(n_1324)
);

INVx5_ASAP7_75t_L g1325 ( 
.A(n_1319),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1308),
.A2(n_1229),
.B1(n_1223),
.B2(n_1225),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1306),
.Y(n_1327)
);

AOI33xp33_ASAP7_75t_L g1328 ( 
.A1(n_1312),
.A2(n_66),
.A3(n_68),
.B1(n_64),
.B2(n_65),
.B3(n_67),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1310),
.B(n_70),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_1314),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1315),
.Y(n_1331)
);

INVxp67_ASAP7_75t_SL g1332 ( 
.A(n_1318),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1316),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1321),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1313),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1305),
.B(n_1237),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1311),
.B(n_73),
.Y(n_1337)
);

AND3x1_ASAP7_75t_L g1338 ( 
.A(n_1317),
.B(n_76),
.C(n_77),
.Y(n_1338)
);

AO21x2_ASAP7_75t_L g1339 ( 
.A1(n_1320),
.A2(n_77),
.B(n_78),
.Y(n_1339)
);

AOI221xp5_ASAP7_75t_L g1340 ( 
.A1(n_1309),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.C(n_82),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1304),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1327),
.B(n_1331),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1341),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1333),
.B(n_1330),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1335),
.B(n_87),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1325),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1336),
.B(n_88),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1325),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1329),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1337),
.B(n_89),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1339),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1328),
.B(n_90),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1324),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1338),
.B(n_91),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1326),
.B(n_92),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1340),
.B(n_94),
.Y(n_1356)
);

INVx4_ASAP7_75t_L g1357 ( 
.A(n_1322),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1332),
.B(n_95),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1323),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1332),
.B(n_98),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1323),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1334),
.B(n_99),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_SL g1363 ( 
.A1(n_1354),
.A2(n_105),
.B1(n_101),
.B2(n_104),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1349),
.B(n_106),
.Y(n_1364)
);

NOR2x1_ASAP7_75t_L g1365 ( 
.A(n_1357),
.B(n_107),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1342),
.Y(n_1366)
);

AO221x2_ASAP7_75t_L g1367 ( 
.A1(n_1351),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.C(n_112),
.Y(n_1367)
);

INVxp67_ASAP7_75t_SL g1368 ( 
.A(n_1346),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1348),
.Y(n_1369)
);

AO221x2_ASAP7_75t_L g1370 ( 
.A1(n_1352),
.A2(n_120),
.B1(n_122),
.B2(n_119),
.C(n_121),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1356),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1343),
.B(n_126),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1355),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1344),
.B(n_136),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1359),
.B(n_138),
.Y(n_1375)
);

OAI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1362),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1361),
.B(n_143),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1347),
.B(n_151),
.Y(n_1378)
);

AO221x2_ASAP7_75t_L g1379 ( 
.A1(n_1358),
.A2(n_155),
.B1(n_152),
.B2(n_153),
.C(n_156),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1360),
.B(n_160),
.Y(n_1380)
);

AO221x2_ASAP7_75t_L g1381 ( 
.A1(n_1350),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.C(n_166),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1345),
.B(n_163),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1342),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1357),
.Y(n_1384)
);

OAI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1353),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_1385)
);

NAND2xp33_ASAP7_75t_R g1386 ( 
.A(n_1354),
.B(n_177),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1384),
.B(n_182),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1374),
.B(n_187),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1372),
.B(n_188),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1375),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1377),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1364),
.B(n_189),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1365),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1378),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1380),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1382),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1379),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1381),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1373),
.B(n_1371),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1376),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1385),
.Y(n_1401)
);

INVxp67_ASAP7_75t_L g1402 ( 
.A(n_1386),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1367),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1366),
.B(n_198),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1384),
.B(n_199),
.Y(n_1405)
);

AOI222xp33_ASAP7_75t_L g1406 ( 
.A1(n_1363),
.A2(n_205),
.B1(n_207),
.B2(n_202),
.C1(n_204),
.C2(n_206),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1369),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1369),
.A2(n_208),
.B(n_209),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1383),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1370),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1369),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1368),
.B(n_214),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1396),
.B(n_214),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1393),
.B(n_215),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1403),
.A2(n_1397),
.B1(n_1398),
.B2(n_1402),
.Y(n_1415)
);

NAND3xp33_ASAP7_75t_L g1416 ( 
.A(n_1406),
.B(n_222),
.C(n_223),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1412),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1395),
.B(n_231),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1407),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1410),
.A2(n_236),
.B1(n_233),
.B2(n_234),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1409),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1399),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_1422)
);

AO22x2_ASAP7_75t_L g1423 ( 
.A1(n_1390),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1391),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1394),
.B(n_249),
.Y(n_1425)
);

INVxp67_ASAP7_75t_L g1426 ( 
.A(n_1400),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1401),
.A2(n_253),
.B1(n_250),
.B2(n_252),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1411),
.B(n_254),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1404),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1387),
.Y(n_1430)
);

CKINVDCx16_ASAP7_75t_R g1431 ( 
.A(n_1415),
.Y(n_1431)
);

INVx2_ASAP7_75t_SL g1432 ( 
.A(n_1417),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1430),
.B(n_1426),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1416),
.A2(n_1389),
.B1(n_1388),
.B2(n_1392),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1429),
.B(n_1405),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1421),
.B(n_1408),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1418),
.B(n_259),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1419),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1425),
.B(n_1428),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1424),
.B(n_262),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1414),
.B(n_264),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1413),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1439),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1431),
.B(n_1432),
.Y(n_1444)
);

CKINVDCx6p67_ASAP7_75t_R g1445 ( 
.A(n_1437),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1438),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1433),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1440),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1436),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1435),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1442),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1434),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1441),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1444),
.Y(n_1454)
);

AOI221xp5_ASAP7_75t_L g1455 ( 
.A1(n_1452),
.A2(n_1422),
.B1(n_1427),
.B2(n_1423),
.C(n_1420),
.Y(n_1455)
);

NAND5xp2_ASAP7_75t_L g1456 ( 
.A(n_1451),
.B(n_270),
.C(n_267),
.D(n_269),
.E(n_271),
.Y(n_1456)
);

NOR3xp33_ASAP7_75t_SL g1457 ( 
.A(n_1447),
.B(n_272),
.C(n_273),
.Y(n_1457)
);

O2A1O1Ixp5_ASAP7_75t_L g1458 ( 
.A1(n_1449),
.A2(n_277),
.B(n_274),
.C(n_275),
.Y(n_1458)
);

NAND4xp25_ASAP7_75t_L g1459 ( 
.A(n_1443),
.B(n_280),
.C(n_278),
.D(n_279),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1445),
.B(n_284),
.Y(n_1460)
);

NAND3xp33_ASAP7_75t_L g1461 ( 
.A(n_1446),
.B(n_291),
.C(n_292),
.Y(n_1461)
);

NAND4xp25_ASAP7_75t_L g1462 ( 
.A(n_1450),
.B(n_294),
.C(n_292),
.D(n_293),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1448),
.B(n_295),
.Y(n_1463)
);

NOR2x1_ASAP7_75t_L g1464 ( 
.A(n_1453),
.B(n_298),
.Y(n_1464)
);

NOR3xp33_ASAP7_75t_L g1465 ( 
.A(n_1454),
.B(n_300),
.C(n_301),
.Y(n_1465)
);

AOI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1455),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.C(n_309),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1457),
.Y(n_1467)
);

AOI21xp33_ASAP7_75t_L g1468 ( 
.A1(n_1460),
.A2(n_316),
.B(n_317),
.Y(n_1468)
);

XOR2xp5_ASAP7_75t_L g1469 ( 
.A(n_1459),
.B(n_319),
.Y(n_1469)
);

NAND4xp25_ASAP7_75t_L g1470 ( 
.A(n_1456),
.B(n_323),
.C(n_320),
.D(n_321),
.Y(n_1470)
);

AO22x1_ASAP7_75t_L g1471 ( 
.A1(n_1464),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_1471)
);

NOR2x1_ASAP7_75t_L g1472 ( 
.A(n_1461),
.B(n_329),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1458),
.B(n_330),
.Y(n_1473)
);

AOI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1462),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.C(n_334),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1463),
.Y(n_1475)
);

XNOR2xp5_ASAP7_75t_L g1476 ( 
.A(n_1469),
.B(n_336),
.Y(n_1476)
);

NAND2x1p5_ASAP7_75t_L g1477 ( 
.A(n_1472),
.B(n_340),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1471),
.B(n_342),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1466),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1470),
.B(n_347),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1467),
.B(n_347),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1473),
.B(n_348),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_R g1483 ( 
.A(n_1476),
.B(n_1475),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_R g1484 ( 
.A(n_1482),
.B(n_1465),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_R g1485 ( 
.A(n_1478),
.B(n_1468),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1484),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1486),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1487),
.A2(n_1477),
.B1(n_1479),
.B2(n_1481),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1488),
.A2(n_1485),
.B1(n_1483),
.B2(n_1480),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1489),
.B(n_1474),
.Y(n_1490)
);

AOI222xp33_ASAP7_75t_L g1491 ( 
.A1(n_1490),
.A2(n_351),
.B1(n_352),
.B2(n_353),
.C1(n_354),
.C2(n_355),
.Y(n_1491)
);

INVxp67_ASAP7_75t_SL g1492 ( 
.A(n_1491),
.Y(n_1492)
);

AOI221xp5_ASAP7_75t_L g1493 ( 
.A1(n_1492),
.A2(n_358),
.B1(n_356),
.B2(n_357),
.C(n_359),
.Y(n_1493)
);

AOI211xp5_ASAP7_75t_L g1494 ( 
.A1(n_1493),
.A2(n_360),
.B(n_357),
.C(n_358),
.Y(n_1494)
);


endmodule