module fake_netlist_6_3104_n_2353 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2353);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2353;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2255;
wire n_2112;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_138),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_14),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_91),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_177),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_190),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_107),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_197),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_82),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_112),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_209),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_80),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_63),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_183),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_49),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_81),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_153),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_152),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_67),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_66),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_172),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_41),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_105),
.Y(n_260)
);

BUFx8_ASAP7_75t_SL g261 ( 
.A(n_223),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_86),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_130),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_65),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_227),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_156),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_229),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_95),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_144),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_191),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_173),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_129),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_103),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_143),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_35),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_125),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_170),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_189),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_121),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_148),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_205),
.Y(n_281)
);

INVxp33_ASAP7_75t_SL g282 ( 
.A(n_149),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_213),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_39),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_184),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_201),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_3),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_117),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_136),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_30),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_222),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_202),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_180),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_237),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_8),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_147),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_41),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_154),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_159),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_176),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_99),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_50),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_18),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_163),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_70),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_139),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_185),
.Y(n_307)
);

BUFx10_ASAP7_75t_L g308 ( 
.A(n_36),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_56),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_13),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_119),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_141),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_31),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_69),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_194),
.Y(n_315)
);

BUFx2_ASAP7_75t_SL g316 ( 
.A(n_1),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_198),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_174),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_65),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_42),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_216),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_76),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_219),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_19),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_45),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_131),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_42),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_124),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_207),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_235),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_203),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_182),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_61),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_66),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_75),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_168),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_97),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_155),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_3),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_76),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_187),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_113),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_192),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_94),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_175),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_218),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_101),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_17),
.Y(n_348)
);

BUFx10_ASAP7_75t_L g349 ( 
.A(n_45),
.Y(n_349)
);

BUFx8_ASAP7_75t_SL g350 ( 
.A(n_208),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_217),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_0),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_14),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_89),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_210),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_225),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_39),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_115),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_79),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_18),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_167),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_110),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_199),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_86),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_61),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_200),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_109),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_106),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_231),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_58),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_123),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_78),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_11),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_162),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_150),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_2),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_80),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_46),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_2),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_74),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_59),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_164),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_29),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_31),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_93),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_22),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_6),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_220),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_10),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_21),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_171),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_59),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_232),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_48),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_51),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_72),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_98),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_55),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_75),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_58),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_46),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_60),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_35),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_27),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_111),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_12),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_166),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_47),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_132),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_4),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_48),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_73),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_146),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_133),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_96),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_62),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_234),
.Y(n_417)
);

BUFx8_ASAP7_75t_SL g418 ( 
.A(n_84),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_52),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_0),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_19),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_23),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_169),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_120),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_211),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_118),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_87),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_90),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_178),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_221),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_60),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_27),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_34),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_85),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_8),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_236),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_204),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_23),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_96),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_15),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_127),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_43),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_212),
.Y(n_443)
);

INVx2_ASAP7_75t_SL g444 ( 
.A(n_32),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_102),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_62),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_47),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_51),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_195),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_26),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_32),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_78),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_10),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_91),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_22),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_81),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_94),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_33),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_186),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_67),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_157),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_104),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_122),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_12),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_93),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_314),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_261),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_314),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_314),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_314),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_350),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_418),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_314),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_422),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_314),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_254),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_411),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_238),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_411),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_271),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_256),
.B(n_1),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_321),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_411),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_411),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_241),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_411),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_411),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_312),
.B(n_4),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_242),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_433),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_433),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_R g492 ( 
.A(n_329),
.B(n_100),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_255),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_433),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_280),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_433),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_293),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_315),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_377),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g500 ( 
.A(n_377),
.B(n_5),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_422),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_433),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_433),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_460),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_321),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_377),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_464),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_282),
.B(n_5),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_464),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_256),
.B(n_6),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_243),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_377),
.Y(n_512)
);

INVxp33_ASAP7_75t_SL g513 ( 
.A(n_399),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_460),
.Y(n_514)
);

BUFx10_ASAP7_75t_L g515 ( 
.A(n_460),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_317),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_460),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_244),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_460),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_247),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_258),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g522 ( 
.A(n_308),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_460),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_260),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_326),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_393),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_386),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_386),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_266),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_386),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_386),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_267),
.B(n_7),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_409),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_327),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_316),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_267),
.B(n_7),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_327),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_239),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_417),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_269),
.Y(n_540)
);

INVxp33_ASAP7_75t_SL g541 ( 
.A(n_248),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_257),
.B(n_9),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_243),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_273),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_274),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_276),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_278),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_279),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_327),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_286),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_289),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_353),
.Y(n_552)
);

CKINVDCx16_ASAP7_75t_R g553 ( 
.A(n_308),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_291),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_316),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_253),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_353),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_294),
.Y(n_558)
);

INVxp67_ASAP7_75t_SL g559 ( 
.A(n_276),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_353),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_264),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_298),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_299),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_240),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_301),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_304),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_257),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_303),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_303),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_322),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_322),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_430),
.B(n_9),
.Y(n_572)
);

BUFx2_ASAP7_75t_SL g573 ( 
.A(n_430),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_311),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_324),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_323),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_331),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_246),
.B(n_11),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_332),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_324),
.Y(n_580)
);

INVxp33_ASAP7_75t_L g581 ( 
.A(n_334),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_334),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_336),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_339),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_339),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_345),
.Y(n_586)
);

INVxp67_ASAP7_75t_SL g587 ( 
.A(n_276),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_344),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_344),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_348),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_346),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_348),
.B(n_13),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_246),
.B(n_15),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_466),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_506),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_507),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_466),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_468),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_468),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_469),
.Y(n_600)
);

AND2x6_ASAP7_75t_L g601 ( 
.A(n_527),
.B(n_250),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_515),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_469),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_556),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_506),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_528),
.B(n_437),
.Y(n_606)
);

BUFx8_ASAP7_75t_L g607 ( 
.A(n_556),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_499),
.B(n_437),
.Y(n_608)
);

OA21x2_ASAP7_75t_L g609 ( 
.A1(n_527),
.A2(n_376),
.B(n_357),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_470),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_549),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_512),
.B(n_437),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_470),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_573),
.B(n_306),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_473),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_473),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_475),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_475),
.Y(n_618)
);

OA21x2_ASAP7_75t_L g619 ( 
.A1(n_530),
.A2(n_376),
.B(n_357),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_528),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_549),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_SL g622 ( 
.A1(n_509),
.A2(n_297),
.B1(n_333),
.B2(n_259),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_477),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_477),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_479),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_546),
.B(n_351),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_573),
.B(n_330),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_559),
.B(n_250),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_587),
.B(n_355),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_530),
.B(n_250),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_479),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_536),
.B(n_356),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_538),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_572),
.B(n_361),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_515),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_483),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_483),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_484),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_476),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_484),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_486),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_486),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_561),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_487),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_487),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_490),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_490),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_491),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_491),
.Y(n_649)
);

NOR2x1_ASAP7_75t_L g650 ( 
.A(n_532),
.B(n_288),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_494),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_494),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_531),
.B(n_288),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_496),
.Y(n_654)
);

AND2x6_ASAP7_75t_L g655 ( 
.A(n_531),
.B(n_288),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_496),
.Y(n_656)
);

AND2x6_ASAP7_75t_L g657 ( 
.A(n_502),
.B(n_300),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_500),
.B(n_300),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_513),
.B(n_445),
.Y(n_659)
);

INVxp33_ASAP7_75t_L g660 ( 
.A(n_474),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_502),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_503),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_511),
.B(n_300),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_488),
.B(n_382),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_547),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_503),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_504),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_504),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_514),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_514),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_517),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_543),
.B(n_443),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_517),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_519),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_519),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_523),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_523),
.B(n_443),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_534),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_515),
.Y(n_679)
);

OAI21x1_ASAP7_75t_L g680 ( 
.A1(n_481),
.A2(n_443),
.B(n_263),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_534),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_567),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_537),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_567),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_548),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_537),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_568),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_568),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_569),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_552),
.B(n_251),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_552),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_557),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_609),
.Y(n_693)
);

INVxp67_ASAP7_75t_SL g694 ( 
.A(n_680),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_609),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_595),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_609),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_SL g698 ( 
.A(n_664),
.B(n_245),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_664),
.B(n_541),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_659),
.B(n_482),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_598),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_595),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_598),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_626),
.B(n_478),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_609),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_598),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_659),
.B(n_505),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_596),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_626),
.B(n_485),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_609),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_L g711 ( 
.A1(n_596),
.A2(n_480),
.B1(n_249),
.B2(n_245),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_629),
.B(n_489),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_629),
.B(n_518),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_606),
.B(n_251),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_632),
.B(n_520),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_614),
.B(n_521),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_632),
.B(n_524),
.Y(n_717)
);

OR2x6_ASAP7_75t_L g718 ( 
.A(n_680),
.B(n_481),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_609),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_619),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_634),
.B(n_529),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_634),
.B(n_540),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_614),
.B(n_544),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_604),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_627),
.B(n_545),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_650),
.A2(n_578),
.B1(n_593),
.B2(n_501),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_598),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_608),
.B(n_550),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_650),
.A2(n_508),
.B1(n_542),
.B2(n_510),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_608),
.B(n_551),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_619),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_600),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_L g733 ( 
.A1(n_660),
.A2(n_249),
.B1(n_455),
.B2(n_262),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_619),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_600),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_639),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_619),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_600),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_L g739 ( 
.A(n_608),
.B(n_492),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_600),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_610),
.Y(n_741)
);

INVxp67_ASAP7_75t_SL g742 ( 
.A(n_680),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_610),
.Y(n_743)
);

INVx4_ASAP7_75t_L g744 ( 
.A(n_595),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_602),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_658),
.A2(n_542),
.B1(n_592),
.B2(n_510),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_595),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_628),
.B(n_554),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_628),
.B(n_558),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_612),
.B(n_562),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_595),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_612),
.B(n_566),
.Y(n_752)
);

INVx4_ASAP7_75t_L g753 ( 
.A(n_595),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_619),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_612),
.B(n_574),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_628),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_658),
.A2(n_592),
.B1(n_444),
.B2(n_268),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_658),
.A2(n_444),
.B1(n_268),
.B2(n_379),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_610),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_619),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_658),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_633),
.B(n_576),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_602),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_610),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_602),
.Y(n_765)
);

OAI22xp33_ASAP7_75t_L g766 ( 
.A1(n_660),
.A2(n_553),
.B1(n_522),
.B2(n_581),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_633),
.B(n_577),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_623),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_602),
.B(n_579),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_597),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_623),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_633),
.B(n_583),
.Y(n_772)
);

OAI22xp33_ASAP7_75t_L g773 ( 
.A1(n_643),
.A2(n_275),
.B1(n_287),
.B2(n_284),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_597),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_643),
.B(n_586),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_663),
.B(n_557),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_639),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_606),
.B(n_263),
.Y(n_778)
);

NAND2x1p5_ASAP7_75t_L g779 ( 
.A(n_658),
.B(n_270),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_635),
.B(n_414),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_622),
.A2(n_370),
.B1(n_401),
.B2(n_380),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_595),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_643),
.B(n_591),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_599),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_599),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_603),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_635),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_623),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_623),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_624),
.Y(n_790)
);

AND3x1_ASAP7_75t_L g791 ( 
.A(n_663),
.B(n_379),
.C(n_378),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_603),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_663),
.B(n_560),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_616),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_635),
.B(n_362),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_624),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_616),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_607),
.B(n_563),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_658),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_635),
.B(n_363),
.Y(n_800)
);

INVxp67_ASAP7_75t_SL g801 ( 
.A(n_679),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_595),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_690),
.A2(n_402),
.B1(n_406),
.B2(n_378),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_605),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_SL g805 ( 
.A1(n_607),
.A2(n_416),
.B1(n_564),
.B2(n_495),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_672),
.B(n_560),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_617),
.Y(n_807)
);

INVx5_ASAP7_75t_L g808 ( 
.A(n_657),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_617),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_604),
.B(n_565),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_624),
.Y(n_811)
);

AND2x6_ASAP7_75t_L g812 ( 
.A(n_630),
.B(n_283),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_618),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_622),
.B(n_252),
.C(n_535),
.Y(n_814)
);

OAI22xp33_ASAP7_75t_L g815 ( 
.A1(n_604),
.A2(n_295),
.B1(n_302),
.B2(n_290),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_679),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_618),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_606),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_624),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_679),
.B(n_467),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_605),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_606),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_625),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_607),
.B(n_471),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_638),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_679),
.B(n_366),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_625),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_605),
.Y(n_828)
);

INVx4_ASAP7_75t_L g829 ( 
.A(n_605),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_638),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_638),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_690),
.A2(n_406),
.B1(n_410),
.B2(n_402),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_644),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_682),
.B(n_555),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_606),
.B(n_270),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_690),
.A2(n_415),
.B1(n_420),
.B2(n_410),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_605),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_638),
.Y(n_838)
);

OR2x6_ASAP7_75t_L g839 ( 
.A(n_606),
.B(n_272),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_607),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_644),
.B(n_367),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_649),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_649),
.Y(n_843)
);

OR2x6_ASAP7_75t_L g844 ( 
.A(n_630),
.B(n_272),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_649),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_649),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_682),
.B(n_472),
.Y(n_847)
);

INVxp33_ASAP7_75t_L g848 ( 
.A(n_672),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_645),
.B(n_368),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_652),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_645),
.B(n_369),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_630),
.Y(n_852)
);

BUFx3_ASAP7_75t_L g853 ( 
.A(n_690),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_647),
.B(n_371),
.Y(n_854)
);

INVx5_ASAP7_75t_L g855 ( 
.A(n_657),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_738),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_715),
.B(n_653),
.Y(n_857)
);

NOR2x1_ASAP7_75t_L g858 ( 
.A(n_820),
.B(n_493),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_756),
.B(n_653),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_699),
.A2(n_498),
.B1(n_516),
.B2(n_497),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_738),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_728),
.A2(n_526),
.B1(n_533),
.B2(n_525),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_776),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_708),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_698),
.B(n_607),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_695),
.A2(n_653),
.B1(n_690),
.B2(n_420),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_756),
.B(n_690),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_738),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_708),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_852),
.B(n_684),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_852),
.B(n_672),
.Y(n_871)
);

AND2x6_ASAP7_75t_SL g872 ( 
.A(n_810),
.B(n_415),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_704),
.B(n_647),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_698),
.A2(n_442),
.B(n_446),
.C(n_431),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_776),
.B(n_684),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_761),
.B(n_651),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_740),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_761),
.A2(n_677),
.B(n_662),
.Y(n_878)
);

OAI221xp5_ASAP7_75t_L g879 ( 
.A1(n_729),
.A2(n_746),
.B1(n_726),
.B2(n_757),
.C(n_758),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_748),
.B(n_607),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_793),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_799),
.B(n_717),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_740),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_799),
.B(n_651),
.Y(n_884)
);

INVx8_ASAP7_75t_L g885 ( 
.A(n_718),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_793),
.B(n_687),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_693),
.B(n_283),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_749),
.B(n_320),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_806),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_SL g890 ( 
.A(n_840),
.B(n_665),
.Y(n_890)
);

OAI221xp5_ASAP7_75t_L g891 ( 
.A1(n_803),
.A2(n_373),
.B1(n_590),
.B2(n_580),
.C(n_456),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_730),
.A2(n_539),
.B1(n_375),
.B2(n_388),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_721),
.B(n_662),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_750),
.A2(n_391),
.B1(n_397),
.B2(n_374),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_806),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_714),
.B(n_687),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_722),
.B(n_668),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_740),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_752),
.B(n_668),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_736),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_755),
.B(n_670),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_693),
.B(n_283),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_818),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_695),
.A2(n_442),
.B(n_446),
.C(n_431),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_853),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_775),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_777),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_848),
.B(n_305),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_739),
.A2(n_712),
.B1(n_713),
.B2(n_709),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_716),
.B(n_309),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_693),
.B(n_283),
.Y(n_911)
);

INVxp33_ASAP7_75t_L g912 ( 
.A(n_783),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_741),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_693),
.B(n_671),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_818),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_822),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_697),
.A2(n_456),
.B(n_448),
.C(n_277),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_697),
.A2(n_448),
.B(n_277),
.C(n_285),
.Y(n_918)
);

NAND3xp33_ASAP7_75t_L g919 ( 
.A(n_814),
.B(n_313),
.C(n_310),
.Y(n_919)
);

NOR3xp33_ASAP7_75t_L g920 ( 
.A(n_700),
.B(n_685),
.C(n_665),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_741),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_822),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_724),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_743),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_718),
.A2(n_407),
.B1(n_413),
.B2(n_405),
.Y(n_925)
);

INVx8_ASAP7_75t_L g926 ( 
.A(n_718),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_693),
.B(n_671),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_723),
.B(n_319),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_720),
.B(n_675),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_720),
.B(n_675),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_725),
.B(n_325),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_720),
.B(n_676),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_743),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_743),
.Y(n_934)
);

INVxp67_ASAP7_75t_SL g935 ( 
.A(n_720),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_853),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_720),
.B(n_676),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_724),
.B(n_685),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_811),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_853),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_760),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_760),
.B(n_677),
.Y(n_942)
);

OAI21xp33_ASAP7_75t_L g943 ( 
.A1(n_834),
.A2(n_570),
.B(n_569),
.Y(n_943)
);

NAND2xp33_ASAP7_75t_L g944 ( 
.A(n_760),
.B(n_423),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_760),
.B(n_705),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_847),
.B(n_688),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_705),
.A2(n_689),
.B(n_688),
.C(n_613),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_760),
.B(n_677),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_707),
.B(n_335),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_710),
.B(n_677),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_762),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_815),
.B(n_340),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_770),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_710),
.B(n_677),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_770),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_719),
.B(n_283),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_719),
.B(n_677),
.Y(n_957)
);

AND2x6_ASAP7_75t_L g958 ( 
.A(n_731),
.B(n_281),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_811),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_811),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_774),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_731),
.B(n_594),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_769),
.B(n_352),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_714),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_773),
.B(n_767),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_734),
.B(n_594),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_734),
.B(n_594),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_774),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_718),
.A2(n_424),
.B1(n_425),
.B2(n_429),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_772),
.B(n_354),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_784),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_780),
.B(n_359),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_714),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_784),
.Y(n_974)
);

XOR2xp5_ASAP7_75t_L g975 ( 
.A(n_805),
.B(n_436),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_737),
.B(n_283),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_714),
.B(n_689),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_785),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_819),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_737),
.B(n_459),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_785),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_841),
.B(n_360),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_754),
.A2(n_347),
.B(n_281),
.C(n_285),
.Y(n_983)
);

AND2x6_ASAP7_75t_SL g984 ( 
.A(n_781),
.B(n_570),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_754),
.B(n_459),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_786),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_786),
.B(n_613),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_766),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_718),
.A2(n_347),
.B1(n_296),
.B2(n_307),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_792),
.B(n_613),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_792),
.B(n_615),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_694),
.A2(n_742),
.B(n_801),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_844),
.A2(n_463),
.B1(n_449),
.B2(n_461),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_779),
.B(n_459),
.Y(n_994)
);

AND2x4_ASAP7_75t_SL g995 ( 
.A(n_844),
.B(n_265),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_794),
.B(n_797),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_794),
.B(n_615),
.Y(n_997)
);

AO221x1_ASAP7_75t_L g998 ( 
.A1(n_711),
.A2(n_733),
.B1(n_840),
.B2(n_459),
.C(n_343),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_819),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_797),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_807),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_778),
.B(n_571),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_779),
.B(n_459),
.Y(n_1003)
);

NOR2xp67_ASAP7_75t_SL g1004 ( 
.A(n_745),
.B(n_459),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_807),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_809),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_779),
.B(n_605),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_809),
.B(n_615),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_849),
.B(n_364),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_781),
.A2(n_338),
.B(n_296),
.C(n_307),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_844),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_844),
.A2(n_341),
.B1(n_292),
.B2(n_318),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_819),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_813),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_813),
.B(n_631),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_817),
.B(n_823),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_778),
.B(n_605),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_851),
.B(n_365),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_817),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_701),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_823),
.B(n_631),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_844),
.B(n_778),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_854),
.B(n_372),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_827),
.B(n_631),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_827),
.B(n_381),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_824),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_701),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_857),
.B(n_816),
.Y(n_1028)
);

AO21x1_ASAP7_75t_L g1029 ( 
.A1(n_989),
.A2(n_835),
.B(n_778),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_945),
.A2(n_800),
.B(n_795),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_942),
.A2(n_826),
.B(n_839),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_863),
.B(n_798),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_909),
.A2(n_835),
.B1(n_839),
.B2(n_791),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_948),
.A2(n_839),
.B(n_835),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_881),
.B(n_791),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_SL g1036 ( 
.A1(n_983),
.A2(n_292),
.B(n_328),
.C(n_318),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_864),
.B(n_835),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_887),
.A2(n_833),
.B(n_706),
.Y(n_1038)
);

NOR3xp33_ASAP7_75t_L g1039 ( 
.A(n_965),
.B(n_337),
.C(n_328),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_935),
.A2(n_839),
.B(n_763),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_887),
.A2(n_839),
.B(n_763),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_953),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_906),
.B(n_745),
.Y(n_1043)
);

AND2x6_ASAP7_75t_L g1044 ( 
.A(n_941),
.B(n_745),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_965),
.A2(n_833),
.B(n_765),
.C(n_787),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_873),
.B(n_763),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_902),
.A2(n_787),
.B(n_765),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_902),
.A2(n_911),
.B(n_914),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_905),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_936),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_869),
.B(n_787),
.Y(n_1051)
);

AO21x1_ASAP7_75t_L g1052 ( 
.A1(n_865),
.A2(n_880),
.B(n_956),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_940),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_911),
.A2(n_751),
.B(n_744),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_946),
.B(n_832),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_882),
.A2(n_751),
.B(n_744),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_905),
.Y(n_1057)
);

OAI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_879),
.A2(n_337),
.B1(n_341),
.B2(n_338),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_927),
.A2(n_751),
.B(n_744),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_893),
.B(n_836),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_929),
.A2(n_751),
.B(n_744),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_875),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_923),
.B(n_951),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_930),
.A2(n_802),
.B(n_753),
.Y(n_1064)
);

AOI21x1_ASAP7_75t_L g1065 ( 
.A1(n_956),
.A2(n_706),
.B(n_703),
.Y(n_1065)
);

BUFx8_ASAP7_75t_L g1066 ( 
.A(n_938),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_932),
.A2(n_802),
.B(n_753),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_875),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_937),
.A2(n_802),
.B(n_753),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_950),
.A2(n_802),
.B(n_753),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_880),
.A2(n_866),
.B1(n_865),
.B2(n_1022),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_888),
.B(n_308),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_912),
.B(n_383),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_888),
.A2(n_462),
.B(n_441),
.C(n_426),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_992),
.A2(n_829),
.B(n_702),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_L g1076 ( 
.A(n_970),
.B(n_343),
.C(n_342),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_897),
.B(n_696),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_886),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_899),
.B(n_696),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_908),
.Y(n_1080)
);

INVx2_ASAP7_75t_SL g1081 ( 
.A(n_886),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_954),
.A2(n_829),
.B(n_702),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_901),
.B(n_696),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_957),
.A2(n_829),
.B(n_702),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_998),
.A2(n_812),
.B1(n_426),
.B2(n_358),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_871),
.B(n_696),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_988),
.B(n_384),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_963),
.A2(n_812),
.B1(n_782),
.B2(n_837),
.Y(n_1088)
);

O2A1O1Ixp5_ASAP7_75t_L g1089 ( 
.A1(n_976),
.A2(n_702),
.B(n_747),
.C(n_782),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_866),
.A2(n_342),
.B1(n_441),
.B2(n_358),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_870),
.B(n_747),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_963),
.B(n_385),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_870),
.B(n_972),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_867),
.A2(n_829),
.B(n_782),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_972),
.B(n_747),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_859),
.B(n_747),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_982),
.B(n_782),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_982),
.B(n_828),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1009),
.B(n_828),
.Y(n_1099)
);

NOR3xp33_ASAP7_75t_L g1100 ( 
.A(n_970),
.B(n_462),
.C(n_389),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_955),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_908),
.B(n_308),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_976),
.A2(n_837),
.B(n_828),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1009),
.B(n_828),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_905),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_900),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_980),
.A2(n_837),
.B(n_727),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_980),
.A2(n_837),
.B(n_727),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_910),
.A2(n_703),
.B(n_850),
.C(n_846),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_961),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1018),
.B(n_732),
.Y(n_1111)
);

INVx4_ASAP7_75t_L g1112 ( 
.A(n_905),
.Y(n_1112)
);

INVx1_ASAP7_75t_SL g1113 ( 
.A(n_907),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_949),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_L g1115 ( 
.A(n_952),
.B(n_390),
.C(n_387),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_985),
.A2(n_735),
.B(n_732),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_952),
.A2(n_812),
.B1(n_601),
.B2(n_655),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_910),
.A2(n_931),
.B(n_928),
.C(n_1018),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_885),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_1023),
.B(n_804),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_889),
.B(n_349),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_968),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_985),
.A2(n_764),
.B(n_759),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_971),
.B(n_759),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_895),
.B(n_571),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_856),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1007),
.A2(n_768),
.B(n_764),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1007),
.A2(n_771),
.B(n_768),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_928),
.A2(n_825),
.B(n_850),
.C(n_846),
.Y(n_1129)
);

OR2x6_ASAP7_75t_L g1130 ( 
.A(n_885),
.B(n_575),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_941),
.A2(n_804),
.B1(n_821),
.B2(n_843),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_861),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_974),
.B(n_771),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_1002),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_931),
.B(n_804),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_896),
.Y(n_1136)
);

OR2x2_ASAP7_75t_L g1137 ( 
.A(n_860),
.B(n_575),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1017),
.A2(n_789),
.B(n_788),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1017),
.A2(n_789),
.B(n_788),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_978),
.B(n_790),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_862),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_981),
.B(n_790),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_896),
.B(n_804),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_892),
.B(n_392),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_986),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_973),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_962),
.A2(n_825),
.B(n_796),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_878),
.A2(n_830),
.B(n_796),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_944),
.A2(n_831),
.B(n_830),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_966),
.A2(n_967),
.B(n_884),
.Y(n_1150)
);

AO21x1_ASAP7_75t_L g1151 ( 
.A1(n_994),
.A2(n_838),
.B(n_831),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_947),
.A2(n_842),
.B(n_838),
.Y(n_1152)
);

OAI321xp33_ASAP7_75t_L g1153 ( 
.A1(n_1010),
.A2(n_588),
.A3(n_585),
.B1(n_584),
.B2(n_582),
.C(n_589),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_949),
.A2(n_845),
.B(n_843),
.C(n_842),
.Y(n_1154)
);

AOI21xp33_ASAP7_75t_L g1155 ( 
.A1(n_925),
.A2(n_395),
.B(n_394),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_919),
.B(n_396),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1000),
.B(n_845),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_996),
.A2(n_812),
.B(n_637),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1001),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_876),
.A2(n_821),
.B(n_804),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_868),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_994),
.A2(n_821),
.B(n_808),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1005),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1006),
.B(n_812),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_977),
.B(n_890),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_885),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1010),
.A2(n_641),
.B(n_636),
.C(n_637),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1011),
.A2(n_821),
.B1(n_404),
.B2(n_408),
.Y(n_1168)
);

NAND3xp33_ASAP7_75t_L g1169 ( 
.A(n_894),
.B(n_400),
.C(n_398),
.Y(n_1169)
);

OAI21xp33_ASAP7_75t_L g1170 ( 
.A1(n_1025),
.A2(n_412),
.B(n_403),
.Y(n_1170)
);

INVx5_ASAP7_75t_L g1171 ( 
.A(n_926),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_926),
.Y(n_1172)
);

NOR2xp67_ASAP7_75t_L g1173 ( 
.A(n_969),
.B(n_582),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1003),
.A2(n_821),
.B(n_808),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1014),
.B(n_812),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1011),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_926),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_977),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1019),
.B(n_812),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1026),
.B(n_265),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_975),
.B(n_419),
.Y(n_1181)
);

AOI21x1_ASAP7_75t_L g1182 ( 
.A1(n_987),
.A2(n_991),
.B(n_990),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_858),
.B(n_421),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_964),
.B(n_584),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1003),
.A2(n_855),
.B(n_808),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1025),
.B(n_265),
.Y(n_1186)
);

AO21x1_ASAP7_75t_L g1187 ( 
.A1(n_1016),
.A2(n_637),
.B(n_636),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_903),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_958),
.A2(n_640),
.B(n_641),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_958),
.A2(n_640),
.B(n_641),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_904),
.A2(n_917),
.B(n_874),
.C(n_918),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_915),
.A2(n_922),
.B1(n_916),
.B2(n_1012),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_995),
.A2(n_993),
.B(n_1024),
.C(n_1021),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_997),
.A2(n_855),
.B(n_808),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_920),
.B(n_349),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1008),
.A2(n_1015),
.B1(n_983),
.B2(n_1020),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_874),
.B(n_585),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_877),
.Y(n_1198)
);

BUFx8_ASAP7_75t_L g1199 ( 
.A(n_958),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_943),
.B(n_349),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_904),
.A2(n_636),
.B(n_640),
.C(n_674),
.Y(n_1201)
);

AOI21x1_ASAP7_75t_L g1202 ( 
.A1(n_883),
.A2(n_656),
.B(n_667),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1027),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_984),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_898),
.B(n_265),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_958),
.B(n_642),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_913),
.A2(n_855),
.B(n_808),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_958),
.B(n_642),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_921),
.A2(n_855),
.B(n_808),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_924),
.B(n_642),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_917),
.B(n_349),
.Y(n_1211)
);

INVx4_ASAP7_75t_L g1212 ( 
.A(n_933),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_934),
.B(n_642),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_939),
.B(n_855),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_959),
.B(n_642),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_960),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_979),
.B(n_855),
.Y(n_1217)
);

AOI21x1_ASAP7_75t_L g1218 ( 
.A1(n_999),
.A2(n_656),
.B(n_652),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1080),
.B(n_872),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1118),
.A2(n_918),
.B1(n_1013),
.B2(n_891),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1042),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_1106),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1114),
.B(n_427),
.Y(n_1223)
);

INVx4_ASAP7_75t_L g1224 ( 
.A(n_1057),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1066),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1071),
.A2(n_428),
.B1(n_440),
.B2(n_447),
.Y(n_1226)
);

INVx4_ASAP7_75t_L g1227 ( 
.A(n_1057),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1216),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1057),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1058),
.A2(n_681),
.B(n_692),
.C(n_691),
.Y(n_1230)
);

NOR4xp25_ASAP7_75t_SL g1231 ( 
.A(n_1186),
.B(n_452),
.C(n_434),
.D(n_435),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1093),
.B(n_432),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1072),
.B(n_588),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1063),
.B(n_589),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1092),
.B(n_438),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_SL g1236 ( 
.A(n_1113),
.B(n_1066),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1150),
.A2(n_605),
.B(n_620),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_1141),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1087),
.B(n_439),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1101),
.Y(n_1240)
);

NOR3xp33_ASAP7_75t_SL g1241 ( 
.A(n_1181),
.B(n_450),
.C(n_451),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1110),
.Y(n_1242)
);

NAND2xp33_ASAP7_75t_L g1243 ( 
.A(n_1044),
.B(n_601),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1172),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1028),
.B(n_1004),
.Y(n_1245)
);

NAND2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1171),
.B(n_620),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1150),
.A2(n_1048),
.B(n_1097),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1122),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1145),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1137),
.B(n_453),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1159),
.Y(n_1251)
);

AO32x1_ASAP7_75t_L g1252 ( 
.A1(n_1090),
.A2(n_1196),
.A3(n_1192),
.B1(n_1211),
.B2(n_1102),
.Y(n_1252)
);

INVx2_ASAP7_75t_SL g1253 ( 
.A(n_1176),
.Y(n_1253)
);

INVx4_ASAP7_75t_L g1254 ( 
.A(n_1172),
.Y(n_1254)
);

OR2x6_ASAP7_75t_L g1255 ( 
.A(n_1130),
.B(n_1119),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1048),
.A2(n_620),
.B(n_621),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1144),
.A2(n_681),
.B1(n_655),
.B2(n_601),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1032),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1098),
.A2(n_620),
.B(n_621),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1172),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1163),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1184),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1184),
.Y(n_1263)
);

O2A1O1Ixp33_ASAP7_75t_SL g1264 ( 
.A1(n_1045),
.A2(n_674),
.B(n_648),
.C(n_669),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1177),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1124),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1073),
.B(n_1183),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1100),
.A2(n_454),
.B(n_457),
.C(n_458),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1046),
.B(n_648),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1099),
.A2(n_1104),
.B(n_1031),
.Y(n_1270)
);

INVxp33_ASAP7_75t_SL g1271 ( 
.A(n_1204),
.Y(n_1271)
);

INVx3_ASAP7_75t_SL g1272 ( 
.A(n_1130),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1055),
.B(n_648),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1032),
.B(n_465),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1125),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1037),
.B(n_692),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1170),
.B(n_16),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1133),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1060),
.B(n_648),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1188),
.B(n_648),
.Y(n_1280)
);

AOI33xp33_ASAP7_75t_L g1281 ( 
.A1(n_1125),
.A2(n_1121),
.A3(n_1195),
.B1(n_1035),
.B2(n_1200),
.B3(n_1197),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1079),
.B(n_654),
.Y(n_1282)
);

NOR2x1_ASAP7_75t_L g1283 ( 
.A(n_1119),
.B(n_654),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1083),
.B(n_654),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1039),
.B(n_654),
.Y(n_1285)
);

INVx5_ASAP7_75t_L g1286 ( 
.A(n_1044),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1216),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1062),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_SL g1289 ( 
.A1(n_1115),
.A2(n_1081),
.B1(n_1130),
.B2(n_1156),
.Y(n_1289)
);

NOR2x1_ASAP7_75t_L g1290 ( 
.A(n_1166),
.B(n_654),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1177),
.Y(n_1291)
);

BUFx4f_ASAP7_75t_L g1292 ( 
.A(n_1177),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1076),
.B(n_1155),
.C(n_1169),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1035),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1146),
.B(n_620),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1126),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1140),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1146),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1031),
.A2(n_620),
.B(n_611),
.Y(n_1299)
);

INVx4_ASAP7_75t_L g1300 ( 
.A(n_1171),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1068),
.Y(n_1301)
);

INVx5_ASAP7_75t_L g1302 ( 
.A(n_1044),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1132),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1193),
.A2(n_620),
.B1(n_669),
.B2(n_674),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1078),
.B(n_108),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1033),
.A2(n_620),
.B1(n_669),
.B2(n_674),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1165),
.A2(n_601),
.B1(n_655),
.B2(n_657),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1111),
.A2(n_669),
.B1(n_673),
.B2(n_674),
.Y(n_1308)
);

OR2x6_ASAP7_75t_L g1309 ( 
.A(n_1166),
.B(n_1136),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1077),
.B(n_669),
.Y(n_1310)
);

AO22x1_ASAP7_75t_L g1311 ( 
.A1(n_1199),
.A2(n_655),
.B1(n_601),
.B2(n_657),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1051),
.B(n_16),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1041),
.A2(n_673),
.B1(n_652),
.B2(n_667),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1034),
.A2(n_673),
.B(n_652),
.Y(n_1314)
);

AOI221xp5_ASAP7_75t_L g1315 ( 
.A1(n_1074),
.A2(n_692),
.B1(n_691),
.B2(n_683),
.C(n_678),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1171),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1095),
.A2(n_621),
.B(n_611),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1134),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1142),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1161),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1112),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1049),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1180),
.B(n_17),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1191),
.A2(n_692),
.B(n_691),
.C(n_683),
.Y(n_1324)
);

O2A1O1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1167),
.A2(n_691),
.B(n_683),
.C(n_678),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1036),
.A2(n_683),
.B(n_678),
.C(n_656),
.Y(n_1326)
);

NAND3xp33_ASAP7_75t_SL g1327 ( 
.A(n_1052),
.B(n_667),
.C(n_656),
.Y(n_1327)
);

AOI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1120),
.A2(n_1135),
.B(n_1040),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1043),
.B(n_20),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1049),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1030),
.A2(n_621),
.B(n_611),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1178),
.B(n_114),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1198),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1157),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1203),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1050),
.Y(n_1336)
);

NOR3xp33_ASAP7_75t_SL g1337 ( 
.A(n_1168),
.B(n_20),
.C(n_21),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1053),
.Y(n_1338)
);

O2A1O1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1153),
.A2(n_1201),
.B(n_1154),
.C(n_1109),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1212),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1112),
.Y(n_1341)
);

AOI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1040),
.A2(n_667),
.B(n_666),
.Y(n_1342)
);

O2A1O1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1129),
.A2(n_673),
.B(n_621),
.C(n_611),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1091),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1030),
.A2(n_611),
.B(n_666),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1173),
.A2(n_655),
.B1(n_601),
.B2(n_657),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1171),
.B(n_686),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1034),
.A2(n_666),
.B(n_661),
.Y(n_1348)
);

OAI21xp33_ASAP7_75t_L g1349 ( 
.A1(n_1197),
.A2(n_686),
.B(n_666),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1105),
.B(n_116),
.Y(n_1350)
);

AO21x2_ASAP7_75t_L g1351 ( 
.A1(n_1187),
.A2(n_601),
.B(n_655),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1105),
.Y(n_1352)
);

AOI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1047),
.A2(n_666),
.B(n_661),
.Y(n_1353)
);

OAI21xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1158),
.A2(n_24),
.B(n_25),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1212),
.B(n_24),
.Y(n_1355)
);

O2A1O1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1086),
.A2(n_655),
.B(n_601),
.C(n_28),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1041),
.A2(n_666),
.B(n_661),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1056),
.A2(n_1075),
.B(n_1061),
.Y(n_1358)
);

O2A1O1Ixp5_ASAP7_75t_L g1359 ( 
.A1(n_1029),
.A2(n_655),
.B(n_601),
.C(n_657),
.Y(n_1359)
);

NAND3xp33_ASAP7_75t_SL g1360 ( 
.A(n_1205),
.B(n_25),
.C(n_26),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1210),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1182),
.B(n_28),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1199),
.B(n_1047),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_R g1364 ( 
.A(n_1065),
.B(n_126),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1075),
.A2(n_666),
.B(n_661),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1096),
.B(n_601),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1088),
.A2(n_686),
.B1(n_666),
.B2(n_661),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1143),
.B(n_29),
.Y(n_1368)
);

INVx2_ASAP7_75t_SL g1369 ( 
.A(n_1214),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1164),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1044),
.B(n_601),
.Y(n_1371)
);

BUFx8_ASAP7_75t_L g1372 ( 
.A(n_1044),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1213),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1215),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1085),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1147),
.B(n_655),
.Y(n_1376)
);

A2O1A1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1089),
.A2(n_686),
.B(n_661),
.C(n_646),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1059),
.A2(n_661),
.B(n_646),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1148),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1189),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1175),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1117),
.B(n_30),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1324),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1342),
.A2(n_1149),
.B(n_1127),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1324),
.Y(n_1385)
);

BUFx10_ASAP7_75t_L g1386 ( 
.A(n_1219),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1267),
.A2(n_1235),
.B(n_1239),
.C(n_1293),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1294),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1270),
.A2(n_1064),
.B(n_1067),
.Y(n_1389)
);

AO32x2_ASAP7_75t_L g1390 ( 
.A1(n_1220),
.A2(n_1131),
.A3(n_1151),
.B1(n_1152),
.B2(n_1038),
.Y(n_1390)
);

A2O1A1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1281),
.A2(n_1179),
.B(n_1190),
.C(n_1160),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1238),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1221),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1234),
.B(n_1160),
.Y(n_1394)
);

AOI21x1_ASAP7_75t_SL g1395 ( 
.A1(n_1245),
.A2(n_1208),
.B(n_1206),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_SL g1396 ( 
.A1(n_1339),
.A2(n_1054),
.B(n_1094),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1240),
.Y(n_1397)
);

AO31x2_ASAP7_75t_L g1398 ( 
.A1(n_1270),
.A2(n_1149),
.A3(n_1094),
.B(n_1054),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1242),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1247),
.A2(n_1069),
.B(n_1070),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1248),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1247),
.A2(n_1084),
.B(n_1082),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1380),
.A2(n_1084),
.B(n_1138),
.Y(n_1403)
);

NAND2x1p5_ASAP7_75t_L g1404 ( 
.A(n_1292),
.B(n_1217),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1249),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1251),
.Y(n_1406)
);

AO31x2_ASAP7_75t_L g1407 ( 
.A1(n_1358),
.A2(n_1127),
.A3(n_1128),
.B(n_1123),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1261),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1365),
.A2(n_1128),
.B(n_1123),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1222),
.Y(n_1410)
);

NAND2xp33_ASAP7_75t_SL g1411 ( 
.A(n_1265),
.B(n_1254),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1233),
.B(n_1138),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1358),
.A2(n_1103),
.B(n_1108),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1266),
.B(n_1139),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1285),
.A2(n_1139),
.B(n_1103),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1379),
.A2(n_1116),
.B(n_1107),
.Y(n_1416)
);

AO31x2_ASAP7_75t_L g1417 ( 
.A1(n_1377),
.A2(n_1116),
.A3(n_1108),
.B(n_1107),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1292),
.Y(n_1418)
);

A2O1A1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1277),
.A2(n_1194),
.B(n_1162),
.C(n_1174),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1271),
.Y(n_1420)
);

INVx5_ASAP7_75t_L g1421 ( 
.A(n_1316),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1223),
.B(n_1162),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1375),
.A2(n_1174),
.B1(n_1194),
.B2(n_1209),
.Y(n_1423)
);

OA22x2_ASAP7_75t_L g1424 ( 
.A1(n_1253),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1258),
.B(n_1202),
.Y(n_1425)
);

AO31x2_ASAP7_75t_L g1426 ( 
.A1(n_1362),
.A2(n_1209),
.A3(n_1185),
.B(n_1207),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1286),
.A2(n_1185),
.B(n_686),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1323),
.A2(n_686),
.B(n_1218),
.C(n_661),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1289),
.A2(n_655),
.B1(n_657),
.B2(n_686),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1365),
.A2(n_657),
.B(n_181),
.Y(n_1430)
);

CKINVDCx14_ASAP7_75t_R g1431 ( 
.A(n_1225),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1353),
.A2(n_657),
.B(n_179),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1378),
.A2(n_657),
.B(n_188),
.Y(n_1433)
);

AO31x2_ASAP7_75t_L g1434 ( 
.A1(n_1362),
.A2(n_657),
.A3(n_38),
.B(n_40),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1329),
.A2(n_686),
.B(n_646),
.C(n_40),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1354),
.A2(n_646),
.B(n_38),
.C(n_43),
.Y(n_1436)
);

AOI221xp5_ASAP7_75t_SL g1437 ( 
.A1(n_1226),
.A2(n_37),
.B1(n_44),
.B2(n_49),
.C(n_50),
.Y(n_1437)
);

BUFx12f_ASAP7_75t_L g1438 ( 
.A(n_1265),
.Y(n_1438)
);

O2A1O1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1268),
.A2(n_37),
.B(n_44),
.C(n_52),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1378),
.A2(n_161),
.B(n_230),
.Y(n_1440)
);

AO32x2_ASAP7_75t_L g1441 ( 
.A1(n_1252),
.A2(n_53),
.A3(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1286),
.A2(n_646),
.B(n_228),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1265),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1335),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1278),
.B(n_53),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1250),
.B(n_54),
.Y(n_1446)
);

AOI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1237),
.A2(n_646),
.B(n_226),
.Y(n_1447)
);

OAI22x1_ASAP7_75t_L g1448 ( 
.A1(n_1272),
.A2(n_57),
.B1(n_63),
.B2(n_64),
.Y(n_1448)
);

AO31x2_ASAP7_75t_L g1449 ( 
.A1(n_1299),
.A2(n_57),
.A3(n_64),
.B(n_68),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1286),
.A2(n_646),
.B1(n_69),
.B2(n_70),
.Y(n_1450)
);

A2O1A1Ixp33_ASAP7_75t_L g1451 ( 
.A1(n_1312),
.A2(n_1368),
.B(n_1319),
.C(n_1334),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1237),
.A2(n_128),
.B(n_224),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1298),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1274),
.A2(n_68),
.B(n_71),
.C(n_72),
.Y(n_1454)
);

A2O1A1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1297),
.A2(n_646),
.B(n_73),
.C(n_74),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1359),
.A2(n_135),
.B(n_214),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1276),
.Y(n_1457)
);

AO31x2_ASAP7_75t_L g1458 ( 
.A1(n_1299),
.A2(n_71),
.A3(n_77),
.B(n_79),
.Y(n_1458)
);

AO31x2_ASAP7_75t_L g1459 ( 
.A1(n_1348),
.A2(n_77),
.A3(n_82),
.B(n_83),
.Y(n_1459)
);

AO32x2_ASAP7_75t_L g1460 ( 
.A1(n_1252),
.A2(n_83),
.A3(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_1460)
);

O2A1O1Ixp5_ASAP7_75t_L g1461 ( 
.A1(n_1363),
.A2(n_1232),
.B(n_1359),
.C(n_1328),
.Y(n_1461)
);

A2O1A1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1339),
.A2(n_88),
.B(n_89),
.C(n_90),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_SL g1463 ( 
.A1(n_1370),
.A2(n_151),
.B(n_206),
.C(n_196),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1286),
.A2(n_142),
.B(n_193),
.Y(n_1464)
);

AO21x2_ASAP7_75t_L g1465 ( 
.A1(n_1327),
.A2(n_140),
.B(n_165),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1302),
.A2(n_137),
.B(n_160),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1302),
.A2(n_134),
.B(n_145),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1302),
.A2(n_88),
.B1(n_92),
.B2(n_95),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1314),
.A2(n_215),
.B(n_158),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1325),
.Y(n_1470)
);

INVx6_ASAP7_75t_L g1471 ( 
.A(n_1254),
.Y(n_1471)
);

BUFx8_ASAP7_75t_L g1472 ( 
.A(n_1244),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1302),
.A2(n_1243),
.B(n_1269),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1279),
.A2(n_1273),
.B(n_1366),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1256),
.A2(n_1331),
.B(n_1345),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1338),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1260),
.Y(n_1477)
);

A2O1A1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1355),
.A2(n_1344),
.B(n_1349),
.C(n_1263),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1291),
.Y(n_1479)
);

NAND2x2_ASAP7_75t_L g1480 ( 
.A(n_1275),
.B(n_1352),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1301),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1288),
.Y(n_1482)
);

BUFx2_ASAP7_75t_R g1483 ( 
.A(n_1272),
.Y(n_1483)
);

BUFx4f_ASAP7_75t_SL g1484 ( 
.A(n_1318),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1262),
.B(n_1336),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1310),
.A2(n_1252),
.B(n_1284),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1256),
.A2(n_1331),
.B(n_1345),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1325),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1316),
.Y(n_1489)
);

BUFx8_ASAP7_75t_L g1490 ( 
.A(n_1316),
.Y(n_1490)
);

AO32x2_ASAP7_75t_L g1491 ( 
.A1(n_1313),
.A2(n_1306),
.A3(n_1304),
.B1(n_1367),
.B2(n_1308),
.Y(n_1491)
);

NAND3xp33_ASAP7_75t_SL g1492 ( 
.A(n_1231),
.B(n_1241),
.C(n_1337),
.Y(n_1492)
);

CKINVDCx16_ASAP7_75t_R g1493 ( 
.A(n_1236),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1361),
.B(n_1373),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1374),
.B(n_1320),
.Y(n_1495)
);

O2A1O1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1360),
.A2(n_1337),
.B(n_1241),
.C(n_1264),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1296),
.B(n_1333),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1282),
.A2(n_1327),
.B(n_1376),
.Y(n_1498)
);

NOR2xp67_ASAP7_75t_L g1499 ( 
.A(n_1303),
.B(n_1300),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1309),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1228),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1317),
.A2(n_1259),
.B(n_1280),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1255),
.B(n_1309),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1357),
.A2(n_1348),
.B(n_1259),
.Y(n_1504)
);

NAND2xp33_ASAP7_75t_L g1505 ( 
.A(n_1340),
.B(n_1287),
.Y(n_1505)
);

AO31x2_ASAP7_75t_L g1506 ( 
.A1(n_1357),
.A2(n_1317),
.A3(n_1326),
.B(n_1371),
.Y(n_1506)
);

INVx4_ASAP7_75t_L g1507 ( 
.A(n_1224),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1255),
.A2(n_1321),
.B1(n_1341),
.B2(n_1309),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1343),
.A2(n_1326),
.B(n_1246),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1343),
.A2(n_1381),
.B(n_1382),
.Y(n_1510)
);

NOR2x1_ASAP7_75t_SL g1511 ( 
.A(n_1300),
.B(n_1255),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1356),
.A2(n_1257),
.B(n_1347),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1322),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1322),
.Y(n_1514)
);

OAI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1360),
.A2(n_1369),
.B1(n_1305),
.B2(n_1332),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1332),
.B(n_1305),
.Y(n_1516)
);

NAND2xp33_ASAP7_75t_L g1517 ( 
.A(n_1321),
.B(n_1341),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1330),
.B(n_1350),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1246),
.A2(n_1283),
.B(n_1290),
.Y(n_1519)
);

OAI22x1_ASAP7_75t_L g1520 ( 
.A1(n_1350),
.A2(n_1295),
.B1(n_1229),
.B2(n_1227),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1229),
.Y(n_1521)
);

AOI211x1_ASAP7_75t_L g1522 ( 
.A1(n_1311),
.A2(n_1356),
.B(n_1364),
.C(n_1351),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1372),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1224),
.B(n_1227),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1230),
.A2(n_1351),
.B(n_1315),
.Y(n_1525)
);

O2A1O1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1230),
.A2(n_1315),
.B(n_1372),
.C(n_1307),
.Y(n_1526)
);

BUFx10_ASAP7_75t_L g1527 ( 
.A(n_1346),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1270),
.A2(n_1118),
.B(n_935),
.Y(n_1528)
);

AND2x6_ASAP7_75t_SL g1529 ( 
.A(n_1219),
.B(n_1181),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1221),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1267),
.B(n_1080),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1300),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1342),
.A2(n_1365),
.B(n_1353),
.Y(n_1533)
);

NOR2xp67_ASAP7_75t_L g1534 ( 
.A(n_1238),
.B(n_864),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1238),
.B(n_708),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1270),
.A2(n_1118),
.B(n_935),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1235),
.A2(n_1118),
.B(n_1267),
.Y(n_1537)
);

AO22x2_ASAP7_75t_L g1538 ( 
.A1(n_1226),
.A2(n_1071),
.B1(n_1360),
.B2(n_1039),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1270),
.A2(n_1118),
.B(n_935),
.Y(n_1539)
);

INVx2_ASAP7_75t_SL g1540 ( 
.A(n_1298),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1292),
.Y(n_1541)
);

INVxp67_ASAP7_75t_SL g1542 ( 
.A(n_1372),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1270),
.A2(n_1118),
.B(n_935),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_SL g1544 ( 
.A1(n_1267),
.A2(n_805),
.B(n_1181),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1221),
.Y(n_1545)
);

AO31x2_ASAP7_75t_L g1546 ( 
.A1(n_1270),
.A2(n_1052),
.A3(n_1187),
.B(n_1247),
.Y(n_1546)
);

A2O1A1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_1267),
.A2(n_1118),
.B(n_1235),
.C(n_1092),
.Y(n_1547)
);

AO31x2_ASAP7_75t_L g1548 ( 
.A1(n_1270),
.A2(n_1052),
.A3(n_1187),
.B(n_1247),
.Y(n_1548)
);

O2A1O1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1235),
.A2(n_1118),
.B(n_1267),
.C(n_699),
.Y(n_1549)
);

AOI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1270),
.A2(n_1118),
.B(n_935),
.Y(n_1550)
);

AO32x2_ASAP7_75t_L g1551 ( 
.A1(n_1220),
.A2(n_1090),
.A3(n_1071),
.B1(n_1226),
.B2(n_989),
.Y(n_1551)
);

AOI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1270),
.A2(n_1118),
.B(n_935),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1270),
.A2(n_1118),
.B(n_935),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1270),
.A2(n_1118),
.B(n_935),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1267),
.B(n_1080),
.Y(n_1555)
);

CKINVDCx8_ASAP7_75t_R g1556 ( 
.A(n_1225),
.Y(n_1556)
);

CKINVDCx11_ASAP7_75t_R g1557 ( 
.A(n_1222),
.Y(n_1557)
);

AO31x2_ASAP7_75t_L g1558 ( 
.A1(n_1270),
.A2(n_1052),
.A3(n_1187),
.B(n_1247),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1270),
.A2(n_1118),
.B(n_935),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1267),
.B(n_1080),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1342),
.A2(n_1365),
.B(n_1353),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1324),
.Y(n_1562)
);

AOI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1342),
.A2(n_1353),
.B(n_1237),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1490),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1406),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1537),
.A2(n_1538),
.B1(n_1492),
.B2(n_1424),
.Y(n_1566)
);

OAI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1544),
.A2(n_1531),
.B1(n_1560),
.B2(n_1555),
.Y(n_1567)
);

OAI22x1_ASAP7_75t_L g1568 ( 
.A1(n_1503),
.A2(n_1422),
.B1(n_1500),
.B2(n_1429),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1547),
.A2(n_1387),
.B1(n_1549),
.B2(n_1535),
.Y(n_1569)
);

OAI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1445),
.A2(n_1448),
.B1(n_1494),
.B2(n_1493),
.Y(n_1570)
);

OAI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1468),
.A2(n_1450),
.B1(n_1394),
.B2(n_1457),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1538),
.A2(n_1446),
.B1(n_1515),
.B2(n_1457),
.Y(n_1572)
);

INVx6_ASAP7_75t_L g1573 ( 
.A(n_1490),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1516),
.A2(n_1412),
.B1(n_1383),
.B2(n_1385),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1392),
.A2(n_1523),
.B1(n_1386),
.B2(n_1456),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_1557),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1383),
.A2(n_1385),
.B1(n_1562),
.B2(n_1444),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1408),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1562),
.A2(n_1530),
.B1(n_1545),
.B2(n_1510),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1451),
.A2(n_1534),
.B1(n_1518),
.B2(n_1481),
.Y(n_1580)
);

CKINVDCx6p67_ASAP7_75t_R g1581 ( 
.A(n_1438),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1478),
.A2(n_1388),
.B1(n_1503),
.B2(n_1482),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1397),
.Y(n_1583)
);

OAI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1485),
.A2(n_1495),
.B1(n_1401),
.B2(n_1405),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1410),
.B(n_1399),
.Y(n_1585)
);

INVx11_ASAP7_75t_L g1586 ( 
.A(n_1472),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1556),
.A2(n_1499),
.B1(n_1480),
.B2(n_1501),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1523),
.A2(n_1386),
.B1(n_1542),
.B2(n_1511),
.Y(n_1588)
);

INVx4_ASAP7_75t_L g1589 ( 
.A(n_1418),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1470),
.A2(n_1488),
.B1(n_1476),
.B2(n_1512),
.Y(n_1590)
);

OAI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1414),
.A2(n_1484),
.B1(n_1513),
.B2(n_1514),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1497),
.Y(n_1592)
);

BUFx12f_ASAP7_75t_L g1593 ( 
.A(n_1472),
.Y(n_1593)
);

BUFx8_ASAP7_75t_L g1594 ( 
.A(n_1541),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1483),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1470),
.A2(n_1488),
.B1(n_1396),
.B2(n_1527),
.Y(n_1596)
);

BUFx6f_ASAP7_75t_SL g1597 ( 
.A(n_1541),
.Y(n_1597)
);

INVx6_ASAP7_75t_L g1598 ( 
.A(n_1421),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1449),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1527),
.A2(n_1469),
.B1(n_1403),
.B2(n_1474),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1453),
.B(n_1540),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1477),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1477),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1529),
.B(n_1479),
.Y(n_1604)
);

BUFx8_ASAP7_75t_L g1605 ( 
.A(n_1477),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1462),
.B(n_1435),
.Y(n_1606)
);

BUFx10_ASAP7_75t_L g1607 ( 
.A(n_1420),
.Y(n_1607)
);

BUFx6f_ASAP7_75t_SL g1608 ( 
.A(n_1443),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1521),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1532),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1421),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1471),
.Y(n_1612)
);

INVx11_ASAP7_75t_L g1613 ( 
.A(n_1471),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1469),
.A2(n_1465),
.B1(n_1525),
.B2(n_1536),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1431),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1449),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1465),
.A2(n_1543),
.B1(n_1539),
.B2(n_1552),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1496),
.B(n_1425),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1449),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1524),
.B(n_1443),
.Y(n_1620)
);

INVx6_ASAP7_75t_L g1621 ( 
.A(n_1421),
.Y(n_1621)
);

OAI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1508),
.A2(n_1441),
.B1(n_1460),
.B2(n_1437),
.Y(n_1622)
);

CKINVDCx20_ASAP7_75t_R g1623 ( 
.A(n_1411),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1443),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1528),
.A2(n_1550),
.B1(n_1559),
.B2(n_1554),
.Y(n_1625)
);

CKINVDCx16_ASAP7_75t_R g1626 ( 
.A(n_1489),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1404),
.A2(n_1391),
.B1(n_1522),
.B2(n_1526),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1458),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_SL g1629 ( 
.A1(n_1517),
.A2(n_1452),
.B1(n_1440),
.B2(n_1505),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1553),
.A2(n_1415),
.B1(n_1423),
.B2(n_1520),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1458),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1489),
.Y(n_1632)
);

INVx6_ASAP7_75t_L g1633 ( 
.A(n_1507),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1532),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_SL g1635 ( 
.A1(n_1551),
.A2(n_1439),
.B1(n_1454),
.B2(n_1467),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1507),
.Y(n_1636)
);

CKINVDCx11_ASAP7_75t_R g1637 ( 
.A(n_1459),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1389),
.A2(n_1400),
.B(n_1402),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1459),
.Y(n_1639)
);

NAND2x1p5_ASAP7_75t_L g1640 ( 
.A(n_1519),
.B(n_1509),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1464),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1498),
.A2(n_1551),
.B1(n_1502),
.B2(n_1466),
.Y(n_1642)
);

AOI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1436),
.A2(n_1455),
.B1(n_1463),
.B2(n_1473),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1434),
.Y(n_1644)
);

BUFx2_ASAP7_75t_SL g1645 ( 
.A(n_1442),
.Y(n_1645)
);

INVx6_ASAP7_75t_L g1646 ( 
.A(n_1395),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1407),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1407),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1486),
.A2(n_1441),
.B1(n_1460),
.B2(n_1413),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1441),
.A2(n_1460),
.B1(n_1487),
.B2(n_1475),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1426),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1447),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1504),
.A2(n_1416),
.B1(n_1430),
.B2(n_1409),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1426),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1416),
.A2(n_1433),
.B1(n_1384),
.B2(n_1533),
.Y(n_1655)
);

INVx6_ASAP7_75t_L g1656 ( 
.A(n_1461),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1419),
.B(n_1558),
.Y(n_1657)
);

BUFx12f_ASAP7_75t_L g1658 ( 
.A(n_1428),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1432),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1427),
.Y(n_1660)
);

INVx4_ASAP7_75t_L g1661 ( 
.A(n_1506),
.Y(n_1661)
);

CKINVDCx20_ASAP7_75t_R g1662 ( 
.A(n_1546),
.Y(n_1662)
);

INVx6_ASAP7_75t_L g1663 ( 
.A(n_1546),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1546),
.Y(n_1664)
);

BUFx8_ASAP7_75t_SL g1665 ( 
.A(n_1563),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1417),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1561),
.A2(n_1491),
.B1(n_1390),
.B2(n_1548),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1491),
.A2(n_1390),
.B1(n_1548),
.B2(n_1558),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1548),
.B(n_1558),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1417),
.Y(n_1670)
);

CKINVDCx11_ASAP7_75t_R g1671 ( 
.A(n_1390),
.Y(n_1671)
);

BUFx12f_ASAP7_75t_L g1672 ( 
.A(n_1506),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1506),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1398),
.Y(n_1674)
);

CKINVDCx11_ASAP7_75t_R g1675 ( 
.A(n_1491),
.Y(n_1675)
);

BUFx10_ASAP7_75t_L g1676 ( 
.A(n_1398),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1398),
.B(n_1234),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1393),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1557),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_SL g1680 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1547),
.A2(n_1118),
.B1(n_1387),
.B2(n_1537),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1393),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_SL g1684 ( 
.A1(n_1493),
.A2(n_805),
.B1(n_1267),
.B2(n_965),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1393),
.Y(n_1685)
);

BUFx4f_ASAP7_75t_L g1686 ( 
.A(n_1418),
.Y(n_1686)
);

OAI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1537),
.A2(n_698),
.B1(n_1544),
.B2(n_781),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1393),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1547),
.A2(n_1118),
.B1(n_1387),
.B2(n_1537),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1393),
.Y(n_1690)
);

BUFx12f_ASAP7_75t_L g1691 ( 
.A(n_1557),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1393),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_SL g1694 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1531),
.B(n_1267),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1696)
);

BUFx10_ASAP7_75t_L g1697 ( 
.A(n_1420),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_SL g1698 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1393),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1393),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1484),
.Y(n_1702)
);

CKINVDCx20_ASAP7_75t_R g1703 ( 
.A(n_1557),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1535),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1706)
);

INVx6_ASAP7_75t_L g1707 ( 
.A(n_1490),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1490),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1393),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1547),
.A2(n_1118),
.B1(n_1387),
.B2(n_1537),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1393),
.Y(n_1711)
);

OAI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1547),
.A2(n_1118),
.B(n_1387),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1484),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1513),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1484),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_SL g1717 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1717)
);

BUFx2_ASAP7_75t_SL g1718 ( 
.A(n_1418),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_SL g1719 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1535),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1393),
.Y(n_1721)
);

OAI22xp5_ASAP7_75t_SL g1722 ( 
.A1(n_1493),
.A2(n_805),
.B1(n_1267),
.B2(n_965),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1393),
.Y(n_1723)
);

INVx8_ASAP7_75t_L g1724 ( 
.A(n_1421),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1547),
.A2(n_1118),
.B1(n_1387),
.B2(n_1537),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_L g1727 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1484),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1393),
.Y(n_1729)
);

BUFx3_ASAP7_75t_L g1730 ( 
.A(n_1490),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1531),
.B(n_1267),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1531),
.B(n_1234),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1484),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1393),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1393),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1393),
.Y(n_1737)
);

INVx4_ASAP7_75t_L g1738 ( 
.A(n_1418),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1393),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1393),
.Y(n_1740)
);

CKINVDCx16_ASAP7_75t_R g1741 ( 
.A(n_1493),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1537),
.A2(n_1267),
.B1(n_865),
.B2(n_698),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1547),
.A2(n_1118),
.B1(n_1387),
.B2(n_1537),
.Y(n_1744)
);

BUFx12f_ASAP7_75t_L g1745 ( 
.A(n_1557),
.Y(n_1745)
);

OR2x6_ASAP7_75t_L g1746 ( 
.A(n_1712),
.B(n_1672),
.Y(n_1746)
);

OAI21x1_ASAP7_75t_L g1747 ( 
.A1(n_1638),
.A2(n_1640),
.B(n_1653),
.Y(n_1747)
);

INVx11_ASAP7_75t_L g1748 ( 
.A(n_1594),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1599),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1616),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1677),
.B(n_1675),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1619),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1657),
.B(n_1669),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1628),
.Y(n_1754)
);

AOI222xp33_ASAP7_75t_L g1755 ( 
.A1(n_1687),
.A2(n_1684),
.B1(n_1722),
.B2(n_1726),
.C1(n_1681),
.C2(n_1744),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1576),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1670),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1631),
.Y(n_1758)
);

AOI21x1_ASAP7_75t_L g1759 ( 
.A1(n_1689),
.A2(n_1710),
.B(n_1644),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1639),
.Y(n_1760)
);

BUFx3_ASAP7_75t_L g1761 ( 
.A(n_1605),
.Y(n_1761)
);

INVx3_ASAP7_75t_L g1762 ( 
.A(n_1646),
.Y(n_1762)
);

OAI21x1_ASAP7_75t_L g1763 ( 
.A1(n_1640),
.A2(n_1653),
.B(n_1625),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1647),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1648),
.Y(n_1765)
);

INVxp33_ASAP7_75t_L g1766 ( 
.A(n_1585),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1674),
.Y(n_1767)
);

OAI21x1_ASAP7_75t_L g1768 ( 
.A1(n_1625),
.A2(n_1655),
.B(n_1617),
.Y(n_1768)
);

OAI21x1_ASAP7_75t_L g1769 ( 
.A1(n_1655),
.A2(n_1617),
.B(n_1614),
.Y(n_1769)
);

BUFx6f_ASAP7_75t_L g1770 ( 
.A(n_1611),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1567),
.B(n_1680),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1664),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1664),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1651),
.B(n_1654),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1675),
.B(n_1671),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1666),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1685),
.B(n_1583),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1646),
.Y(n_1778)
);

INVx2_ASAP7_75t_SL g1779 ( 
.A(n_1715),
.Y(n_1779)
);

NAND2x1_ASAP7_75t_L g1780 ( 
.A(n_1656),
.B(n_1646),
.Y(n_1780)
);

OR2x6_ASAP7_75t_L g1781 ( 
.A(n_1656),
.B(n_1568),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1663),
.Y(n_1782)
);

INVx3_ASAP7_75t_L g1783 ( 
.A(n_1663),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1663),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1671),
.B(n_1596),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1618),
.B(n_1596),
.Y(n_1786)
);

INVxp67_ASAP7_75t_L g1787 ( 
.A(n_1705),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1582),
.Y(n_1788)
);

INVx4_ASAP7_75t_L g1789 ( 
.A(n_1724),
.Y(n_1789)
);

AOI221xp5_ASAP7_75t_L g1790 ( 
.A1(n_1687),
.A2(n_1733),
.B1(n_1727),
.B2(n_1706),
.C(n_1700),
.Y(n_1790)
);

OAI21x1_ASAP7_75t_L g1791 ( 
.A1(n_1614),
.A2(n_1673),
.B(n_1630),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1662),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1676),
.Y(n_1793)
);

INVxp67_ASAP7_75t_SL g1794 ( 
.A(n_1584),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1673),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1650),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1565),
.Y(n_1797)
);

OA21x2_ASAP7_75t_L g1798 ( 
.A1(n_1650),
.A2(n_1649),
.B(n_1667),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1661),
.Y(n_1799)
);

INVx2_ASAP7_75t_SL g1800 ( 
.A(n_1598),
.Y(n_1800)
);

INVx2_ASAP7_75t_SL g1801 ( 
.A(n_1598),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1649),
.B(n_1566),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1661),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1637),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1656),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1578),
.Y(n_1806)
);

BUFx3_ASAP7_75t_L g1807 ( 
.A(n_1605),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1637),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1667),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1566),
.B(n_1572),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1567),
.A2(n_1569),
.B1(n_1717),
.B2(n_1698),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1682),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1668),
.B(n_1572),
.Y(n_1813)
);

OAI21x1_ASAP7_75t_L g1814 ( 
.A1(n_1630),
.A2(n_1642),
.B(n_1600),
.Y(n_1814)
);

AOI21x1_ASAP7_75t_L g1815 ( 
.A1(n_1627),
.A2(n_1606),
.B(n_1580),
.Y(n_1815)
);

BUFx2_ASAP7_75t_L g1816 ( 
.A(n_1665),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1688),
.Y(n_1817)
);

BUFx2_ASAP7_75t_L g1818 ( 
.A(n_1591),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1668),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1577),
.B(n_1574),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1720),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1577),
.Y(n_1822)
);

INVx4_ASAP7_75t_L g1823 ( 
.A(n_1724),
.Y(n_1823)
);

INVx3_ASAP7_75t_L g1824 ( 
.A(n_1659),
.Y(n_1824)
);

AO21x1_ASAP7_75t_L g1825 ( 
.A1(n_1622),
.A2(n_1571),
.B(n_1584),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1690),
.Y(n_1826)
);

OA21x2_ASAP7_75t_L g1827 ( 
.A1(n_1642),
.A2(n_1600),
.B(n_1574),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1692),
.Y(n_1828)
);

BUFx3_ASAP7_75t_L g1829 ( 
.A(n_1686),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1694),
.A2(n_1719),
.B(n_1727),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1699),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1701),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1709),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1721),
.Y(n_1834)
);

OAI21x1_ASAP7_75t_L g1835 ( 
.A1(n_1643),
.A2(n_1590),
.B(n_1579),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1729),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_SL g1837 ( 
.A1(n_1641),
.A2(n_1658),
.B1(n_1741),
.B2(n_1732),
.Y(n_1837)
);

OAI21x1_ASAP7_75t_L g1838 ( 
.A1(n_1590),
.A2(n_1579),
.B(n_1740),
.Y(n_1838)
);

INVx4_ASAP7_75t_L g1839 ( 
.A(n_1724),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1735),
.Y(n_1840)
);

OR2x6_ASAP7_75t_L g1841 ( 
.A(n_1645),
.B(n_1652),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1736),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1739),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1622),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1678),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1683),
.B(n_1693),
.Y(n_1846)
);

BUFx6f_ASAP7_75t_L g1847 ( 
.A(n_1611),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1711),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1723),
.B(n_1737),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1695),
.B(n_1731),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1592),
.Y(n_1851)
);

BUFx2_ASAP7_75t_L g1852 ( 
.A(n_1591),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1652),
.Y(n_1853)
);

INVx1_ASAP7_75t_SL g1854 ( 
.A(n_1609),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1660),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1620),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1683),
.B(n_1693),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1659),
.Y(n_1858)
);

AOI21x1_ASAP7_75t_L g1859 ( 
.A1(n_1610),
.A2(n_1632),
.B(n_1624),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1634),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1696),
.B(n_1700),
.Y(n_1861)
);

INVx2_ASAP7_75t_SL g1862 ( 
.A(n_1598),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1714),
.B(n_1728),
.Y(n_1863)
);

AO21x1_ASAP7_75t_L g1864 ( 
.A1(n_1571),
.A2(n_1570),
.B(n_1733),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1629),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1696),
.B(n_1713),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1635),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1575),
.Y(n_1868)
);

BUFx6f_ASAP7_75t_L g1869 ( 
.A(n_1611),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1703),
.Y(n_1870)
);

A2O1A1Ixp33_ASAP7_75t_L g1871 ( 
.A1(n_1704),
.A2(n_1743),
.B(n_1742),
.C(n_1725),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1570),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1704),
.A2(n_1713),
.B1(n_1706),
.B2(n_1743),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1725),
.B(n_1742),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1621),
.Y(n_1875)
);

AO21x2_ASAP7_75t_L g1876 ( 
.A1(n_1587),
.A2(n_1604),
.B(n_1601),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1621),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1626),
.B(n_1602),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1621),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1588),
.B(n_1603),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1608),
.Y(n_1881)
);

OAI21x1_ASAP7_75t_L g1882 ( 
.A1(n_1608),
.A2(n_1633),
.B(n_1597),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1636),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1636),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1633),
.Y(n_1885)
);

NAND2x1p5_ASAP7_75t_L g1886 ( 
.A(n_1589),
.B(n_1738),
.Y(n_1886)
);

OAI21x1_ASAP7_75t_L g1887 ( 
.A1(n_1633),
.A2(n_1597),
.B(n_1573),
.Y(n_1887)
);

INVx1_ASAP7_75t_SL g1888 ( 
.A(n_1716),
.Y(n_1888)
);

BUFx3_ASAP7_75t_L g1889 ( 
.A(n_1686),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1718),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1612),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_1679),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1594),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1573),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_1564),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1871),
.A2(n_1623),
.B(n_1595),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1792),
.B(n_1856),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_L g1898 ( 
.A(n_1850),
.B(n_1702),
.Y(n_1898)
);

INVxp67_ASAP7_75t_SL g1899 ( 
.A(n_1855),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1794),
.B(n_1707),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1822),
.B(n_1707),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1782),
.B(n_1564),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1888),
.B(n_1766),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1820),
.B(n_1573),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1751),
.B(n_1730),
.Y(n_1905)
);

A2O1A1Ixp33_ASAP7_75t_L g1906 ( 
.A1(n_1811),
.A2(n_1708),
.B(n_1730),
.C(n_1734),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1751),
.B(n_1708),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1753),
.B(n_1707),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1804),
.B(n_1697),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1782),
.B(n_1615),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1753),
.B(n_1581),
.Y(n_1911)
);

HB1xp67_ASAP7_75t_L g1912 ( 
.A(n_1779),
.Y(n_1912)
);

BUFx2_ASAP7_75t_SL g1913 ( 
.A(n_1761),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1804),
.B(n_1607),
.Y(n_1914)
);

BUFx4f_ASAP7_75t_SL g1915 ( 
.A(n_1761),
.Y(n_1915)
);

O2A1O1Ixp33_ASAP7_75t_SL g1916 ( 
.A1(n_1771),
.A2(n_1586),
.B(n_1593),
.C(n_1691),
.Y(n_1916)
);

BUFx2_ASAP7_75t_L g1917 ( 
.A(n_1821),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1808),
.B(n_1607),
.Y(n_1918)
);

AOI221xp5_ASAP7_75t_SL g1919 ( 
.A1(n_1830),
.A2(n_1613),
.B1(n_1697),
.B2(n_1745),
.C(n_1790),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1878),
.B(n_1775),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1846),
.A2(n_1768),
.B(n_1873),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1844),
.B(n_1855),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1756),
.Y(n_1923)
);

BUFx3_ASAP7_75t_L g1924 ( 
.A(n_1807),
.Y(n_1924)
);

A2O1A1Ixp33_ASAP7_75t_L g1925 ( 
.A1(n_1835),
.A2(n_1866),
.B(n_1857),
.C(n_1874),
.Y(n_1925)
);

A2O1A1Ixp33_ASAP7_75t_L g1926 ( 
.A1(n_1835),
.A2(n_1866),
.B(n_1857),
.C(n_1874),
.Y(n_1926)
);

OAI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1755),
.A2(n_1815),
.B(n_1861),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1777),
.Y(n_1928)
);

AOI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1864),
.A2(n_1810),
.B1(n_1876),
.B2(n_1837),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1863),
.B(n_1787),
.Y(n_1930)
);

A2O1A1Ixp33_ASAP7_75t_L g1931 ( 
.A1(n_1818),
.A2(n_1852),
.B(n_1814),
.C(n_1810),
.Y(n_1931)
);

AO21x2_ASAP7_75t_L g1932 ( 
.A1(n_1825),
.A2(n_1747),
.B(n_1769),
.Y(n_1932)
);

A2O1A1Ixp33_ASAP7_75t_L g1933 ( 
.A1(n_1818),
.A2(n_1852),
.B(n_1814),
.C(n_1867),
.Y(n_1933)
);

NAND4xp25_ASAP7_75t_L g1934 ( 
.A(n_1872),
.B(n_1867),
.C(n_1786),
.D(n_1844),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1783),
.B(n_1887),
.Y(n_1935)
);

O2A1O1Ixp33_ASAP7_75t_SL g1936 ( 
.A1(n_1780),
.A2(n_1881),
.B(n_1872),
.C(n_1786),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1854),
.B(n_1756),
.Y(n_1937)
);

OAI21x1_ASAP7_75t_L g1938 ( 
.A1(n_1747),
.A2(n_1763),
.B(n_1768),
.Y(n_1938)
);

OAI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1759),
.A2(n_1788),
.B(n_1838),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1785),
.B(n_1868),
.Y(n_1940)
);

A2O1A1Ixp33_ASAP7_75t_L g1941 ( 
.A1(n_1868),
.A2(n_1865),
.B(n_1802),
.C(n_1769),
.Y(n_1941)
);

OAI21xp33_ASAP7_75t_L g1942 ( 
.A1(n_1802),
.A2(n_1865),
.B(n_1746),
.Y(n_1942)
);

A2O1A1Ixp33_ASAP7_75t_L g1943 ( 
.A1(n_1791),
.A2(n_1864),
.B(n_1816),
.C(n_1838),
.Y(n_1943)
);

OA21x2_ASAP7_75t_L g1944 ( 
.A1(n_1791),
.A2(n_1763),
.B(n_1825),
.Y(n_1944)
);

AO32x2_ASAP7_75t_L g1945 ( 
.A1(n_1800),
.A2(n_1862),
.A3(n_1801),
.B1(n_1798),
.B2(n_1796),
.Y(n_1945)
);

OAI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1813),
.A2(n_1816),
.B1(n_1746),
.B2(n_1851),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1851),
.B(n_1819),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1876),
.A2(n_1746),
.B1(n_1781),
.B2(n_1894),
.Y(n_1948)
);

A2O1A1Ixp33_ASAP7_75t_L g1949 ( 
.A1(n_1813),
.A2(n_1805),
.B(n_1829),
.C(n_1889),
.Y(n_1949)
);

AO32x1_ASAP7_75t_L g1950 ( 
.A1(n_1795),
.A2(n_1773),
.A3(n_1772),
.B1(n_1749),
.B2(n_1750),
.Y(n_1950)
);

A2O1A1Ixp33_ASAP7_75t_L g1951 ( 
.A1(n_1805),
.A2(n_1889),
.B(n_1829),
.C(n_1762),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1870),
.B(n_1892),
.Y(n_1952)
);

OAI21x1_ASAP7_75t_L g1953 ( 
.A1(n_1759),
.A2(n_1887),
.B(n_1824),
.Y(n_1953)
);

OAI211xp5_ASAP7_75t_L g1954 ( 
.A1(n_1827),
.A2(n_1796),
.B(n_1891),
.C(n_1798),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_1870),
.Y(n_1955)
);

NAND2x1_ASAP7_75t_L g1956 ( 
.A(n_1805),
.B(n_1841),
.Y(n_1956)
);

NAND3xp33_ASAP7_75t_L g1957 ( 
.A(n_1827),
.B(n_1891),
.C(n_1817),
.Y(n_1957)
);

AOI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1876),
.A2(n_1781),
.B1(n_1894),
.B2(n_1762),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1783),
.B(n_1882),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1781),
.B(n_1797),
.Y(n_1960)
);

A2O1A1Ixp33_ASAP7_75t_L g1961 ( 
.A1(n_1762),
.A2(n_1778),
.B(n_1882),
.C(n_1881),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1809),
.B(n_1826),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1806),
.B(n_1812),
.Y(n_1963)
);

AOI22xp33_ASAP7_75t_L g1964 ( 
.A1(n_1880),
.A2(n_1827),
.B1(n_1778),
.B2(n_1895),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1826),
.B(n_1828),
.Y(n_1965)
);

AO21x1_ASAP7_75t_L g1966 ( 
.A1(n_1880),
.A2(n_1884),
.B(n_1883),
.Y(n_1966)
);

AND2x6_ASAP7_75t_L g1967 ( 
.A(n_1778),
.B(n_1784),
.Y(n_1967)
);

AOI22xp33_ASAP7_75t_SL g1968 ( 
.A1(n_1827),
.A2(n_1798),
.B1(n_1895),
.B2(n_1807),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1892),
.B(n_1893),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1749),
.Y(n_1970)
);

INVx1_ASAP7_75t_SL g1971 ( 
.A(n_1860),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_1748),
.Y(n_1972)
);

OAI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1853),
.A2(n_1859),
.B(n_1841),
.Y(n_1973)
);

AND2x4_ASAP7_75t_L g1974 ( 
.A(n_1828),
.B(n_1831),
.Y(n_1974)
);

A2O1A1Ixp33_ASAP7_75t_L g1975 ( 
.A1(n_1890),
.A2(n_1879),
.B(n_1893),
.C(n_1801),
.Y(n_1975)
);

AND2x2_ASAP7_75t_SL g1976 ( 
.A(n_1789),
.B(n_1823),
.Y(n_1976)
);

AO32x2_ASAP7_75t_L g1977 ( 
.A1(n_1800),
.A2(n_1862),
.A3(n_1798),
.B1(n_1839),
.B2(n_1823),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1833),
.B(n_1834),
.Y(n_1978)
);

OA21x2_ASAP7_75t_L g1979 ( 
.A1(n_1750),
.A2(n_1758),
.B(n_1752),
.Y(n_1979)
);

AO32x2_ASAP7_75t_L g1980 ( 
.A1(n_1789),
.A2(n_1823),
.A3(n_1839),
.B1(n_1754),
.B2(n_1758),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1754),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1831),
.B(n_1832),
.Y(n_1982)
);

HB1xp67_ASAP7_75t_L g1983 ( 
.A(n_1836),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_L g1984 ( 
.A(n_1877),
.B(n_1748),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1832),
.B(n_1843),
.Y(n_1985)
);

INVxp67_ASAP7_75t_SL g1986 ( 
.A(n_1776),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1979),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1979),
.Y(n_1988)
);

BUFx2_ASAP7_75t_L g1989 ( 
.A(n_1980),
.Y(n_1989)
);

HB1xp67_ASAP7_75t_L g1990 ( 
.A(n_1912),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1970),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1971),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1981),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1965),
.Y(n_1994)
);

NAND3xp33_ASAP7_75t_L g1995 ( 
.A(n_1919),
.B(n_1842),
.C(n_1840),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1965),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1982),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1899),
.B(n_1760),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1960),
.B(n_1928),
.Y(n_1999)
);

AND2x4_ASAP7_75t_L g2000 ( 
.A(n_1935),
.B(n_1858),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1935),
.B(n_1959),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1922),
.B(n_1767),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1983),
.Y(n_2003)
);

INVx3_ASAP7_75t_L g2004 ( 
.A(n_1959),
.Y(n_2004)
);

AOI22xp33_ASAP7_75t_L g2005 ( 
.A1(n_1927),
.A2(n_1877),
.B1(n_1841),
.B2(n_1793),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1977),
.B(n_1803),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1977),
.B(n_1799),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1977),
.B(n_1793),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1974),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1985),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1985),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1950),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1963),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1971),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1957),
.B(n_1757),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1978),
.Y(n_2016)
);

BUFx3_ASAP7_75t_L g2017 ( 
.A(n_1956),
.Y(n_2017)
);

BUFx6f_ASAP7_75t_L g2018 ( 
.A(n_1976),
.Y(n_2018)
);

AOI22xp5_ASAP7_75t_L g2019 ( 
.A1(n_1919),
.A2(n_1849),
.B1(n_1879),
.B2(n_1885),
.Y(n_2019)
);

AOI22xp33_ASAP7_75t_L g2020 ( 
.A1(n_1927),
.A2(n_1896),
.B1(n_1942),
.B2(n_1921),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1945),
.B(n_1764),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1898),
.B(n_1885),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1945),
.B(n_1764),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_1917),
.Y(n_2024)
);

OAI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1929),
.A2(n_1845),
.B1(n_1848),
.B2(n_1879),
.Y(n_2025)
);

AOI22xp33_ASAP7_75t_SL g2026 ( 
.A1(n_1896),
.A2(n_1875),
.B1(n_1770),
.B2(n_1847),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1957),
.B(n_1774),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1897),
.B(n_1774),
.Y(n_2028)
);

INVx4_ASAP7_75t_L g2029 ( 
.A(n_1967),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1962),
.Y(n_2030)
);

INVxp33_ASAP7_75t_L g2031 ( 
.A(n_1952),
.Y(n_2031)
);

BUFx2_ASAP7_75t_L g2032 ( 
.A(n_1980),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1945),
.B(n_1765),
.Y(n_2033)
);

INVxp67_ASAP7_75t_SL g2034 ( 
.A(n_1986),
.Y(n_2034)
);

INVxp67_ASAP7_75t_SL g2035 ( 
.A(n_1947),
.Y(n_2035)
);

OAI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_2020),
.A2(n_1906),
.B1(n_1931),
.B2(n_1933),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1987),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1993),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1992),
.B(n_1925),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2014),
.B(n_1926),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_2018),
.B(n_2019),
.Y(n_2041)
);

OR2x2_ASAP7_75t_L g2042 ( 
.A(n_2028),
.B(n_2027),
.Y(n_2042)
);

NOR2x1_ASAP7_75t_L g2043 ( 
.A(n_2017),
.B(n_1995),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_2018),
.B(n_1958),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_2018),
.B(n_1948),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_2024),
.B(n_1941),
.Y(n_2046)
);

NOR2xp33_ASAP7_75t_L g2047 ( 
.A(n_2031),
.B(n_1911),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_2035),
.B(n_1921),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_2028),
.B(n_1954),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1987),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1990),
.B(n_2013),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_2027),
.B(n_1954),
.Y(n_2052)
);

OR2x6_ASAP7_75t_SL g2053 ( 
.A(n_2025),
.B(n_1904),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1987),
.Y(n_2054)
);

OAI221xp5_ASAP7_75t_SL g2055 ( 
.A1(n_2019),
.A2(n_1943),
.B1(n_2005),
.B2(n_1964),
.C(n_1934),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_2001),
.B(n_1968),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2001),
.B(n_1980),
.Y(n_2057)
);

BUFx3_ASAP7_75t_L g2058 ( 
.A(n_2017),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_R g2059 ( 
.A(n_2018),
.B(n_1923),
.Y(n_2059)
);

OAI31xp33_ASAP7_75t_L g2060 ( 
.A1(n_2025),
.A2(n_1946),
.A3(n_1949),
.B(n_1961),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2009),
.B(n_1920),
.Y(n_2061)
);

AOI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_2022),
.A2(n_1946),
.B1(n_1934),
.B2(n_1900),
.Y(n_2062)
);

AOI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_2018),
.A2(n_1940),
.B1(n_1904),
.B2(n_1909),
.Y(n_2063)
);

INVx3_ASAP7_75t_L g2064 ( 
.A(n_2017),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_2009),
.B(n_1944),
.Y(n_2065)
);

AOI221xp5_ASAP7_75t_L g2066 ( 
.A1(n_1989),
.A2(n_1901),
.B1(n_1900),
.B2(n_1936),
.C(n_1939),
.Y(n_2066)
);

OR2x2_ASAP7_75t_SL g2067 ( 
.A(n_2018),
.B(n_1944),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_2003),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_2004),
.B(n_1953),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_1995),
.A2(n_1916),
.B(n_1951),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1988),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2015),
.B(n_1932),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2004),
.B(n_1999),
.Y(n_2073)
);

OR2x2_ASAP7_75t_L g2074 ( 
.A(n_2015),
.B(n_1932),
.Y(n_2074)
);

OR2x6_ASAP7_75t_L g2075 ( 
.A(n_2029),
.B(n_1938),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1999),
.B(n_1939),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1988),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1991),
.Y(n_2078)
);

OR2x6_ASAP7_75t_L g2079 ( 
.A(n_2029),
.B(n_1973),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1989),
.B(n_1914),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2032),
.B(n_1918),
.Y(n_2081)
);

NAND2x1_ASAP7_75t_L g2082 ( 
.A(n_2029),
.B(n_1967),
.Y(n_2082)
);

BUFx6f_ASAP7_75t_L g2083 ( 
.A(n_2000),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_2032),
.B(n_1962),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_SL g2085 ( 
.A(n_2034),
.B(n_1955),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_2010),
.B(n_1908),
.Y(n_2086)
);

AOI21xp5_ASAP7_75t_L g2087 ( 
.A1(n_1998),
.A2(n_1975),
.B(n_1973),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2016),
.B(n_1911),
.Y(n_2088)
);

INVxp67_ASAP7_75t_SL g2089 ( 
.A(n_2002),
.Y(n_2089)
);

INVx1_ASAP7_75t_SL g2090 ( 
.A(n_2049),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2057),
.B(n_2008),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2057),
.B(n_2008),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2037),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2071),
.Y(n_2094)
);

NAND4xp25_ASAP7_75t_L g2095 ( 
.A(n_2055),
.B(n_1930),
.C(n_1901),
.D(n_1903),
.Y(n_2095)
);

INVx1_ASAP7_75t_SL g2096 ( 
.A(n_2049),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2037),
.Y(n_2097)
);

OR2x2_ASAP7_75t_L g2098 ( 
.A(n_2072),
.B(n_2012),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2071),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2050),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2038),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2048),
.B(n_2030),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2089),
.B(n_2030),
.Y(n_2103)
);

NAND2xp33_ASAP7_75t_R g2104 ( 
.A(n_2059),
.B(n_1972),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2038),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2065),
.B(n_2006),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2076),
.B(n_2073),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2042),
.B(n_1994),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2076),
.B(n_2007),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2056),
.B(n_2021),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2056),
.B(n_2021),
.Y(n_2111)
);

AND2x4_ASAP7_75t_L g2112 ( 
.A(n_2075),
.B(n_2069),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_2072),
.B(n_2074),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2080),
.B(n_2023),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2080),
.B(n_2023),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2042),
.B(n_1994),
.Y(n_2116)
);

AND2x4_ASAP7_75t_L g2117 ( 
.A(n_2075),
.B(n_2033),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_2054),
.Y(n_2118)
);

INVx2_ASAP7_75t_SL g2119 ( 
.A(n_2083),
.Y(n_2119)
);

BUFx3_ASAP7_75t_L g2120 ( 
.A(n_2082),
.Y(n_2120)
);

INVx4_ASAP7_75t_L g2121 ( 
.A(n_2079),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2068),
.B(n_1996),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2081),
.B(n_2033),
.Y(n_2123)
);

INVx2_ASAP7_75t_SL g2124 ( 
.A(n_2083),
.Y(n_2124)
);

HB1xp67_ASAP7_75t_L g2125 ( 
.A(n_2077),
.Y(n_2125)
);

A2O1A1Ixp33_ASAP7_75t_SL g2126 ( 
.A1(n_2036),
.A2(n_1984),
.B(n_1937),
.C(n_1969),
.Y(n_2126)
);

AOI22xp33_ASAP7_75t_L g2127 ( 
.A1(n_2039),
.A2(n_2026),
.B1(n_1966),
.B2(n_1910),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2081),
.B(n_2010),
.Y(n_2128)
);

CKINVDCx5p33_ASAP7_75t_R g2129 ( 
.A(n_2058),
.Y(n_2129)
);

AND2x4_ASAP7_75t_L g2130 ( 
.A(n_2075),
.B(n_2012),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2053),
.B(n_2011),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2053),
.B(n_2011),
.Y(n_2132)
);

OR2x2_ASAP7_75t_L g2133 ( 
.A(n_2074),
.B(n_2052),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2077),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2087),
.B(n_1996),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2078),
.B(n_1997),
.Y(n_2136)
);

OR2x2_ASAP7_75t_L g2137 ( 
.A(n_2090),
.B(n_2052),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_2090),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2110),
.B(n_2064),
.Y(n_2139)
);

OR2x6_ASAP7_75t_L g2140 ( 
.A(n_2121),
.B(n_2043),
.Y(n_2140)
);

NOR2xp33_ASAP7_75t_L g2141 ( 
.A(n_2095),
.B(n_1915),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2094),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2094),
.Y(n_2143)
);

NAND2x1p5_ASAP7_75t_L g2144 ( 
.A(n_2120),
.B(n_2043),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2135),
.B(n_2040),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2094),
.Y(n_2146)
);

INVx3_ASAP7_75t_SL g2147 ( 
.A(n_2129),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_2096),
.B(n_2084),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2110),
.B(n_2064),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2135),
.B(n_2046),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_2096),
.B(n_2084),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2134),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2134),
.Y(n_2153)
);

BUFx3_ASAP7_75t_L g2154 ( 
.A(n_2129),
.Y(n_2154)
);

INVxp67_ASAP7_75t_L g2155 ( 
.A(n_2095),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2099),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2099),
.Y(n_2157)
);

OAI21xp33_ASAP7_75t_L g2158 ( 
.A1(n_2127),
.A2(n_2132),
.B(n_2131),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2110),
.B(n_2064),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2099),
.Y(n_2160)
);

AOI221xp5_ASAP7_75t_L g2161 ( 
.A1(n_2126),
.A2(n_2066),
.B1(n_2041),
.B2(n_2044),
.C(n_2045),
.Y(n_2161)
);

INVxp67_ASAP7_75t_L g2162 ( 
.A(n_2102),
.Y(n_2162)
);

OAI31xp33_ASAP7_75t_L g2163 ( 
.A1(n_2126),
.A2(n_2070),
.A3(n_2060),
.B(n_2085),
.Y(n_2163)
);

INVxp67_ASAP7_75t_SL g2164 ( 
.A(n_2102),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2131),
.B(n_2086),
.Y(n_2165)
);

INVx1_ASAP7_75t_SL g2166 ( 
.A(n_2120),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2131),
.B(n_2086),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2136),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2136),
.Y(n_2169)
);

INVx2_ASAP7_75t_SL g2170 ( 
.A(n_2120),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2125),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2125),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2111),
.B(n_2058),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2122),
.Y(n_2174)
);

OR2x2_ASAP7_75t_L g2175 ( 
.A(n_2133),
.B(n_2067),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2122),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2101),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2101),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2134),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2132),
.B(n_2088),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2101),
.Y(n_2181)
);

NOR2xp33_ASAP7_75t_L g2182 ( 
.A(n_2121),
.B(n_2047),
.Y(n_2182)
);

HB1xp67_ASAP7_75t_L g2183 ( 
.A(n_2132),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_SL g2184 ( 
.A(n_2127),
.B(n_2062),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2111),
.B(n_2061),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2111),
.B(n_2061),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2105),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2120),
.B(n_2079),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2150),
.B(n_2107),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2139),
.B(n_2149),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2143),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2143),
.Y(n_2192)
);

OR2x2_ASAP7_75t_L g2193 ( 
.A(n_2137),
.B(n_2133),
.Y(n_2193)
);

HB1xp67_ASAP7_75t_L g2194 ( 
.A(n_2183),
.Y(n_2194)
);

NOR2xp67_ASAP7_75t_L g2195 ( 
.A(n_2138),
.B(n_2121),
.Y(n_2195)
);

INVxp67_ASAP7_75t_SL g2196 ( 
.A(n_2144),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2139),
.B(n_2119),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2149),
.B(n_2119),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2145),
.B(n_2107),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2159),
.B(n_2119),
.Y(n_2200)
);

NOR2x1_ASAP7_75t_L g2201 ( 
.A(n_2154),
.B(n_2140),
.Y(n_2201)
);

OR2x6_ASAP7_75t_L g2202 ( 
.A(n_2140),
.B(n_1913),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2142),
.Y(n_2203)
);

NOR2x1_ASAP7_75t_L g2204 ( 
.A(n_2154),
.B(n_1924),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2159),
.Y(n_2205)
);

OAI22xp5_ASAP7_75t_L g2206 ( 
.A1(n_2184),
.A2(n_2062),
.B1(n_2067),
.B2(n_2079),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2173),
.B(n_2119),
.Y(n_2207)
);

NAND2x1_ASAP7_75t_L g2208 ( 
.A(n_2140),
.B(n_2117),
.Y(n_2208)
);

INVxp67_ASAP7_75t_SL g2209 ( 
.A(n_2144),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2146),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2173),
.B(n_2091),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2155),
.B(n_2107),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2188),
.B(n_2091),
.Y(n_2213)
);

OR2x2_ASAP7_75t_L g2214 ( 
.A(n_2137),
.B(n_2133),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2156),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2161),
.B(n_2103),
.Y(n_2216)
);

OR2x2_ASAP7_75t_L g2217 ( 
.A(n_2148),
.B(n_2098),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_SL g2218 ( 
.A(n_2163),
.B(n_2121),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2184),
.B(n_2103),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2157),
.Y(n_2220)
);

NAND2xp33_ASAP7_75t_R g2221 ( 
.A(n_2140),
.B(n_2141),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2158),
.B(n_2128),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2162),
.B(n_2128),
.Y(n_2223)
);

INVx2_ASAP7_75t_SL g2224 ( 
.A(n_2170),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_L g2225 ( 
.A(n_2147),
.B(n_1910),
.Y(n_2225)
);

INVx1_ASAP7_75t_SL g2226 ( 
.A(n_2147),
.Y(n_2226)
);

AND3x2_ASAP7_75t_L g2227 ( 
.A(n_2188),
.B(n_2104),
.C(n_1907),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2164),
.B(n_2128),
.Y(n_2228)
);

OAI221xp5_ASAP7_75t_L g2229 ( 
.A1(n_2182),
.A2(n_2121),
.B1(n_2063),
.B2(n_2104),
.C(n_2079),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_L g2230 ( 
.A(n_2180),
.B(n_2121),
.Y(n_2230)
);

NOR2xp33_ASAP7_75t_L g2231 ( 
.A(n_2226),
.B(n_2216),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2194),
.Y(n_2232)
);

XOR2x2_ASAP7_75t_L g2233 ( 
.A(n_2204),
.B(n_2144),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2219),
.B(n_2174),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_2218),
.B(n_2166),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2211),
.Y(n_2236)
);

NAND3xp33_ASAP7_75t_L g2237 ( 
.A(n_2201),
.B(n_2175),
.C(n_2170),
.Y(n_2237)
);

OAI221xp5_ASAP7_75t_L g2238 ( 
.A1(n_2206),
.A2(n_2175),
.B1(n_2176),
.B2(n_2151),
.C(n_2148),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2191),
.Y(n_2239)
);

AOI22xp5_ASAP7_75t_L g2240 ( 
.A1(n_2221),
.A2(n_2229),
.B1(n_2227),
.B2(n_2230),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2212),
.B(n_2165),
.Y(n_2241)
);

OAI22xp33_ASAP7_75t_L g2242 ( 
.A1(n_2222),
.A2(n_2195),
.B1(n_2214),
.B2(n_2193),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2213),
.B(n_2167),
.Y(n_2243)
);

BUFx3_ASAP7_75t_L g2244 ( 
.A(n_2225),
.Y(n_2244)
);

AOI221xp5_ASAP7_75t_L g2245 ( 
.A1(n_2213),
.A2(n_2168),
.B1(n_2169),
.B2(n_2171),
.C(n_2172),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2191),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_SL g2247 ( 
.A(n_2193),
.B(n_2214),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2192),
.Y(n_2248)
);

INVxp67_ASAP7_75t_L g2249 ( 
.A(n_2196),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2203),
.Y(n_2250)
);

AOI222xp33_ASAP7_75t_L g2251 ( 
.A1(n_2228),
.A2(n_2130),
.B1(n_2186),
.B2(n_2185),
.C1(n_2117),
.C2(n_2092),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2211),
.B(n_2151),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_2189),
.B(n_2108),
.Y(n_2253)
);

NAND2xp33_ASAP7_75t_R g2254 ( 
.A(n_2202),
.B(n_1905),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_SL g2255 ( 
.A(n_2199),
.B(n_2124),
.Y(n_2255)
);

AOI22xp5_ASAP7_75t_L g2256 ( 
.A1(n_2207),
.A2(n_2075),
.B1(n_2117),
.B2(n_2130),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2207),
.B(n_2091),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2190),
.B(n_2092),
.Y(n_2258)
);

NOR2xp33_ASAP7_75t_L g2259 ( 
.A(n_2209),
.B(n_2108),
.Y(n_2259)
);

INVxp67_ASAP7_75t_L g2260 ( 
.A(n_2224),
.Y(n_2260)
);

OAI221xp5_ASAP7_75t_L g2261 ( 
.A1(n_2238),
.A2(n_2208),
.B1(n_2202),
.B2(n_2224),
.C(n_2205),
.Y(n_2261)
);

NOR2x1_ASAP7_75t_L g2262 ( 
.A(n_2237),
.B(n_2202),
.Y(n_2262)
);

AOI221xp5_ASAP7_75t_L g2263 ( 
.A1(n_2231),
.A2(n_2205),
.B1(n_2208),
.B2(n_2203),
.C(n_2210),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2239),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2246),
.Y(n_2265)
);

INVx2_ASAP7_75t_SL g2266 ( 
.A(n_2233),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2257),
.B(n_2190),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_2247),
.B(n_2217),
.Y(n_2268)
);

HB1xp67_ASAP7_75t_L g2269 ( 
.A(n_2260),
.Y(n_2269)
);

BUFx2_ASAP7_75t_L g2270 ( 
.A(n_2249),
.Y(n_2270)
);

AOI22xp33_ASAP7_75t_L g2271 ( 
.A1(n_2231),
.A2(n_2202),
.B1(n_2223),
.B2(n_2200),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2232),
.B(n_2197),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2258),
.Y(n_2273)
);

INVxp67_ASAP7_75t_SL g2274 ( 
.A(n_2235),
.Y(n_2274)
);

NOR3xp33_ASAP7_75t_SL g2275 ( 
.A(n_2242),
.B(n_2210),
.C(n_2215),
.Y(n_2275)
);

INVxp67_ASAP7_75t_SL g2276 ( 
.A(n_2235),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2250),
.Y(n_2277)
);

INVx2_ASAP7_75t_SL g2278 ( 
.A(n_2236),
.Y(n_2278)
);

OAI22xp33_ASAP7_75t_L g2279 ( 
.A1(n_2240),
.A2(n_2217),
.B1(n_2082),
.B2(n_2124),
.Y(n_2279)
);

AOI21xp5_ASAP7_75t_L g2280 ( 
.A1(n_2242),
.A2(n_2220),
.B(n_2198),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2248),
.Y(n_2281)
);

AND2x4_ASAP7_75t_L g2282 ( 
.A(n_2244),
.B(n_2197),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_2241),
.B(n_2198),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2274),
.B(n_2245),
.Y(n_2284)
);

INVxp33_ASAP7_75t_L g2285 ( 
.A(n_2275),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2268),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_2268),
.Y(n_2287)
);

AOI21xp5_ASAP7_75t_L g2288 ( 
.A1(n_2276),
.A2(n_2234),
.B(n_2255),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2270),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2270),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2269),
.B(n_2252),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2278),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2282),
.B(n_2200),
.Y(n_2293)
);

OR2x2_ASAP7_75t_L g2294 ( 
.A(n_2272),
.B(n_2243),
.Y(n_2294)
);

AOI221xp5_ASAP7_75t_L g2295 ( 
.A1(n_2263),
.A2(n_2259),
.B1(n_2253),
.B2(n_2256),
.C(n_2130),
.Y(n_2295)
);

OAI321xp33_ASAP7_75t_L g2296 ( 
.A1(n_2261),
.A2(n_2259),
.A3(n_2253),
.B1(n_2251),
.B2(n_2254),
.C(n_2124),
.Y(n_2296)
);

HAxp5_ASAP7_75t_SL g2297 ( 
.A(n_2281),
.B(n_2160),
.CON(n_2297),
.SN(n_2297)
);

OAI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_2266),
.A2(n_2098),
.B1(n_2113),
.B2(n_2130),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_2293),
.B(n_2282),
.Y(n_2299)
);

INVx1_ASAP7_75t_SL g2300 ( 
.A(n_2286),
.Y(n_2300)
);

AOI21xp33_ASAP7_75t_SL g2301 ( 
.A1(n_2285),
.A2(n_2266),
.B(n_2279),
.Y(n_2301)
);

AOI221xp5_ASAP7_75t_L g2302 ( 
.A1(n_2285),
.A2(n_2284),
.B1(n_2289),
.B2(n_2290),
.C(n_2286),
.Y(n_2302)
);

AOI222xp33_ASAP7_75t_L g2303 ( 
.A1(n_2296),
.A2(n_2262),
.B1(n_2283),
.B2(n_2271),
.C1(n_2265),
.C2(n_2264),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2292),
.Y(n_2304)
);

AOI21xp5_ASAP7_75t_L g2305 ( 
.A1(n_2288),
.A2(n_2280),
.B(n_2282),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2287),
.B(n_2278),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2287),
.Y(n_2307)
);

NOR2xp33_ASAP7_75t_SL g2308 ( 
.A(n_2291),
.B(n_2273),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2294),
.B(n_2273),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2295),
.B(n_2267),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2298),
.B(n_2267),
.Y(n_2311)
);

AOI321xp33_ASAP7_75t_L g2312 ( 
.A1(n_2302),
.A2(n_2297),
.A3(n_2277),
.B1(n_2298),
.B2(n_2130),
.C(n_2117),
.Y(n_2312)
);

OAI32xp33_ASAP7_75t_L g2313 ( 
.A1(n_2300),
.A2(n_2277),
.A3(n_2098),
.B1(n_2113),
.B2(n_2178),
.Y(n_2313)
);

XOR2xp5_ASAP7_75t_L g2314 ( 
.A(n_2310),
.B(n_1902),
.Y(n_2314)
);

NAND4xp75_ASAP7_75t_L g2315 ( 
.A(n_2302),
.B(n_2187),
.C(n_2181),
.D(n_2178),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2305),
.B(n_2092),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2299),
.B(n_2109),
.Y(n_2317)
);

OAI221xp5_ASAP7_75t_L g2318 ( 
.A1(n_2303),
.A2(n_2152),
.B1(n_2153),
.B2(n_2179),
.C(n_2187),
.Y(n_2318)
);

OAI221xp5_ASAP7_75t_L g2319 ( 
.A1(n_2308),
.A2(n_2179),
.B1(n_2153),
.B2(n_2152),
.C(n_2181),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2306),
.Y(n_2320)
);

AOI21xp33_ASAP7_75t_SL g2321 ( 
.A1(n_2311),
.A2(n_2113),
.B(n_2130),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2307),
.Y(n_2322)
);

INVxp67_ASAP7_75t_L g2323 ( 
.A(n_2316),
.Y(n_2323)
);

OAI211xp5_ASAP7_75t_L g2324 ( 
.A1(n_2312),
.A2(n_2301),
.B(n_2304),
.C(n_2309),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2317),
.B(n_2109),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2322),
.B(n_2109),
.Y(n_2326)
);

OAI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_2314),
.A2(n_2117),
.B1(n_2112),
.B2(n_2177),
.Y(n_2327)
);

NAND3xp33_ASAP7_75t_SL g2328 ( 
.A(n_2312),
.B(n_1886),
.C(n_1839),
.Y(n_2328)
);

NAND5xp2_ASAP7_75t_SL g2329 ( 
.A(n_2318),
.B(n_2319),
.C(n_2315),
.D(n_2321),
.E(n_2313),
.Y(n_2329)
);

OAI22xp5_ASAP7_75t_L g2330 ( 
.A1(n_2320),
.A2(n_2117),
.B1(n_2112),
.B2(n_2116),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2326),
.Y(n_2331)
);

NOR2x1_ASAP7_75t_L g2332 ( 
.A(n_2324),
.B(n_2112),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2325),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2323),
.Y(n_2334)
);

NAND4xp75_ASAP7_75t_L g2335 ( 
.A(n_2329),
.B(n_2115),
.C(n_2114),
.D(n_2123),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2328),
.Y(n_2336)
);

OR2x2_ASAP7_75t_L g2337 ( 
.A(n_2333),
.B(n_2327),
.Y(n_2337)
);

NOR4xp75_ASAP7_75t_L g2338 ( 
.A(n_2335),
.B(n_2330),
.C(n_2116),
.D(n_2051),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2332),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2336),
.B(n_2134),
.Y(n_2340)
);

XNOR2xp5_ASAP7_75t_L g2341 ( 
.A(n_2338),
.B(n_2334),
.Y(n_2341)
);

AND2x4_ASAP7_75t_L g2342 ( 
.A(n_2341),
.B(n_2339),
.Y(n_2342)
);

OAI22xp5_ASAP7_75t_SL g2343 ( 
.A1(n_2342),
.A2(n_2331),
.B1(n_2337),
.B2(n_2340),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2342),
.Y(n_2344)
);

OAI22xp5_ASAP7_75t_SL g2345 ( 
.A1(n_2343),
.A2(n_2331),
.B1(n_1886),
.B2(n_2112),
.Y(n_2345)
);

OAI22xp5_ASAP7_75t_SL g2346 ( 
.A1(n_2344),
.A2(n_1886),
.B1(n_2112),
.B2(n_1789),
.Y(n_2346)
);

BUFx2_ASAP7_75t_L g2347 ( 
.A(n_2345),
.Y(n_2347)
);

OAI21x1_ASAP7_75t_SL g2348 ( 
.A1(n_2346),
.A2(n_2100),
.B(n_2093),
.Y(n_2348)
);

OAI21xp5_ASAP7_75t_L g2349 ( 
.A1(n_2347),
.A2(n_2112),
.B(n_2106),
.Y(n_2349)
);

AOI21xp5_ASAP7_75t_L g2350 ( 
.A1(n_2349),
.A2(n_2348),
.B(n_2097),
.Y(n_2350)
);

OAI22xp33_ASAP7_75t_L g2351 ( 
.A1(n_2350),
.A2(n_2093),
.B1(n_2097),
.B2(n_2118),
.Y(n_2351)
);

OAI221xp5_ASAP7_75t_R g2352 ( 
.A1(n_2351),
.A2(n_2097),
.B1(n_2093),
.B2(n_2100),
.C(n_2118),
.Y(n_2352)
);

AOI211xp5_ASAP7_75t_L g2353 ( 
.A1(n_2352),
.A2(n_1770),
.B(n_1869),
.C(n_1847),
.Y(n_2353)
);


endmodule