module real_jpeg_15503_n_20 (n_17, n_8, n_0, n_648, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_648;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_599;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_586;
wire n_155;
wire n_120;
wire n_405;
wire n_572;
wire n_412;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_602;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_636;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_597;
wire n_42;
wire n_313;
wire n_268;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_0),
.A2(n_21),
.B(n_644),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_0),
.B(n_645),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_1),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_1),
.Y(n_175)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_1),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g556 ( 
.A(n_1),
.Y(n_556)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_2),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_3),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_3),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_3),
.A2(n_256),
.B1(n_276),
.B2(n_279),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_3),
.A2(n_256),
.B1(n_330),
.B2(n_336),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_3),
.A2(n_256),
.B1(n_406),
.B2(n_407),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_4),
.A2(n_130),
.B1(n_187),
.B2(n_190),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_4),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_4),
.A2(n_190),
.B1(n_290),
.B2(n_294),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_4),
.A2(n_190),
.B1(n_463),
.B2(n_468),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_SL g522 ( 
.A1(n_4),
.A2(n_190),
.B1(n_523),
.B2(n_528),
.Y(n_522)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_5),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_5),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_5),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g510 ( 
.A(n_5),
.Y(n_510)
);

AOI22x1_ASAP7_75t_L g64 ( 
.A1(n_6),
.A2(n_65),
.B1(n_68),
.B2(n_70),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_6),
.A2(n_70),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_6),
.A2(n_70),
.B1(n_245),
.B2(n_396),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_6),
.A2(n_70),
.B1(n_603),
.B2(n_606),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_7),
.A2(n_52),
.B1(n_58),
.B2(n_61),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_7),
.A2(n_61),
.B1(n_155),
.B2(n_197),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_7),
.A2(n_61),
.B1(n_351),
.B2(n_356),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_7),
.A2(n_61),
.B1(n_590),
.B2(n_593),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_8),
.A2(n_178),
.B1(n_179),
.B2(n_182),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_8),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_8),
.A2(n_178),
.B1(n_322),
.B2(n_325),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_8),
.A2(n_178),
.B1(n_457),
.B2(n_461),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_8),
.A2(n_178),
.B1(n_541),
.B2(n_545),
.Y(n_544)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_9),
.A2(n_84),
.B1(n_88),
.B2(n_89),
.Y(n_83)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_9),
.A2(n_88),
.B1(n_270),
.B2(n_273),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_9),
.A2(n_88),
.B1(n_396),
.B2(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_9),
.A2(n_88),
.B1(n_474),
.B2(n_475),
.Y(n_473)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_10),
.Y(n_151)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_10),
.Y(n_158)
);

BUFx4f_ASAP7_75t_L g210 ( 
.A(n_10),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_10),
.Y(n_527)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_11),
.A2(n_154),
.B1(n_159),
.B2(n_160),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_11),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_11),
.A2(n_159),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_11),
.A2(n_159),
.B1(n_368),
.B2(n_370),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g583 ( 
.A1(n_11),
.A2(n_159),
.B1(n_584),
.B2(n_586),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_12),
.A2(n_165),
.B1(n_170),
.B2(n_172),
.Y(n_164)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_12),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_12),
.A2(n_172),
.B1(n_227),
.B2(n_230),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_12),
.A2(n_172),
.B1(n_385),
.B2(n_388),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_SL g598 ( 
.A1(n_12),
.A2(n_53),
.B1(n_172),
.B2(n_599),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_13),
.Y(n_99)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_13),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_14),
.A2(n_116),
.B1(n_121),
.B2(n_122),
.Y(n_115)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_14),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_14),
.A2(n_121),
.B1(n_306),
.B2(n_309),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_14),
.A2(n_55),
.B1(n_121),
.B2(n_182),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_14),
.A2(n_121),
.B1(n_443),
.B2(n_445),
.Y(n_442)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_15),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_15),
.B(n_63),
.Y(n_339)
);

OAI32xp33_ASAP7_75t_L g431 ( 
.A1(n_15),
.A2(n_101),
.A3(n_136),
.B1(n_432),
.B2(n_435),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_15),
.B(n_125),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_SL g489 ( 
.A1(n_15),
.A2(n_129),
.B1(n_490),
.B2(n_491),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_15),
.A2(n_144),
.B1(n_544),
.B2(n_551),
.Y(n_543)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_16),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_17),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_17),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_17),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_17),
.Y(n_249)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_17),
.Y(n_261)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_17),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_17),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g189 ( 
.A(n_19),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g587 ( 
.A(n_19),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_74),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_73),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_71),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_24),
.B(n_71),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_24),
.B(n_636),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_24),
.B(n_636),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_51),
.B1(n_62),
.B2(n_64),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_25),
.A2(n_62),
.B1(n_186),
.B2(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_25),
.A2(n_62),
.B1(n_269),
.B2(n_365),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_25),
.A2(n_62),
.B1(n_365),
.B2(n_405),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_25),
.A2(n_62),
.B1(n_405),
.B2(n_583),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_25),
.A2(n_51),
.B1(n_62),
.B2(n_629),
.Y(n_628)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_26),
.A2(n_63),
.B(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_26),
.A2(n_63),
.B1(n_177),
.B2(n_185),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_26),
.A2(n_63),
.B1(n_177),
.B2(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_26),
.A2(n_63),
.B1(n_597),
.B2(n_598),
.Y(n_596)
);

OA21x2_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_39),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_32),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_32),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_33),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_35),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

AOI22x1_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_43),
.B1(n_46),
.B2(n_50),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_44),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_45),
.Y(n_137)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_45),
.Y(n_278)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_45),
.Y(n_392)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_45),
.Y(n_493)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_48),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_49),
.Y(n_120)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_49),
.Y(n_293)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_57),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_57),
.Y(n_408)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_57),
.Y(n_585)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_69),
.Y(n_406)
);

AO21x1_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_574),
.B(n_637),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_413),
.B(n_569),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_343),
.C(n_376),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_281),
.B(n_313),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_78),
.B(n_281),
.C(n_571),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_191),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_79),
.B(n_192),
.C(n_250),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_126),
.C(n_176),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_81),
.B(n_176),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_94),
.B1(n_115),
.B2(n_124),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_83),
.A2(n_125),
.B1(n_289),
.B2(n_301),
.Y(n_288)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_87),
.Y(n_327)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_91),
.Y(n_593)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_93),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_94),
.A2(n_115),
.B1(n_124),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_94),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_94),
.A2(n_124),
.B1(n_275),
.B2(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_94),
.A2(n_124),
.B1(n_321),
.B2(n_489),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_94),
.A2(n_124),
.B1(n_384),
.B2(n_589),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_94),
.A2(n_124),
.B1(n_589),
.B2(n_602),
.Y(n_601)
);

AO21x1_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_101),
.B(n_107),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_108),
.B1(n_110),
.B2(n_112),
.Y(n_107)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_104),
.Y(n_387)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_105),
.Y(n_369)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_106),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_108),
.Y(n_255)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_108),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx6_ASAP7_75t_L g355 ( 
.A(n_109),
.Y(n_355)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_109),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_111),
.Y(n_229)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_111),
.Y(n_434)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_120),
.Y(n_592)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_125),
.A2(n_289),
.B1(n_301),
.B2(n_320),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_125),
.A2(n_301),
.B1(n_382),
.B2(n_383),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g626 ( 
.A1(n_125),
.A2(n_301),
.B(n_627),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_126),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_143),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_127),
.B(n_143),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_133),
.B1(n_138),
.B2(n_142),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_SL g303 ( 
.A1(n_128),
.A2(n_129),
.B(n_273),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_129),
.B(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_129),
.B(n_504),
.Y(n_503)
);

OAI21xp33_ASAP7_75t_SL g514 ( 
.A1(n_129),
.A2(n_503),
.B(n_515),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_129),
.B(n_173),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_R g557 ( 
.A(n_129),
.B(n_214),
.Y(n_557)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx6_ASAP7_75t_L g606 ( 
.A(n_136),
.Y(n_606)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_152),
.B1(n_164),
.B2(n_173),
.Y(n_143)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_144),
.A2(n_164),
.B1(n_196),
.B2(n_263),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_144),
.A2(n_206),
.B(n_360),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_144),
.A2(n_473),
.B1(n_476),
.B2(n_480),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_144),
.A2(n_522),
.B1(n_544),
.B2(n_554),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_150),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_145),
.A2(n_194),
.B1(n_329),
.B2(n_442),
.Y(n_441)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_148),
.Y(n_266)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_151),
.Y(n_219)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_151),
.Y(n_541)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_153),
.A2(n_194),
.B1(n_329),
.B2(n_337),
.Y(n_328)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_154),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_157),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_158),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_170),
.Y(n_207)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_174),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_175),
.Y(n_479)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g273 ( 
.A(n_189),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_250),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_211),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_193),
.A2(n_212),
.B(n_234),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_200),
.B2(n_205),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_194),
.A2(n_521),
.B1(n_530),
.B2(n_532),
.Y(n_520)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_204),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_209),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_234),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_225),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_213),
.A2(n_235),
.B1(n_305),
.B2(n_312),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_213),
.A2(n_235),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_213),
.A2(n_235),
.B1(n_456),
.B2(n_462),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_213),
.A2(n_235),
.B1(n_423),
.B2(n_462),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_213),
.A2(n_235),
.B1(n_456),
.B2(n_514),
.Y(n_513)
);

OA21x2_ASAP7_75t_L g580 ( 
.A1(n_213),
.A2(n_235),
.B(n_395),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_214),
.A2(n_244),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_214),
.A2(n_226),
.B1(n_253),
.B2(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_214),
.A2(n_253),
.B1(n_422),
.B2(n_428),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_219),
.B1(n_220),
.B2(n_222),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_221),
.Y(n_444)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_229),
.Y(n_233)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_243),
.Y(n_234)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g242 ( 
.A(n_238),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_238),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_241),
.Y(n_502)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_267),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_251),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_262),
.Y(n_251)
);

XOR2x2_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_262),
.Y(n_285)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_261),
.Y(n_311)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_261),
.Y(n_439)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_261),
.Y(n_506)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_265),
.Y(n_264)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_274),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_268),
.B(n_274),
.C(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_273),
.Y(n_599)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.C(n_286),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_282),
.A2(n_283),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_285),
.B(n_287),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_302),
.C(n_304),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_304),
.Y(n_316)
);

INVx8_ASAP7_75t_L g490 ( 
.A(n_290),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_293),
.Y(n_373)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_316),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_305),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_308),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_340),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_314),
.B(n_340),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_317),
.C(n_318),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_315),
.B(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_317),
.B(n_318),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_328),
.C(n_339),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_319),
.B(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_SL g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_328),
.B(n_339),
.Y(n_420)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_334),
.Y(n_474)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_335),
.Y(n_475)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_337),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx6_ASAP7_75t_L g531 ( 
.A(n_338),
.Y(n_531)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_341),
.Y(n_342)
);

A2O1A1O1Ixp25_ASAP7_75t_L g569 ( 
.A1(n_343),
.A2(n_376),
.B(n_570),
.C(n_572),
.D(n_573),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_375),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_SL g572 ( 
.A(n_344),
.B(n_375),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_347),
.Y(n_344)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_362),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_348),
.B(n_411),
.C(n_412),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_349),
.A2(n_358),
.B1(n_359),
.B2(n_361),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g361 ( 
.A(n_349),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_349),
.B(n_359),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_350),
.Y(n_394)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_354),
.Y(n_501)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_355),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_358),
.A2(n_359),
.B1(n_403),
.B2(n_404),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_358),
.A2(n_409),
.B1(n_615),
.B2(n_648),
.Y(n_614)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_362),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_374),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_366),
.C(n_374),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_367),
.Y(n_382)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_410),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_377),
.B(n_410),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_378),
.B(n_618),
.C(n_619),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_399),
.Y(n_379)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_380),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_381),
.A2(n_393),
.B(n_398),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_393),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_398),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_398),
.A2(n_610),
.B1(n_613),
.B2(n_622),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_399),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_400),
.A2(n_401),
.B1(n_402),
.B2(n_409),
.Y(n_399)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_400),
.Y(n_409)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_403),
.Y(n_615)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx3_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

AOI21x1_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_450),
.B(n_568),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_417),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_415),
.B(n_417),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_421),
.C(n_429),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g563 ( 
.A(n_419),
.B(n_564),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_421),
.A2(n_429),
.B1(n_430),
.B2(n_565),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_421),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_440),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_431),
.A2(n_440),
.B1(n_441),
.B2(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_431),
.Y(n_485)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_442),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_562),
.B(n_567),
.Y(n_450)
);

AOI21x1_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_496),
.B(n_561),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_483),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_453),
.B(n_483),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_472),
.C(n_481),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_454),
.A2(n_455),
.B1(n_481),
.B2(n_482),
.Y(n_517)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_470),
.Y(n_515)
);

INVx5_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_472),
.B(n_517),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_473),
.Y(n_532)
);

OAI32xp33_ASAP7_75t_L g499 ( 
.A1(n_475),
.A2(n_500),
.A3(n_502),
.B1(n_503),
.B2(n_507),
.Y(n_499)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_475),
.Y(n_511)
);

BUFx5_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_486),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_484),
.B(n_487),
.C(n_495),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_487),
.A2(n_488),
.B1(n_494),
.B2(n_495),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_497),
.A2(n_518),
.B(n_560),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_516),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_498),
.B(n_516),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_512),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_499),
.A2(n_512),
.B1(n_513),
.B2(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_499),
.Y(n_534)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_511),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_519),
.A2(n_535),
.B(n_559),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_533),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_520),
.B(n_533),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_527),
.Y(n_550)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_529),
.Y(n_528)
);

INVx6_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_536),
.A2(n_552),
.B(n_558),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_543),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_542),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_539),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_553),
.B(n_557),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_553),
.B(n_557),
.Y(n_558)
);

INVx6_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

BUFx12f_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

NOR2xp67_ASAP7_75t_SL g562 ( 
.A(n_563),
.B(n_566),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_563),
.B(n_566),
.Y(n_567)
);

NOR3xp33_ASAP7_75t_L g574 ( 
.A(n_575),
.B(n_623),
.C(n_634),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_576),
.B(n_616),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_577),
.A2(n_640),
.B(n_641),
.Y(n_639)
);

NOR2x1_ASAP7_75t_L g577 ( 
.A(n_578),
.B(n_608),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_578),
.B(n_608),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_579),
.B(n_594),
.Y(n_578)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_579),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_580),
.B(n_581),
.C(n_588),
.Y(n_579)
);

XNOR2x1_ASAP7_75t_L g600 ( 
.A(n_580),
.B(n_601),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_580),
.B(n_588),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_580),
.B(n_596),
.C(n_631),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_581),
.A2(n_582),
.B1(n_595),
.B2(n_607),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_581),
.A2(n_582),
.B1(n_611),
.B2(n_612),
.Y(n_610)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_582),
.B(n_595),
.C(n_633),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_583),
.Y(n_597)
);

INVx6_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_595),
.Y(n_607)
);

XNOR2x1_ASAP7_75t_L g595 ( 
.A(n_596),
.B(n_600),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g629 ( 
.A(n_598),
.Y(n_629)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_601),
.Y(n_631)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_602),
.Y(n_627)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_609),
.B(n_613),
.C(n_614),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_610),
.Y(n_622)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_611),
.Y(n_612)
);

XOR2xp5_ASAP7_75t_L g620 ( 
.A(n_614),
.B(n_621),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_617),
.B(n_620),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_617),
.B(n_620),
.Y(n_640)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_624),
.Y(n_623)
);

A2O1A1O1Ixp25_ASAP7_75t_L g638 ( 
.A1(n_624),
.A2(n_635),
.B(n_639),
.C(n_642),
.D(n_643),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_625),
.B(n_632),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_625),
.B(n_632),
.Y(n_642)
);

BUFx24_ASAP7_75t_SL g646 ( 
.A(n_625),
.Y(n_646)
);

FAx1_ASAP7_75t_SL g625 ( 
.A(n_626),
.B(n_628),
.CI(n_630),
.CON(n_625),
.SN(n_625)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_626),
.B(n_628),
.C(n_630),
.Y(n_636)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_635),
.Y(n_634)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);


endmodule