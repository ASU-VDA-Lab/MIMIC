module fake_jpeg_6299_n_301 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NAND2x1_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_0),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_37),
.B(n_24),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_39),
.Y(n_47)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_57),
.Y(n_86)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_23),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_54),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_19),
.B1(n_32),
.B2(n_18),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_55),
.B1(n_64),
.B2(n_66),
.Y(n_68)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_53),
.B(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_30),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_19),
.B1(n_32),
.B2(n_18),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_19),
.B1(n_34),
.B2(n_21),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_33),
.B1(n_17),
.B2(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_62),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_34),
.C(n_21),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_42),
.C(n_40),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_23),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_28),
.B1(n_31),
.B2(n_18),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_38),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_27),
.B1(n_30),
.B2(n_23),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_33),
.B1(n_17),
.B2(n_29),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_42),
.B1(n_40),
.B2(n_37),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_80),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_31),
.B1(n_41),
.B2(n_27),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_29),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_41),
.B1(n_26),
.B2(n_37),
.Y(n_73)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_78),
.Y(n_95)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_42),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_85),
.B(n_54),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_45),
.A2(n_41),
.B1(n_26),
.B2(n_37),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_33),
.A3(n_17),
.B1(n_24),
.B2(n_43),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_64),
.C(n_29),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_82),
.B(n_83),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_24),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_45),
.A2(n_33),
.B1(n_17),
.B2(n_14),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_90),
.B1(n_73),
.B2(n_80),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_52),
.B(n_0),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_17),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_93),
.Y(n_115)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_0),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_47),
.C(n_51),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_102),
.C(n_93),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_116),
.B1(n_106),
.B2(n_99),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_55),
.C(n_50),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_104),
.B(n_107),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_45),
.B1(n_56),
.B2(n_66),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_68),
.B1(n_89),
.B2(n_71),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_74),
.B(n_63),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_118),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_49),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_110),
.B(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_67),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_113),
.B(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_65),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_79),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_48),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_57),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_121),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_83),
.B(n_0),
.Y(n_121)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_130),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_129),
.B1(n_131),
.B2(n_149),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_68),
.B1(n_70),
.B2(n_89),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_106),
.A2(n_89),
.B1(n_75),
.B2(n_72),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_132),
.B(n_137),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_133),
.A2(n_58),
.B1(n_77),
.B2(n_101),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_102),
.A2(n_75),
.B(n_69),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_134),
.A2(n_121),
.B(n_105),
.Y(n_162)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_108),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_142),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_140),
.C(n_143),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_75),
.C(n_72),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_117),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_94),
.C(n_87),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_144),
.B(n_11),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_88),
.B1(n_78),
.B2(n_85),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_111),
.B1(n_120),
.B2(n_118),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_78),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_107),
.B(n_1),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_110),
.B(n_114),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_106),
.A2(n_84),
.B1(n_65),
.B2(n_58),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_111),
.Y(n_150)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_155),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_102),
.C(n_119),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_162),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_156),
.A2(n_173),
.B1(n_176),
.B2(n_180),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_148),
.A2(n_126),
.B1(n_103),
.B2(n_109),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_158),
.Y(n_182)
);

NOR3xp33_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_104),
.C(n_113),
.Y(n_160)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_141),
.C(n_123),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_99),
.B1(n_97),
.B2(n_119),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_161),
.A2(n_172),
.B1(n_140),
.B2(n_135),
.Y(n_192)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_167),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_105),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_154),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_148),
.A2(n_109),
.B1(n_58),
.B2(n_77),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_174),
.B(n_132),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_145),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_171),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_129),
.B1(n_131),
.B2(n_143),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_98),
.B(n_92),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_60),
.B1(n_43),
.B2(n_98),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_178),
.Y(n_200)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_179),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_122),
.A2(n_43),
.B1(n_98),
.B2(n_29),
.Y(n_180)
);

NAND5xp2_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_163),
.C(n_161),
.D(n_171),
.E(n_159),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_183),
.B(n_192),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_189),
.B(n_197),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_134),
.B(n_122),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_202),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_198),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_123),
.B1(n_141),
.B2(n_135),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_174),
.B1(n_169),
.B2(n_155),
.Y(n_219)
);

BUFx12f_ASAP7_75t_SL g197 ( 
.A(n_160),
.Y(n_197)
);

NOR3xp33_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_147),
.C(n_137),
.Y(n_199)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

NAND2xp33_ASAP7_75t_SL g201 ( 
.A(n_153),
.B(n_124),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_206),
.B(n_3),
.Y(n_225)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_151),
.B(n_128),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_151),
.C(n_157),
.Y(n_212)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_180),
.Y(n_220)
);

AO22x1_ASAP7_75t_L g206 ( 
.A1(n_173),
.A2(n_128),
.B1(n_124),
.B2(n_43),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_191),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_208),
.Y(n_236)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_216),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_215),
.C(n_218),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_204),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_214),
.B(n_4),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_159),
.C(n_165),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_177),
.B1(n_175),
.B2(n_157),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_222),
.B1(n_226),
.B2(n_206),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_167),
.C(n_156),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_219),
.B(n_185),
.Y(n_240)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_176),
.C(n_178),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_223),
.C(n_12),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_182),
.A2(n_136),
.B1(n_2),
.B2(n_3),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_1),
.C(n_2),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_1),
.Y(n_224)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_229),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_183),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_186),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_248),
.C(n_221),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_227),
.A2(n_181),
.B1(n_196),
.B2(n_197),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_237),
.B1(n_219),
.B2(n_209),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_181),
.B1(n_201),
.B2(n_188),
.Y(n_237)
);

OAI22x1_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_184),
.B1(n_185),
.B2(n_195),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_238),
.A2(n_229),
.B1(n_216),
.B2(n_220),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_245),
.Y(n_249)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_243),
.B(n_246),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_227),
.B(n_11),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_224),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_254),
.B(n_238),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_256),
.C(n_261),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_232),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_212),
.C(n_218),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_233),
.A2(n_211),
.B1(n_228),
.B2(n_223),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_240),
.B1(n_245),
.B2(n_4),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_211),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_259),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_228),
.C(n_213),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_248),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_236),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_263),
.B(n_265),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_231),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_273),
.C(n_251),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_241),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_269),
.B(n_270),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_241),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_268),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_230),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_233),
.B(n_235),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_271),
.A2(n_10),
.B(n_15),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_272),
.A2(n_254),
.B1(n_249),
.B2(n_261),
.Y(n_275)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_282),
.C(n_274),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_269),
.A2(n_256),
.B1(n_257),
.B2(n_249),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_278),
.B(n_276),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_266),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_284),
.Y(n_288)
);

NOR2xp67_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_260),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_7),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_270),
.A2(n_10),
.B1(n_15),
.B2(n_7),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_277),
.B(n_274),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_287),
.B(n_291),
.Y(n_293)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_281),
.A3(n_279),
.B1(n_9),
.B2(n_13),
.C1(n_14),
.C2(n_16),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_9),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_283),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_295),
.B1(n_296),
.B2(n_4),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_294),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_283),
.B1(n_278),
.B2(n_9),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_288),
.A2(n_13),
.B(n_16),
.Y(n_296)
);

AOI321xp33_ASAP7_75t_L g299 ( 
.A1(n_297),
.A2(n_6),
.A3(n_285),
.B1(n_293),
.B2(n_199),
.C(n_76),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_298),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_6),
.Y(n_301)
);


endmodule