module real_jpeg_16952_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_8),
.B1(n_15),
.B2(n_16),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

AND2x4_ASAP7_75t_L g35 ( 
.A(n_1),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_1),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_1),
.B(n_62),
.Y(n_61)
);

AND2x4_ASAP7_75t_SL g73 ( 
.A(n_1),
.B(n_74),
.Y(n_73)
);

AND2x4_ASAP7_75t_L g99 ( 
.A(n_1),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_1),
.B(n_56),
.Y(n_117)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_1),
.Y(n_140)
);

NAND2x1p5_ASAP7_75t_L g181 ( 
.A(n_1),
.B(n_182),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_2),
.Y(n_323)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_3),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_4),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_4),
.B(n_224),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_4),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_4),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_4),
.B(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_5),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_5),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_6),
.B(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_6),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_6),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_6),
.B(n_40),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_6),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_6),
.B(n_182),
.Y(n_241)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_7),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_9),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_9),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_9),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_9),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_9),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_9),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_9),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_9),
.B(n_220),
.Y(n_219)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_10),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_10),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_11),
.Y(n_137)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_12),
.Y(n_87)
);

BUFx4f_ASAP7_75t_L g226 ( 
.A(n_12),
.Y(n_226)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_13),
.Y(n_182)
);

BUFx8_ASAP7_75t_L g220 ( 
.A(n_13),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_302),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_270),
.B(n_300),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_232),
.B(n_264),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_197),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_159),
.B(n_196),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_126),
.B(n_158),
.Y(n_22)
);

OAI21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_96),
.B(n_125),
.Y(n_23)
);

NOR2xp67_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_78),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_25),
.B(n_78),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_57),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_42),
.B2(n_43),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_27),
.B(n_43),
.C(n_57),
.Y(n_127)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.B1(n_34),
.B2(n_41),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_29),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_29),
.B(n_35),
.C(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_29),
.B(n_45),
.C(n_170),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_29),
.A2(n_41),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_35),
.A2(n_256),
.B1(n_257),
.B2(n_259),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_35),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_35),
.B(n_257),
.C(n_260),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_35),
.B(n_218),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_35),
.A2(n_180),
.B1(n_181),
.B2(n_256),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_38),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_38),
.A2(n_155),
.B1(n_169),
.B2(n_175),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_41),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.C(n_53),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_44),
.A2(n_45),
.B1(n_53),
.B2(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_44),
.A2(n_45),
.B1(n_170),
.B2(n_174),
.Y(n_248)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_45),
.B(n_209),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g244 ( 
.A1(n_45),
.A2(n_245),
.B(n_246),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_49),
.B1(n_80),
.B2(n_82),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_48),
.A2(n_49),
.B1(n_148),
.B2(n_151),
.Y(n_147)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_49),
.A2(n_108),
.B(n_117),
.C(n_149),
.Y(n_165)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_53),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_53),
.A2(n_81),
.B1(n_132),
.B2(n_144),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_53),
.B(n_293),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_90),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_54),
.B(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_69),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_59),
.A2(n_114),
.B(n_118),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_59),
.A2(n_70),
.B(n_77),
.Y(n_145)
);

NOR2x1_ASAP7_75t_R g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_60),
.A2(n_61),
.B1(n_88),
.B2(n_89),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_60),
.A2(n_61),
.B1(n_116),
.B2(n_117),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_60),
.B(n_73),
.C(n_139),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_73),
.B(n_75),
.Y(n_72)
);

NAND2x1p5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_73),
.Y(n_75)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_65),
.A2(n_103),
.B1(n_106),
.B2(n_107),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_72),
.B1(n_76),
.B2(n_77),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_99),
.B(n_102),
.C(n_108),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_99),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_70),
.A2(n_76),
.B1(n_99),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_72),
.A2(n_77),
.B1(n_138),
.B2(n_139),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_84),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_73),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_73),
.B(n_103),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_73),
.A2(n_94),
.B1(n_103),
.B2(n_106),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_73),
.A2(n_103),
.B(n_241),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_75),
.B(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_75),
.B(n_132),
.C(n_139),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.C(n_92),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_81),
.B(n_144),
.C(n_204),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_81),
.B(n_149),
.C(n_294),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_92),
.B1(n_93),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_83),
.A2(n_84),
.B(n_88),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_88),
.A2(n_89),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_89),
.B(n_219),
.C(n_223),
.Y(n_260)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_112),
.B(n_124),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_109),
.Y(n_97)
);

NOR2xp67_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_109),
.Y(n_124)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_99),
.B(n_116),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_99),
.B(n_117),
.C(n_181),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_99),
.A2(n_122),
.B1(n_208),
.B2(n_212),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_99),
.B(n_210),
.Y(n_246)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_103),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_103),
.A2(n_106),
.B1(n_170),
.B2(n_174),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_103),
.B(n_155),
.C(n_170),
.Y(n_229)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_120),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_119),
.B(n_123),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_116),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_116),
.A2(n_117),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_122),
.B(n_209),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_128),
.Y(n_158)
);

XOR2x2_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_146),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_145),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_130),
.B(n_145),
.C(n_146),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_138),
.B1(n_139),
.B2(n_144),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_136),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_138),
.A2(n_139),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_143),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_152),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_153),
.C(n_157),
.Y(n_162)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

AO22x1_ASAP7_75t_L g293 ( 
.A1(n_149),
.A2(n_150),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_195),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_195),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_176),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_163),
.C(n_176),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_168),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_166),
.B(n_168),
.C(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_167),
.B(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_194),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_184),
.C(n_194),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_183),
.Y(n_178)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_179),
.Y(n_183)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_191),
.B(n_193),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_191),
.Y(n_193)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_191),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_191),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_193),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_198),
.B(n_199),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_215),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_200),
.B(n_216),
.C(n_231),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_213),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_206),
.B2(n_207),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_206),
.C(n_213),
.Y(n_234)
);

XNOR2x2_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_208),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_231),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_227),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_229),
.C(n_230),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_218),
.B(n_256),
.C(n_280),
.Y(n_331)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_263),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_263),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_234),
.B(n_237),
.C(n_249),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_249),
.B2(n_250),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2x2_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_247),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_243),
.B2(n_244),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_239),
.B(n_244),
.C(n_247),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2x1_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_261),
.B2(n_262),
.Y(n_252)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_262),
.C(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_254),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_260),
.Y(n_254)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_299),
.Y(n_271)
);

NOR2x1_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_299),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_276),
.C(n_287),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_287),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_286),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_284),
.B2(n_285),
.Y(n_277)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_285),
.C(n_286),
.Y(n_307)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_290),
.C(n_292),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_332),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_306),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_325),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_314),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_324),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_331),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);


endmodule