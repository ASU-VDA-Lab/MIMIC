module fake_jpeg_11583_n_38 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_38);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

INVx3_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_20),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_0),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g21 ( 
.A1(n_16),
.A2(n_13),
.B1(n_12),
.B2(n_9),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_15),
.B1(n_14),
.B2(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_1),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_2),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_14),
.B(n_15),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.C(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_18),
.C(n_3),
.Y(n_31)
);

XOR2x2_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_8),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.C(n_31),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_24),
.B(n_4),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_34),
.Y(n_36)
);

INVxp33_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_35)
);

NAND5xp2_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_5),
.C(n_6),
.D(n_7),
.E(n_36),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_35),
.Y(n_38)
);


endmodule