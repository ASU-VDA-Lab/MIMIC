module fake_jpeg_24250_n_108 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVxp67_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVxp33_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_16),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx9p33_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_25),
.A2(n_13),
.B1(n_17),
.B2(n_16),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_13),
.B1(n_9),
.B2(n_18),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_13),
.B1(n_17),
.B2(n_15),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_28),
.B(n_21),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_25),
.B1(n_33),
.B2(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_44),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_43),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

AOI22x1_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_34),
.B1(n_27),
.B2(n_26),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_49),
.B1(n_41),
.B2(n_42),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_25),
.B1(n_33),
.B2(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_43),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_15),
.B1(n_14),
.B2(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_66),
.Y(n_75)
);

AOI221xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_62),
.B1(n_51),
.B2(n_49),
.C(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_43),
.C(n_39),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_52),
.C(n_14),
.Y(n_73)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_39),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_46),
.B1(n_48),
.B2(n_52),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_30),
.B1(n_10),
.B2(n_20),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_15),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_47),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_73),
.C(n_63),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_70),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_71),
.B1(n_76),
.B2(n_62),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_64),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_0),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_79),
.C(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_81),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_22),
.C(n_20),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_76),
.B1(n_22),
.B2(n_20),
.Y(n_89)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_87),
.C(n_83),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_79),
.B(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_16),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_94),
.C(n_95),
.Y(n_98)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_88),
.A2(n_7),
.B(n_8),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_7),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_22),
.C(n_20),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_22),
.C(n_16),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_86),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_99),
.B1(n_0),
.B2(n_2),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_6),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_99),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_101),
.B(n_102),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_103),
.Y(n_106)
);

AOI221xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_100),
.B1(n_5),
.B2(n_3),
.C(n_30),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_5),
.Y(n_108)
);


endmodule