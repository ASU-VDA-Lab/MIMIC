module fake_jpeg_588_n_105 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_105);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_43),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_32),
.C(n_36),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_34),
.C(n_29),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_37),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_49),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_53),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_31),
.B1(n_30),
.B2(n_37),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_44),
.B1(n_43),
.B2(n_11),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_50),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_45),
.B1(n_46),
.B2(n_43),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_26),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_1),
.C(n_2),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_66),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_51),
.B(n_48),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_70),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_19),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_17),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_54),
.B1(n_61),
.B2(n_59),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_80),
.B1(n_7),
.B2(n_8),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_83),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_18),
.C(n_16),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_70),
.C(n_12),
.Y(n_85)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_68),
.B1(n_8),
.B2(n_9),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_86),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_81),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_13),
.B1(n_15),
.B2(n_9),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_10),
.B1(n_78),
.B2(n_77),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

XNOR2x1_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_83),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_93),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_96),
.B(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_98),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_94),
.CI(n_85),
.CON(n_103),
.SN(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_10),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_103),
.Y(n_105)
);


endmodule