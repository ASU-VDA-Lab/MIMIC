module fake_jpeg_28753_n_451 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_451);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_451;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_48),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_51),
.Y(n_123)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

BUFx12f_ASAP7_75t_SL g55 ( 
.A(n_15),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g133 ( 
.A(n_55),
.Y(n_133)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_59),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_72),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_26),
.B(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_68),
.B(n_83),
.Y(n_92)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_26),
.B(n_7),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_79),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_80),
.Y(n_122)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_82),
.Y(n_127)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_85),
.Y(n_118)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_87),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_89),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_17),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_20),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g142 ( 
.A(n_95),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_49),
.B(n_40),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_104),
.B(n_110),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_52),
.A2(n_38),
.B1(n_22),
.B2(n_41),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_105),
.A2(n_107),
.B1(n_112),
.B2(n_95),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_63),
.A2(n_22),
.B1(n_17),
.B2(n_41),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_106),
.A2(n_129),
.B1(n_35),
.B2(n_61),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_76),
.A2(n_22),
.B1(n_41),
.B2(n_25),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g110 ( 
.A1(n_49),
.A2(n_45),
.B(n_44),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_25),
.B1(n_37),
.B2(n_29),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_33),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_130),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_85),
.A2(n_17),
.B1(n_28),
.B2(n_40),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_57),
.B(n_33),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_58),
.B(n_43),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_134),
.B(n_43),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_53),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_54),
.B(n_28),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_138),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_54),
.B(n_32),
.Y(n_138)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_151),
.Y(n_197)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_148),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_120),
.A2(n_71),
.B1(n_77),
.B2(n_87),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_149),
.A2(n_150),
.B1(n_179),
.B2(n_106),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_66),
.B1(n_86),
.B2(n_81),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_92),
.B(n_42),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_152),
.B(n_155),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_98),
.B(n_42),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_153),
.B(n_174),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_108),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_181),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_133),
.B(n_45),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_160),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_129),
.A2(n_35),
.B1(n_44),
.B2(n_80),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_158),
.B(n_163),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_159),
.A2(n_158),
.B1(n_151),
.B2(n_143),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_135),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_133),
.A2(n_88),
.B1(n_79),
.B2(n_74),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

OA22x2_ASAP7_75t_SL g164 ( 
.A1(n_108),
.A2(n_89),
.B1(n_72),
.B2(n_59),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_165),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_109),
.B(n_0),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_125),
.C(n_126),
.Y(n_206)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_122),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_173),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_118),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_102),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_180),
.Y(n_205)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_124),
.A2(n_89),
.B1(n_72),
.B2(n_59),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_127),
.B(n_140),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_116),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_182),
.A2(n_184),
.B1(n_185),
.B2(n_123),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_123),
.Y(n_199)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_SL g187 ( 
.A1(n_181),
.A2(n_128),
.B(n_100),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_199),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_188),
.A2(n_218),
.B1(n_142),
.B2(n_101),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_147),
.A2(n_127),
.B1(n_94),
.B2(n_116),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_193),
.A2(n_198),
.B1(n_211),
.B2(n_168),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_128),
.B1(n_93),
.B2(n_91),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_200),
.A2(n_220),
.B1(n_197),
.B2(n_216),
.Y(n_242)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_143),
.B(n_127),
.C(n_139),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_207),
.C(n_217),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_119),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_212),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_142),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_144),
.B(n_117),
.C(n_96),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_210),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_149),
.A2(n_93),
.B1(n_91),
.B2(n_115),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_96),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_146),
.B(n_154),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_164),
.A2(n_115),
.B1(n_101),
.B2(n_111),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_175),
.A2(n_111),
.B1(n_117),
.B2(n_46),
.Y(n_220)
);

INVx11_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_145),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_225),
.B(n_226),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_165),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_196),
.A2(n_159),
.B1(n_183),
.B2(n_150),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_227),
.A2(n_241),
.B1(n_252),
.B2(n_254),
.Y(n_260)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_228),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_195),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_229),
.B(n_236),
.Y(n_271)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_231),
.Y(n_284)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_234),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_146),
.B(n_164),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_235),
.A2(n_217),
.B(n_197),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_178),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_237),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_194),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_239),
.Y(n_272)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_244),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_242),
.A2(n_255),
.B1(n_141),
.B2(n_148),
.Y(n_286)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_247),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_248),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_179),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_246),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_189),
.B(n_156),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_191),
.B(n_169),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_199),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_257),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_201),
.Y(n_273)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_253),
.B(n_256),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_188),
.A2(n_176),
.B1(n_182),
.B2(n_180),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_185),
.B1(n_177),
.B2(n_172),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_189),
.B(n_202),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_203),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_191),
.A2(n_171),
.B1(n_173),
.B2(n_184),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_213),
.B1(n_186),
.B2(n_209),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_232),
.A2(n_235),
.B(n_249),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_259),
.A2(n_277),
.B(n_279),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_216),
.B1(n_222),
.B2(n_211),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_263),
.A2(n_286),
.B1(n_20),
.B2(n_9),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_268),
.A2(n_276),
.B(n_288),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_197),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_269),
.B(n_285),
.C(n_246),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_270),
.A2(n_255),
.B1(n_224),
.B2(n_228),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_273),
.B(n_280),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_229),
.A2(n_209),
.B1(n_213),
.B2(n_223),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_274),
.A2(n_275),
.B1(n_231),
.B2(n_245),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_238),
.A2(n_239),
.B1(n_230),
.B2(n_234),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_233),
.A2(n_212),
.B(n_207),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_232),
.A2(n_206),
.B(n_193),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_232),
.A2(n_113),
.B(n_132),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_251),
.B(n_205),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_132),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_242),
.A2(n_37),
.B(n_29),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_287),
.A2(n_289),
.B(n_246),
.Y(n_306)
);

MAJx3_ASAP7_75t_L g288 ( 
.A(n_233),
.B(n_20),
.C(n_37),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_247),
.A2(n_37),
.B(n_29),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_284),
.Y(n_292)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_292),
.Y(n_327)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_284),
.Y(n_293)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_290),
.B(n_262),
.Y(n_294)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_294),
.Y(n_339)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_264),
.Y(n_296)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_296),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_253),
.Y(n_297)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_264),
.Y(n_298)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_298),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_244),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_299),
.B(n_316),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_243),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_303),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_266),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_315),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_304),
.B(n_283),
.Y(n_346)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_265),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_305),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_306),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_260),
.A2(n_227),
.B1(n_254),
.B2(n_241),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_309),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_308),
.A2(n_312),
.B1(n_320),
.B2(n_321),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_260),
.A2(n_257),
.B1(n_258),
.B2(n_231),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_291),
.A2(n_240),
.B1(n_237),
.B2(n_20),
.Y(n_311)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_311),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_291),
.A2(n_37),
.B1(n_29),
.B2(n_20),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_278),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_313),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_314),
.A2(n_317),
.B1(n_289),
.B2(n_283),
.Y(n_344)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_278),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_271),
.B(n_18),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_263),
.A2(n_286),
.B1(n_268),
.B2(n_285),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_262),
.B(n_0),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_319),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_259),
.A2(n_279),
.B(n_276),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_277),
.A2(n_9),
.B(n_2),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_265),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_269),
.C(n_273),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_326),
.C(n_336),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_280),
.C(n_288),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_304),
.B(n_288),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_328),
.B(n_331),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_295),
.B(n_287),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_314),
.A2(n_272),
.B1(n_281),
.B2(n_270),
.Y(n_332)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_332),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_300),
.B(n_261),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_301),
.B(n_272),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_318),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_344),
.A2(n_307),
.B1(n_309),
.B2(n_303),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_346),
.B(n_347),
.C(n_348),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_300),
.B(n_18),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_18),
.C(n_1),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_297),
.Y(n_350)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_350),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_351),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_357),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_329),
.A2(n_317),
.B1(n_294),
.B2(n_302),
.Y(n_353)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_339),
.B(n_315),
.Y(n_354)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_354),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_336),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_369),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_320),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_327),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_358),
.B(n_359),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_313),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_323),
.B(n_295),
.C(n_306),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_361),
.C(n_362),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_298),
.C(n_296),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_311),
.C(n_312),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_329),
.A2(n_321),
.B1(n_293),
.B2(n_305),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_363),
.B(n_365),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_292),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_364),
.B(n_368),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_343),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_347),
.B(n_18),
.C(n_1),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_366),
.B(n_331),
.C(n_333),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_343),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_3),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_322),
.B(n_4),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_348),
.Y(n_381)
);

OA21x2_ASAP7_75t_L g375 ( 
.A1(n_371),
.A2(n_345),
.B(n_333),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_375),
.A2(n_385),
.B(n_388),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_381),
.B(n_4),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_383),
.B(n_356),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_344),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_384),
.B(n_387),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_359),
.A2(n_345),
.B(n_341),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_325),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_352),
.A2(n_341),
.B(n_334),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_355),
.B(n_360),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_389),
.B(n_390),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_334),
.C(n_324),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_391),
.B(n_401),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_356),
.C(n_367),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_395),
.C(n_396),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_367),
.C(n_362),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_389),
.C(n_387),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_382),
.B(n_374),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_397),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_373),
.A2(n_350),
.B(n_324),
.Y(n_398)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_398),
.Y(n_415)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_377),
.Y(n_399)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_399),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_390),
.B(n_380),
.C(n_379),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_400),
.B(n_403),
.C(n_5),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_378),
.B(n_358),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_388),
.A2(n_342),
.B(n_366),
.Y(n_402)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_402),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_368),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_405),
.B(n_381),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_404),
.A2(n_375),
.B(n_385),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_10),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_407),
.B(n_411),
.Y(n_420)
);

OAI321xp33_ASAP7_75t_L g410 ( 
.A1(n_397),
.A2(n_375),
.A3(n_372),
.B1(n_386),
.B2(n_379),
.C(n_11),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_410),
.A2(n_414),
.B1(n_5),
.B2(n_10),
.Y(n_423)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_404),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_400),
.B(n_4),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_412),
.B(n_419),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_403),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_416),
.B(n_393),
.C(n_392),
.Y(n_424)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_394),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_409),
.B(n_395),
.Y(n_421)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_421),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_416),
.B(n_394),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_422),
.B(n_429),
.Y(n_432)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_423),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_424),
.B(n_428),
.Y(n_433)
);

INVxp33_ASAP7_75t_L g425 ( 
.A(n_413),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_426),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_417),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_396),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_408),
.B(n_393),
.Y(n_429)
);

OAI21xp33_ASAP7_75t_L g434 ( 
.A1(n_430),
.A2(n_418),
.B(n_415),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_425),
.B(n_408),
.Y(n_431)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_431),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_434),
.A2(n_435),
.B(n_436),
.Y(n_443)
);

FAx1_ASAP7_75t_SL g437 ( 
.A(n_428),
.B(n_406),
.CI(n_414),
.CON(n_437),
.SN(n_437)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_437),
.B(n_420),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_439),
.B(n_441),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_433),
.A2(n_427),
.B(n_419),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_440),
.A2(n_443),
.B(n_438),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_433),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_442),
.A2(n_422),
.B(n_430),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_444),
.A2(n_446),
.B1(n_432),
.B2(n_407),
.Y(n_447)
);

NAND4xp25_ASAP7_75t_SL g448 ( 
.A(n_447),
.B(n_445),
.C(n_11),
.D(n_13),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_10),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_449),
.A2(n_13),
.B(n_14),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_450),
.B(n_18),
.Y(n_451)
);


endmodule