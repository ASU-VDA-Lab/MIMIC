module fake_netlist_6_612_n_1486 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_350, n_78, n_84, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_376, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_364, n_295, n_385, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1486);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_364;
input n_295;
input n_385;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1486;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_1094;
wire n_953;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_811;
wire n_683;
wire n_1207;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1483;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_1437;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_1037;
wire n_621;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_1485;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_1408;
wire n_1196;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1109;
wire n_712;
wire n_1276;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

INVx2_ASAP7_75t_L g388 ( 
.A(n_329),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_360),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_47),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_284),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_13),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_385),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_112),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_132),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_231),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_253),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_357),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_274),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_26),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_83),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_354),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_100),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_178),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_22),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_268),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_380),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_194),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_133),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_191),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_287),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_312),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_108),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_5),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_31),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_382),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_41),
.Y(n_418)
);

INVxp33_ASAP7_75t_R g419 ( 
.A(n_230),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_264),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_179),
.Y(n_421)
);

BUFx10_ASAP7_75t_L g422 ( 
.A(n_307),
.Y(n_422)
);

BUFx5_ASAP7_75t_L g423 ( 
.A(n_110),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_318),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_371),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_105),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_169),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_146),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_252),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_189),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_11),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_59),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_41),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_85),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_365),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_372),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_99),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_279),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_259),
.Y(n_439)
);

BUFx8_ASAP7_75t_SL g440 ( 
.A(n_321),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_376),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_286),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_153),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_340),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_75),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_149),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_87),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_9),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_320),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_317),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_54),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_134),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_55),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_277),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_229),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_347),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_366),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_313),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_322),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_197),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_293),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_20),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_350),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_63),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_204),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_225),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_294),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_209),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_222),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_251),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_155),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_124),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_260),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_59),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_160),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_78),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_128),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_1),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_301),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_364),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_68),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_343),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_182),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_205),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_131),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_82),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_161),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_338),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_374),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_117),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_96),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_54),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_249),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_306),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_316),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_18),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_184),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_235),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_198),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_136),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_373),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_44),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_202),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_361),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_256),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_45),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_23),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_168),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_37),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_218),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_14),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_185),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_101),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_71),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_83),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_152),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_115),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_342),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_65),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_21),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_94),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_332),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_30),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_323),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_309),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_265),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_27),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_220),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_87),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_22),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_305),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_122),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_288),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_346),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_24),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_171),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_280),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_240),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_56),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_227),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_226),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_304),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_145),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_223),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_369),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_266),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_358),
.Y(n_547)
);

CKINVDCx14_ASAP7_75t_R g548 ( 
.A(n_192),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_84),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_143),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_167),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_351),
.Y(n_552)
);

INVx1_ASAP7_75t_SL g553 ( 
.A(n_324),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_2),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_172),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_137),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_200),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_38),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_311),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_334),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_181),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_127),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_377),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_355),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_368),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_290),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_120),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_384),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_88),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_314),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_272),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_98),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_378),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_85),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_163),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_291),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_236),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_345),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_42),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_138),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_282),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_65),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_75),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_86),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_319),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_11),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_352),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_370),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_423),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_562),
.B(n_0),
.Y(n_590)
);

INVx5_ASAP7_75t_L g591 ( 
.A(n_501),
.Y(n_591)
);

BUFx8_ASAP7_75t_SL g592 ( 
.A(n_584),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_562),
.B(n_0),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_562),
.B(n_1),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_530),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_511),
.B(n_2),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_389),
.Y(n_597)
);

BUFx12f_ASAP7_75t_L g598 ( 
.A(n_422),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_410),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_501),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_423),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_423),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_391),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_388),
.B(n_3),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_392),
.B(n_401),
.Y(n_605)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_501),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_530),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_501),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_410),
.Y(n_609)
);

BUFx12f_ASAP7_75t_L g610 ( 
.A(n_422),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_409),
.B(n_553),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_548),
.B(n_3),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_524),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_453),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_388),
.B(n_4),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_524),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_393),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_524),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_523),
.B(n_4),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_539),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_524),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_573),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_453),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_573),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_417),
.B(n_5),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_458),
.B(n_6),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_573),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_390),
.B(n_6),
.Y(n_628)
);

INVx5_ASAP7_75t_L g629 ( 
.A(n_573),
.Y(n_629)
);

BUFx12f_ASAP7_75t_L g630 ( 
.A(n_422),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_458),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_491),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_491),
.B(n_7),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_544),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_544),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_492),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_547),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_417),
.B(n_7),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_427),
.B(n_475),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_539),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_547),
.B(n_8),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_427),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_475),
.B(n_8),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_479),
.B(n_9),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_479),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_548),
.B(n_10),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_492),
.B(n_10),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_418),
.Y(n_648)
);

BUFx8_ASAP7_75t_SL g649 ( 
.A(n_584),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_528),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_434),
.Y(n_651)
);

INVx5_ASAP7_75t_L g652 ( 
.A(n_528),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_528),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_396),
.B(n_12),
.Y(n_654)
);

INVx5_ASAP7_75t_L g655 ( 
.A(n_440),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_440),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_481),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_505),
.B(n_12),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_505),
.B(n_13),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_486),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_506),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_508),
.Y(n_662)
);

NOR2x1_ASAP7_75t_L g663 ( 
.A(n_508),
.B(n_395),
.Y(n_663)
);

BUFx8_ASAP7_75t_SL g664 ( 
.A(n_586),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_516),
.B(n_14),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_462),
.B(n_15),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_482),
.B(n_15),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_423),
.Y(n_668)
);

BUFx12f_ASAP7_75t_L g669 ( 
.A(n_400),
.Y(n_669)
);

NOR2x1_ASAP7_75t_L g670 ( 
.A(n_397),
.B(n_90),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_406),
.Y(n_671)
);

BUFx8_ASAP7_75t_L g672 ( 
.A(n_507),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_557),
.B(n_16),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_529),
.B(n_16),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_549),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_423),
.Y(n_676)
);

BUFx12f_ASAP7_75t_L g677 ( 
.A(n_415),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_554),
.B(n_402),
.Y(n_678)
);

BUFx12f_ASAP7_75t_L g679 ( 
.A(n_416),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_403),
.B(n_17),
.Y(n_680)
);

INVx5_ASAP7_75t_L g681 ( 
.A(n_423),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_405),
.Y(n_682)
);

BUFx8_ASAP7_75t_L g683 ( 
.A(n_423),
.Y(n_683)
);

BUFx8_ASAP7_75t_SL g684 ( 
.A(n_586),
.Y(n_684)
);

INVx5_ASAP7_75t_L g685 ( 
.A(n_394),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_408),
.B(n_17),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_464),
.B(n_527),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_431),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_398),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_411),
.Y(n_690)
);

BUFx12f_ASAP7_75t_L g691 ( 
.A(n_432),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_413),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_611),
.A2(n_665),
.B1(n_654),
.B2(n_646),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_636),
.B(n_433),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_600),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_R g696 ( 
.A1(n_619),
.A2(n_514),
.B1(n_569),
.B2(n_519),
.Y(n_696)
);

AO22x2_ASAP7_75t_L g697 ( 
.A1(n_596),
.A2(n_425),
.B1(n_442),
.B2(n_428),
.Y(n_697)
);

OAI22xp33_ASAP7_75t_L g698 ( 
.A1(n_596),
.A2(n_447),
.B1(n_448),
.B2(n_445),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_611),
.A2(n_612),
.B1(n_687),
.B2(n_605),
.Y(n_699)
);

OAI22xp33_ASAP7_75t_L g700 ( 
.A1(n_653),
.A2(n_474),
.B1(n_476),
.B2(n_451),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_669),
.A2(n_545),
.B1(n_456),
.B2(n_424),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_653),
.B(n_399),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_655),
.B(n_404),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_R g704 ( 
.A1(n_628),
.A2(n_419),
.B1(n_446),
.B2(n_443),
.Y(n_704)
);

AO22x2_ASAP7_75t_L g705 ( 
.A1(n_626),
.A2(n_450),
.B1(n_457),
.B2(n_449),
.Y(n_705)
);

OAI22xp33_ASAP7_75t_L g706 ( 
.A1(n_673),
.A2(n_496),
.B1(n_502),
.B2(n_478),
.Y(n_706)
);

AO22x2_ASAP7_75t_L g707 ( 
.A1(n_626),
.A2(n_465),
.B1(n_467),
.B2(n_460),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_677),
.A2(n_456),
.B1(n_545),
.B2(n_525),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_650),
.Y(n_709)
);

OAI22xp33_ASAP7_75t_L g710 ( 
.A1(n_673),
.A2(n_509),
.B1(n_520),
.B2(n_515),
.Y(n_710)
);

XNOR2xp5_ASAP7_75t_L g711 ( 
.A(n_656),
.B(n_414),
.Y(n_711)
);

OA22x2_ASAP7_75t_L g712 ( 
.A1(n_614),
.A2(n_558),
.B1(n_574),
.B2(n_535),
.Y(n_712)
);

OAI22xp33_ASAP7_75t_L g713 ( 
.A1(n_590),
.A2(n_582),
.B1(n_583),
.B2(n_579),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_679),
.A2(n_570),
.B1(n_575),
.B2(n_555),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_691),
.A2(n_412),
.B1(n_420),
.B2(n_407),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_597),
.B(n_484),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_655),
.B(n_421),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_600),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_603),
.B(n_490),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_655),
.B(n_426),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_617),
.B(n_493),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_666),
.A2(n_430),
.B1(n_435),
.B2(n_429),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_652),
.B(n_497),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_688),
.A2(n_437),
.B1(n_438),
.B2(n_436),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_655),
.B(n_439),
.Y(n_725)
);

OAI22xp33_ASAP7_75t_L g726 ( 
.A1(n_590),
.A2(n_521),
.B1(n_533),
.B2(n_500),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_688),
.A2(n_444),
.B1(n_452),
.B2(n_441),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_671),
.B(n_454),
.Y(n_728)
);

AO22x2_ASAP7_75t_L g729 ( 
.A1(n_633),
.A2(n_540),
.B1(n_546),
.B2(n_534),
.Y(n_729)
);

OAI22xp33_ASAP7_75t_L g730 ( 
.A1(n_594),
.A2(n_551),
.B1(n_559),
.B2(n_550),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_R g731 ( 
.A1(n_592),
.A2(n_566),
.B1(n_567),
.B2(n_560),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_642),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_L g733 ( 
.A1(n_594),
.A2(n_585),
.B1(n_588),
.B2(n_581),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_598),
.A2(n_610),
.B1(n_630),
.B2(n_593),
.Y(n_734)
);

AO22x2_ASAP7_75t_L g735 ( 
.A1(n_633),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_593),
.A2(n_459),
.B1(n_461),
.B2(n_455),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_689),
.B(n_463),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_599),
.B(n_609),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_641),
.A2(n_468),
.B1(n_469),
.B2(n_466),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_652),
.B(n_470),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_652),
.B(n_632),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_652),
.B(n_471),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_600),
.Y(n_743)
);

AO22x2_ASAP7_75t_L g744 ( 
.A1(n_641),
.A2(n_23),
.B1(n_19),
.B2(n_21),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_608),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_667),
.B(n_472),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_632),
.B(n_473),
.Y(n_747)
);

OAI22xp33_ASAP7_75t_L g748 ( 
.A1(n_667),
.A2(n_480),
.B1(n_483),
.B2(n_477),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_685),
.B(n_485),
.Y(n_749)
);

AO22x2_ASAP7_75t_L g750 ( 
.A1(n_680),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_680),
.A2(n_488),
.B1(n_489),
.B2(n_487),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_685),
.B(n_587),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_686),
.A2(n_495),
.B1(n_498),
.B2(n_494),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_686),
.A2(n_503),
.B1(n_504),
.B2(n_499),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_604),
.A2(n_512),
.B1(n_513),
.B2(n_510),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_623),
.B(n_517),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_642),
.Y(n_757)
);

CKINVDCx6p67_ASAP7_75t_R g758 ( 
.A(n_631),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_674),
.B(n_25),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_608),
.Y(n_760)
);

AO22x2_ASAP7_75t_L g761 ( 
.A1(n_647),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_642),
.Y(n_762)
);

OAI22xp33_ASAP7_75t_L g763 ( 
.A1(n_604),
.A2(n_522),
.B1(n_526),
.B2(n_518),
.Y(n_763)
);

OAI22xp33_ASAP7_75t_SL g764 ( 
.A1(n_615),
.A2(n_532),
.B1(n_536),
.B2(n_531),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_631),
.B(n_537),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_625),
.A2(n_541),
.B1(n_542),
.B2(n_538),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_631),
.B(n_28),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_634),
.B(n_543),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_674),
.B(n_29),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_645),
.Y(n_770)
);

AO22x2_ASAP7_75t_L g771 ( 
.A1(n_615),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_L g772 ( 
.A1(n_644),
.A2(n_556),
.B1(n_561),
.B2(n_552),
.Y(n_772)
);

OAI22xp33_ASAP7_75t_SL g773 ( 
.A1(n_644),
.A2(n_564),
.B1(n_565),
.B2(n_563),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_685),
.B(n_568),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_634),
.B(n_571),
.Y(n_775)
);

OA22x2_ASAP7_75t_L g776 ( 
.A1(n_648),
.A2(n_576),
.B1(n_577),
.B2(n_572),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_625),
.A2(n_580),
.B1(n_578),
.B2(n_34),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_634),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_635),
.B(n_91),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_695),
.Y(n_780)
);

OR2x6_ASAP7_75t_L g781 ( 
.A(n_761),
.B(n_648),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_738),
.Y(n_782)
);

CKINVDCx20_ASAP7_75t_R g783 ( 
.A(n_711),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_778),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_732),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_757),
.Y(n_786)
);

BUFx6f_ASAP7_75t_SL g787 ( 
.A(n_709),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_762),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_770),
.Y(n_789)
);

OR2x6_ASAP7_75t_L g790 ( 
.A(n_761),
.B(n_651),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_718),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_746),
.B(n_589),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_743),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_714),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_745),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_760),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_767),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_765),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_768),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_775),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_779),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_SL g802 ( 
.A(n_698),
.B(n_638),
.Y(n_802)
);

INVx4_ASAP7_75t_SL g803 ( 
.A(n_741),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_694),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_756),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_758),
.Y(n_806)
);

AND2x6_ASAP7_75t_L g807 ( 
.A(n_693),
.B(n_670),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_699),
.B(n_635),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_702),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_747),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_723),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_721),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_712),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_705),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_759),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_705),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_707),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_701),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_766),
.B(n_635),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_708),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_715),
.Y(n_821)
);

XOR2x2_ASAP7_75t_L g822 ( 
.A(n_696),
.B(n_592),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_707),
.Y(n_823)
);

INVxp67_ASAP7_75t_SL g824 ( 
.A(n_726),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_729),
.Y(n_825)
);

INVxp33_ASAP7_75t_L g826 ( 
.A(n_716),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_728),
.B(n_637),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_749),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_729),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_697),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_697),
.Y(n_831)
);

NAND2x1p5_ASAP7_75t_L g832 ( 
.A(n_703),
.B(n_663),
.Y(n_832)
);

INVxp33_ASAP7_75t_L g833 ( 
.A(n_719),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_776),
.Y(n_834)
);

INVxp33_ASAP7_75t_SL g835 ( 
.A(n_734),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_735),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_737),
.B(n_740),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_717),
.Y(n_838)
);

XNOR2xp5_ASAP7_75t_L g839 ( 
.A(n_764),
.B(n_773),
.Y(n_839)
);

XNOR2xp5_ASAP7_75t_SL g840 ( 
.A(n_704),
.B(n_649),
.Y(n_840)
);

INVxp33_ASAP7_75t_L g841 ( 
.A(n_724),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_727),
.B(n_637),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_720),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_730),
.B(n_601),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_722),
.B(n_685),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_739),
.B(n_637),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_725),
.B(n_742),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_736),
.B(n_595),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_774),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_755),
.A2(n_659),
.B(n_643),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_752),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_751),
.B(n_595),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_759),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_769),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_735),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_769),
.Y(n_856)
);

INVx4_ASAP7_75t_SL g857 ( 
.A(n_744),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_744),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_733),
.B(n_602),
.Y(n_859)
);

CKINVDCx20_ASAP7_75t_R g860 ( 
.A(n_753),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_754),
.B(n_700),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_777),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_748),
.B(n_659),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_763),
.B(n_690),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_731),
.B(n_591),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_750),
.Y(n_866)
);

INVxp33_ASAP7_75t_L g867 ( 
.A(n_750),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_771),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_771),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_772),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_713),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_706),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_710),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_828),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_812),
.B(n_645),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_782),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_826),
.B(n_651),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_792),
.B(n_645),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_780),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_791),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_798),
.B(n_661),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_828),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_830),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_792),
.B(n_662),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_837),
.B(n_662),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_785),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_828),
.Y(n_887)
);

INVx2_ASAP7_75t_SL g888 ( 
.A(n_827),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_793),
.Y(n_889)
);

OAI21x1_ASAP7_75t_L g890 ( 
.A1(n_801),
.A2(n_639),
.B(n_668),
.Y(n_890)
);

NOR2xp67_ASAP7_75t_L g891 ( 
.A(n_806),
.B(n_639),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_795),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_849),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_847),
.B(n_662),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_799),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_796),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_863),
.B(n_682),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_786),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_833),
.B(n_607),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_788),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_789),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_808),
.B(n_607),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_831),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_784),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_800),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_873),
.B(n_620),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_809),
.B(n_682),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_838),
.B(n_692),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_843),
.Y(n_909)
);

AND2x2_ASAP7_75t_SL g910 ( 
.A(n_802),
.B(n_638),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_797),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_851),
.B(n_682),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_811),
.B(n_682),
.Y(n_913)
);

INVx4_ASAP7_75t_L g914 ( 
.A(n_803),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_850),
.A2(n_658),
.B(n_643),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_848),
.B(n_620),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_807),
.B(n_683),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_807),
.B(n_683),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_807),
.B(n_658),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_804),
.B(n_640),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_805),
.Y(n_921)
);

INVxp33_ASAP7_75t_L g922 ( 
.A(n_864),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_807),
.B(n_676),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_819),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_802),
.B(n_591),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_857),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_810),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_844),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_813),
.B(n_657),
.Y(n_929)
);

AND2x2_ASAP7_75t_SL g930 ( 
.A(n_861),
.B(n_678),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_870),
.B(n_591),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_850),
.B(n_591),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_841),
.B(n_678),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_834),
.B(n_657),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_844),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_832),
.Y(n_936)
);

NOR2xp67_ASAP7_75t_R g937 ( 
.A(n_814),
.B(n_660),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_783),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_872),
.B(n_871),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_832),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_859),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_859),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_824),
.B(n_846),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_853),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_824),
.B(n_606),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_816),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_803),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_803),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_852),
.B(n_640),
.Y(n_949)
);

AND2x2_ASAP7_75t_SL g950 ( 
.A(n_845),
.B(n_613),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_817),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_842),
.B(n_606),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_815),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_823),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_854),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_862),
.B(n_606),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_825),
.B(n_606),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_857),
.B(n_829),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_815),
.B(n_660),
.Y(n_959)
);

INVxp67_ASAP7_75t_L g960 ( 
.A(n_856),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_781),
.B(n_675),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_869),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_868),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_857),
.Y(n_964)
);

AND2x6_ASAP7_75t_L g965 ( 
.A(n_858),
.B(n_613),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_866),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_821),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_781),
.B(n_675),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_836),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_781),
.B(n_608),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_787),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_839),
.B(n_616),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_790),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_790),
.Y(n_974)
);

OR2x6_ASAP7_75t_L g975 ( 
.A(n_940),
.B(n_790),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_882),
.Y(n_976)
);

INVx4_ASAP7_75t_L g977 ( 
.A(n_882),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_941),
.B(n_836),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_886),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_874),
.B(n_865),
.Y(n_980)
);

INVxp67_ASAP7_75t_SL g981 ( 
.A(n_882),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_963),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_922),
.B(n_867),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_942),
.Y(n_984)
);

NAND2x1p5_ASAP7_75t_L g985 ( 
.A(n_874),
.B(n_855),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_941),
.B(n_855),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_933),
.B(n_860),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_899),
.Y(n_988)
);

NAND2x1p5_ASAP7_75t_L g989 ( 
.A(n_882),
.B(n_622),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_930),
.B(n_835),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_886),
.Y(n_991)
);

AND2x2_ASAP7_75t_SL g992 ( 
.A(n_910),
.B(n_840),
.Y(n_992)
);

NAND2x1p5_ASAP7_75t_L g993 ( 
.A(n_887),
.B(n_622),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_901),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_930),
.B(n_622),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_901),
.Y(n_996)
);

CKINVDCx6p67_ASAP7_75t_R g997 ( 
.A(n_967),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_938),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_963),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_933),
.B(n_794),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_898),
.Y(n_1001)
);

BUFx12f_ASAP7_75t_L g1002 ( 
.A(n_971),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_943),
.B(n_822),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_928),
.B(n_624),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_900),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_888),
.B(n_887),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_920),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_877),
.B(n_818),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_938),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_887),
.B(n_820),
.Y(n_1010)
);

OR2x6_ASAP7_75t_L g1011 ( 
.A(n_940),
.B(n_649),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_887),
.B(n_92),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_SL g1013 ( 
.A(n_910),
.B(n_787),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_942),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_942),
.B(n_613),
.Y(n_1015)
);

NAND2x1p5_ASAP7_75t_L g1016 ( 
.A(n_940),
.B(n_624),
.Y(n_1016)
);

OR2x6_ASAP7_75t_L g1017 ( 
.A(n_940),
.B(n_664),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_967),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_916),
.B(n_949),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_893),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_942),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_902),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_922),
.B(n_664),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_951),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_924),
.B(n_684),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_959),
.B(n_684),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_935),
.B(n_624),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_897),
.B(n_613),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_944),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_895),
.B(n_93),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_906),
.B(n_32),
.Y(n_1031)
);

AND2x6_ASAP7_75t_L g1032 ( 
.A(n_947),
.B(n_618),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_895),
.B(n_95),
.Y(n_1033)
);

INVx5_ASAP7_75t_L g1034 ( 
.A(n_914),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_951),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_893),
.B(n_97),
.Y(n_1036)
);

INVx6_ASAP7_75t_SL g1037 ( 
.A(n_934),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_971),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_893),
.B(n_102),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_893),
.Y(n_1040)
);

NOR2x1_ASAP7_75t_R g1041 ( 
.A(n_936),
.B(n_681),
.Y(n_1041)
);

OR2x6_ASAP7_75t_SL g1042 ( 
.A(n_917),
.B(n_672),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_974),
.B(n_103),
.Y(n_1043)
);

INVx4_ASAP7_75t_L g1044 ( 
.A(n_914),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_974),
.B(n_104),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_911),
.B(n_33),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_894),
.B(n_618),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_963),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_891),
.B(n_33),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_969),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_SL g1051 ( 
.A(n_998),
.Y(n_1051)
);

BUFx12f_ASAP7_75t_L g1052 ( 
.A(n_1009),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1024),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_SL g1054 ( 
.A(n_1011),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_1038),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_1007),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_1018),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_982),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_1020),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_1029),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1024),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_1020),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_1020),
.Y(n_1063)
);

INVx5_ASAP7_75t_L g1064 ( 
.A(n_976),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1035),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_976),
.Y(n_1066)
);

INVxp67_ASAP7_75t_SL g1067 ( 
.A(n_976),
.Y(n_1067)
);

INVx5_ASAP7_75t_L g1068 ( 
.A(n_1040),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_999),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_1048),
.Y(n_1070)
);

INVx5_ASAP7_75t_L g1071 ( 
.A(n_1040),
.Y(n_1071)
);

BUFx2_ASAP7_75t_SL g1072 ( 
.A(n_1048),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_1010),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_1007),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1035),
.Y(n_1075)
);

INVx5_ASAP7_75t_L g1076 ( 
.A(n_1040),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_1010),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_1048),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_1034),
.Y(n_1079)
);

INVx8_ASAP7_75t_L g1080 ( 
.A(n_1034),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_997),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_979),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_991),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_994),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_996),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_988),
.B(n_909),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_1034),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_985),
.Y(n_1088)
);

OR2x6_ASAP7_75t_L g1089 ( 
.A(n_975),
.B(n_936),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_984),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1001),
.Y(n_1091)
);

BUFx8_ASAP7_75t_L g1092 ( 
.A(n_1002),
.Y(n_1092)
);

BUFx12f_ASAP7_75t_SL g1093 ( 
.A(n_1011),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1019),
.B(n_885),
.Y(n_1094)
);

NAND2x1p5_ASAP7_75t_L g1095 ( 
.A(n_1044),
.B(n_947),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1005),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_977),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_977),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_1030),
.B(n_958),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_984),
.B(n_909),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_1044),
.Y(n_1101)
);

INVx4_ASAP7_75t_L g1102 ( 
.A(n_1006),
.Y(n_1102)
);

BUFx2_ASAP7_75t_SL g1103 ( 
.A(n_980),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1014),
.Y(n_1104)
);

INVxp67_ASAP7_75t_SL g1105 ( 
.A(n_981),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1014),
.Y(n_1106)
);

BUFx8_ASAP7_75t_L g1107 ( 
.A(n_1026),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_1008),
.Y(n_1108)
);

NAND2x1p5_ASAP7_75t_L g1109 ( 
.A(n_1036),
.B(n_948),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1021),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_1017),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_1050),
.Y(n_1112)
);

BUFx12f_ASAP7_75t_L g1113 ( 
.A(n_1092),
.Y(n_1113)
);

INVx6_ASAP7_75t_L g1114 ( 
.A(n_1080),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1061),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1053),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_SL g1117 ( 
.A1(n_1079),
.A2(n_1039),
.B(n_1036),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1075),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_1055),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1061),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_SL g1121 ( 
.A1(n_1054),
.A2(n_987),
.B1(n_1000),
.B2(n_1013),
.Y(n_1121)
);

INVx8_ASAP7_75t_L g1122 ( 
.A(n_1080),
.Y(n_1122)
);

CKINVDCx11_ASAP7_75t_R g1123 ( 
.A(n_1052),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1094),
.A2(n_915),
.B1(n_1049),
.B2(n_919),
.Y(n_1124)
);

NAND2x1p5_ASAP7_75t_L g1125 ( 
.A(n_1068),
.B(n_1012),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_1079),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1065),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1086),
.A2(n_939),
.B1(n_950),
.B2(n_990),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_1056),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1086),
.A2(n_950),
.B1(n_1031),
.B2(n_992),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1109),
.A2(n_1022),
.B1(n_1021),
.B2(n_986),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1108),
.B(n_1022),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1065),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_1057),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1073),
.A2(n_1023),
.B1(n_1013),
.B2(n_988),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1082),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_1091),
.A2(n_925),
.B1(n_1003),
.B2(n_1046),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_1057),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1082),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1099),
.B(n_978),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1079),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_SL g1142 ( 
.A1(n_1054),
.A2(n_1030),
.B1(n_1033),
.B2(n_1039),
.Y(n_1142)
);

OAI22x1_ASAP7_75t_L g1143 ( 
.A1(n_1077),
.A2(n_1033),
.B1(n_1045),
.B2(n_1043),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1096),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_1081),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_1109),
.A2(n_1105),
.B1(n_1099),
.B2(n_986),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1090),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_1056),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1090),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_SL g1150 ( 
.A1(n_1052),
.A2(n_1012),
.B1(n_1025),
.B2(n_1017),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1083),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1084),
.A2(n_925),
.B1(n_905),
.B2(n_921),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1099),
.B(n_978),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1085),
.A2(n_927),
.B1(n_995),
.B2(n_876),
.Y(n_1154)
);

CKINVDCx11_ASAP7_75t_R g1155 ( 
.A(n_1081),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1104),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1106),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1105),
.A2(n_983),
.B1(n_1006),
.B2(n_972),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1110),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_SL g1160 ( 
.A1(n_1111),
.A2(n_1045),
.B1(n_1043),
.B2(n_918),
.Y(n_1160)
);

INVx4_ASAP7_75t_L g1161 ( 
.A(n_1080),
.Y(n_1161)
);

INVxp67_ASAP7_75t_SL g1162 ( 
.A(n_1067),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1100),
.A2(n_908),
.B1(n_881),
.B2(n_932),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_1058),
.Y(n_1164)
);

BUFx2_ASAP7_75t_SL g1165 ( 
.A(n_1051),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1100),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_1058),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_1055),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1112),
.Y(n_1169)
);

BUFx8_ASAP7_75t_L g1170 ( 
.A(n_1051),
.Y(n_1170)
);

CKINVDCx20_ASAP7_75t_R g1171 ( 
.A(n_1092),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1116),
.Y(n_1172)
);

BUFx12f_ASAP7_75t_L g1173 ( 
.A(n_1123),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1121),
.A2(n_908),
.B1(n_881),
.B2(n_923),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1164),
.Y(n_1175)
);

AOI222xp33_ASAP7_75t_L g1176 ( 
.A1(n_1130),
.A2(n_881),
.B1(n_672),
.B2(n_1074),
.C1(n_908),
.C2(n_960),
.Y(n_1176)
);

INVxp67_ASAP7_75t_L g1177 ( 
.A(n_1129),
.Y(n_1177)
);

BUFx12f_ASAP7_75t_L g1178 ( 
.A(n_1123),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1118),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1121),
.A2(n_1093),
.B1(n_962),
.B2(n_1107),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1130),
.A2(n_1093),
.B1(n_1107),
.B2(n_875),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1165),
.A2(n_1111),
.B1(n_1088),
.B2(n_1092),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1128),
.A2(n_955),
.B1(n_907),
.B2(n_889),
.Y(n_1183)
);

BUFx12f_ASAP7_75t_L g1184 ( 
.A(n_1113),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_SL g1185 ( 
.A1(n_1158),
.A2(n_1088),
.B1(n_1103),
.B2(n_1060),
.Y(n_1185)
);

OAI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1135),
.A2(n_1089),
.B1(n_975),
.B2(n_1102),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_SL g1187 ( 
.A1(n_1150),
.A2(n_980),
.B(n_968),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1157),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1160),
.A2(n_1069),
.B1(n_970),
.B2(n_892),
.Y(n_1189)
);

OAI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1140),
.A2(n_1089),
.B1(n_1102),
.B2(n_963),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1132),
.B(n_1069),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_SL g1192 ( 
.A1(n_1150),
.A2(n_961),
.B(n_973),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1160),
.A2(n_1137),
.B1(n_1128),
.B2(n_1142),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1137),
.A2(n_880),
.B1(n_1089),
.B2(n_896),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1153),
.B(n_883),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1159),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1144),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1168),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1115),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1142),
.A2(n_896),
.B1(n_904),
.B2(n_879),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1138),
.B(n_973),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1162),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_SL g1203 ( 
.A1(n_1124),
.A2(n_960),
.B(n_934),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1170),
.A2(n_953),
.B1(n_1087),
.B2(n_1079),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_SL g1205 ( 
.A1(n_1170),
.A2(n_1087),
.B1(n_1072),
.B2(n_1067),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1143),
.A2(n_931),
.B1(n_912),
.B2(n_956),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_SL g1207 ( 
.A1(n_1134),
.A2(n_1167),
.B1(n_1171),
.B2(n_1146),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1147),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1145),
.Y(n_1209)
);

NAND3xp33_ASAP7_75t_L g1210 ( 
.A(n_1124),
.B(n_952),
.C(n_913),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1151),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1152),
.A2(n_903),
.B1(n_883),
.B2(n_884),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1148),
.B(n_903),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_SL g1214 ( 
.A1(n_1119),
.A2(n_1087),
.B1(n_1068),
.B2(n_1076),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1149),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1156),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1152),
.A2(n_878),
.B1(n_1027),
.B2(n_1004),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1154),
.A2(n_934),
.B1(n_929),
.B2(n_945),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1139),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1141),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1154),
.A2(n_929),
.B1(n_954),
.B2(n_946),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1136),
.Y(n_1222)
);

AOI222xp33_ASAP7_75t_L g1223 ( 
.A1(n_1131),
.A2(n_929),
.B1(n_937),
.B2(n_1041),
.C1(n_946),
.C2(n_954),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1169),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1117),
.A2(n_1071),
.B1(n_1076),
.B2(n_1068),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1163),
.A2(n_965),
.B1(n_1037),
.B2(n_1070),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1122),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1163),
.A2(n_965),
.B1(n_1037),
.B2(n_1070),
.Y(n_1228)
);

BUFx8_ASAP7_75t_SL g1229 ( 
.A(n_1141),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1120),
.A2(n_1047),
.B1(n_1015),
.B2(n_1028),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1162),
.A2(n_1125),
.B1(n_1114),
.B2(n_1166),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1127),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1133),
.A2(n_965),
.B1(n_1078),
.B2(n_1015),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1155),
.A2(n_965),
.B1(n_1078),
.B2(n_1062),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1126),
.B(n_966),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1126),
.Y(n_1236)
);

NOR2xp67_ASAP7_75t_L g1237 ( 
.A(n_1161),
.B(n_1064),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_SL g1238 ( 
.A1(n_1125),
.A2(n_1042),
.B(n_966),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1155),
.A2(n_1047),
.B1(n_1028),
.B2(n_890),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1114),
.A2(n_1161),
.B1(n_1071),
.B2(n_1076),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1114),
.A2(n_1071),
.B1(n_1076),
.B2(n_1068),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1176),
.A2(n_1231),
.B1(n_1192),
.B2(n_1173),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_SL g1243 ( 
.A1(n_1178),
.A2(n_1122),
.B1(n_1141),
.B2(n_1087),
.Y(n_1243)
);

AOI222xp33_ASAP7_75t_L g1244 ( 
.A1(n_1193),
.A2(n_1041),
.B1(n_681),
.B2(n_957),
.C1(n_37),
.C2(n_38),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1181),
.A2(n_1141),
.B1(n_1062),
.B2(n_1063),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1181),
.A2(n_1063),
.B1(n_1059),
.B2(n_1122),
.Y(n_1246)
);

OAI221xp5_ASAP7_75t_L g1247 ( 
.A1(n_1180),
.A2(n_1016),
.B1(n_1095),
.B2(n_1059),
.C(n_964),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1186),
.A2(n_1180),
.B1(n_1207),
.B2(n_1185),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1191),
.B(n_926),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1186),
.A2(n_965),
.B1(n_1097),
.B2(n_1101),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1189),
.A2(n_1097),
.B1(n_1101),
.B2(n_1098),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1194),
.A2(n_1095),
.B1(n_1071),
.B2(n_1098),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_SL g1253 ( 
.A1(n_1182),
.A2(n_1097),
.B1(n_1101),
.B2(n_1064),
.Y(n_1253)
);

NAND3xp33_ASAP7_75t_L g1254 ( 
.A(n_1203),
.B(n_1101),
.C(n_1097),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1177),
.B(n_1066),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1174),
.A2(n_1066),
.B1(n_890),
.B2(n_1032),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1183),
.A2(n_1066),
.B1(n_1032),
.B2(n_989),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_SL g1258 ( 
.A1(n_1175),
.A2(n_1064),
.B1(n_1066),
.B2(n_958),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1183),
.A2(n_1032),
.B1(n_993),
.B2(n_1064),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1225),
.A2(n_948),
.B(n_627),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_SL g1261 ( 
.A1(n_1202),
.A2(n_1195),
.B1(n_1240),
.B2(n_1241),
.Y(n_1261)
);

AOI222xp33_ASAP7_75t_L g1262 ( 
.A1(n_1187),
.A2(n_681),
.B1(n_35),
.B2(n_36),
.C1(n_39),
.C2(n_40),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1210),
.A2(n_1032),
.B(n_958),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1223),
.A2(n_681),
.B1(n_627),
.B2(n_618),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1200),
.A2(n_627),
.B1(n_618),
.B2(n_621),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1204),
.A2(n_629),
.B1(n_616),
.B2(n_621),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_SL g1267 ( 
.A1(n_1202),
.A2(n_621),
.B1(n_36),
.B2(n_34),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1212),
.A2(n_629),
.B1(n_616),
.B2(n_621),
.Y(n_1268)
);

AOI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1238),
.A2(n_629),
.B1(n_616),
.B2(n_40),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1206),
.A2(n_1190),
.B1(n_1201),
.B2(n_1218),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1190),
.A2(n_629),
.B1(n_42),
.B2(n_35),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1198),
.B(n_106),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1218),
.A2(n_44),
.B1(n_39),
.B2(n_43),
.Y(n_1273)
);

NAND2xp33_ASAP7_75t_SL g1274 ( 
.A(n_1227),
.B(n_43),
.Y(n_1274)
);

NOR3xp33_ASAP7_75t_L g1275 ( 
.A(n_1205),
.B(n_45),
.C(n_46),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1212),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1184),
.A2(n_1226),
.B1(n_1228),
.B2(n_1216),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1224),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1219),
.B(n_107),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1209),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1197),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1211),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1172),
.B(n_56),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1199),
.B(n_57),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1234),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1232),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1214),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1179),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1188),
.A2(n_1196),
.B1(n_1221),
.B2(n_1232),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1221),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1213),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1217),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_1292)
);

OAI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1222),
.A2(n_1208),
.B1(n_1215),
.B2(n_1236),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1230),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1233),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_1295)
);

AOI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1217),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1230),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1235),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1220),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1239),
.A2(n_1229),
.B1(n_1220),
.B2(n_1237),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1239),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1220),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1220),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1176),
.A2(n_82),
.B1(n_84),
.B2(n_86),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1255),
.B(n_88),
.Y(n_1305)
);

OAI221xp5_ASAP7_75t_SL g1306 ( 
.A1(n_1304),
.A2(n_1291),
.B1(n_1262),
.B2(n_1242),
.C(n_1280),
.Y(n_1306)
);

OAI221xp5_ASAP7_75t_SL g1307 ( 
.A1(n_1269),
.A2(n_89),
.B1(n_109),
.B2(n_111),
.C(n_113),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1286),
.B(n_1289),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_SL g1309 ( 
.A1(n_1254),
.A2(n_1268),
.B(n_1297),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1249),
.B(n_1270),
.Y(n_1310)
);

NAND3xp33_ASAP7_75t_L g1311 ( 
.A(n_1275),
.B(n_89),
.C(n_114),
.Y(n_1311)
);

NAND3xp33_ASAP7_75t_L g1312 ( 
.A(n_1273),
.B(n_116),
.C(n_118),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1292),
.A2(n_119),
.B1(n_121),
.B2(n_123),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1248),
.B(n_125),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1273),
.B(n_126),
.C(n_129),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1296),
.B(n_130),
.C(n_135),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1303),
.B(n_139),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1261),
.B(n_140),
.Y(n_1318)
);

AOI221xp5_ASAP7_75t_L g1319 ( 
.A1(n_1276),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.C(n_147),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1293),
.B(n_148),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1244),
.A2(n_150),
.B(n_151),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1300),
.B(n_387),
.Y(n_1322)
);

NOR3xp33_ASAP7_75t_SL g1323 ( 
.A(n_1274),
.B(n_154),
.C(n_156),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_1284),
.Y(n_1324)
);

OAI221xp5_ASAP7_75t_L g1325 ( 
.A1(n_1294),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.C(n_162),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1277),
.B(n_164),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1293),
.B(n_165),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1283),
.B(n_166),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1247),
.B(n_1253),
.Y(n_1329)
);

NOR3xp33_ASAP7_75t_L g1330 ( 
.A(n_1302),
.B(n_170),
.C(n_173),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1294),
.B(n_174),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1279),
.B(n_175),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1301),
.A2(n_176),
.B1(n_177),
.B2(n_180),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1281),
.B(n_1282),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1288),
.B(n_183),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1278),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1299),
.B(n_190),
.Y(n_1337)
);

NAND3xp33_ASAP7_75t_L g1338 ( 
.A(n_1267),
.B(n_193),
.C(n_195),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1299),
.B(n_386),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1299),
.B(n_196),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_SL g1341 ( 
.A1(n_1287),
.A2(n_199),
.B(n_201),
.Y(n_1341)
);

OAI221xp5_ASAP7_75t_L g1342 ( 
.A1(n_1298),
.A2(n_203),
.B1(n_206),
.B2(n_207),
.C(n_208),
.Y(n_1342)
);

AOI221xp5_ASAP7_75t_L g1343 ( 
.A1(n_1285),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.C(n_213),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1299),
.B(n_214),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1251),
.B(n_215),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1245),
.B(n_216),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_SL g1347 ( 
.A1(n_1290),
.A2(n_217),
.B(n_219),
.Y(n_1347)
);

NOR3xp33_ASAP7_75t_L g1348 ( 
.A(n_1295),
.B(n_221),
.C(n_224),
.Y(n_1348)
);

NAND3xp33_ASAP7_75t_L g1349 ( 
.A(n_1271),
.B(n_228),
.C(n_232),
.Y(n_1349)
);

NAND3xp33_ASAP7_75t_L g1350 ( 
.A(n_1246),
.B(n_233),
.C(n_234),
.Y(n_1350)
);

NAND3xp33_ASAP7_75t_L g1351 ( 
.A(n_1250),
.B(n_237),
.C(n_238),
.Y(n_1351)
);

NAND3xp33_ASAP7_75t_L g1352 ( 
.A(n_1263),
.B(n_239),
.C(n_241),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1329),
.A2(n_1310),
.B1(n_1311),
.B2(n_1334),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1305),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1324),
.B(n_1272),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1308),
.B(n_1256),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1329),
.B(n_1257),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1320),
.B(n_1259),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1348),
.A2(n_1264),
.B1(n_1252),
.B2(n_1266),
.Y(n_1359)
);

NOR3xp33_ASAP7_75t_L g1360 ( 
.A(n_1306),
.B(n_1243),
.C(n_1258),
.Y(n_1360)
);

AND2x2_ASAP7_75t_SL g1361 ( 
.A(n_1318),
.B(n_1265),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1327),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1327),
.B(n_1260),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1337),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1344),
.Y(n_1365)
);

NAND3xp33_ASAP7_75t_L g1366 ( 
.A(n_1307),
.B(n_1316),
.C(n_1321),
.Y(n_1366)
);

AOI221xp5_ASAP7_75t_L g1367 ( 
.A1(n_1313),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.C(n_245),
.Y(n_1367)
);

NAND4xp25_ASAP7_75t_L g1368 ( 
.A(n_1312),
.B(n_246),
.C(n_247),
.D(n_248),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1328),
.B(n_250),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1326),
.B(n_1322),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1339),
.B(n_254),
.Y(n_1371)
);

OA211x2_ASAP7_75t_L g1372 ( 
.A1(n_1352),
.A2(n_255),
.B(n_257),
.C(n_258),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1340),
.B(n_261),
.Y(n_1373)
);

NAND3xp33_ASAP7_75t_SL g1374 ( 
.A(n_1341),
.B(n_262),
.C(n_263),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1317),
.B(n_267),
.Y(n_1375)
);

NOR3xp33_ASAP7_75t_L g1376 ( 
.A(n_1315),
.B(n_269),
.C(n_270),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1319),
.B(n_1323),
.C(n_1343),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1309),
.B(n_271),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1309),
.B(n_273),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1331),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1332),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1323),
.B(n_275),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1330),
.B(n_276),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1345),
.Y(n_1384)
);

AO21x2_ASAP7_75t_L g1385 ( 
.A1(n_1313),
.A2(n_278),
.B(n_281),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1364),
.Y(n_1386)
);

NOR3xp33_ASAP7_75t_L g1387 ( 
.A(n_1366),
.B(n_1325),
.C(n_1338),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1364),
.B(n_1314),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1354),
.B(n_1346),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1365),
.Y(n_1390)
);

NAND4xp75_ASAP7_75t_SL g1391 ( 
.A(n_1379),
.B(n_1347),
.C(n_1350),
.D(n_1351),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1365),
.B(n_1349),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1377),
.A2(n_1342),
.B1(n_1333),
.B2(n_1336),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1381),
.Y(n_1394)
);

NAND4xp75_ASAP7_75t_L g1395 ( 
.A(n_1379),
.B(n_1335),
.C(n_1336),
.D(n_289),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1380),
.B(n_283),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1354),
.B(n_285),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1381),
.Y(n_1398)
);

XOR2x2_ASAP7_75t_L g1399 ( 
.A(n_1355),
.B(n_292),
.Y(n_1399)
);

NAND4xp75_ASAP7_75t_L g1400 ( 
.A(n_1372),
.B(n_295),
.C(n_296),
.D(n_297),
.Y(n_1400)
);

NAND4xp75_ASAP7_75t_SL g1401 ( 
.A(n_1382),
.B(n_298),
.C(n_299),
.D(n_300),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1380),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1356),
.B(n_302),
.Y(n_1403)
);

NAND4xp75_ASAP7_75t_L g1404 ( 
.A(n_1367),
.B(n_1362),
.C(n_1382),
.D(n_1361),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1356),
.B(n_303),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1402),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1386),
.Y(n_1407)
);

XOR2x2_ASAP7_75t_L g1408 ( 
.A(n_1399),
.B(n_1370),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1402),
.Y(n_1409)
);

AO22x2_ASAP7_75t_L g1410 ( 
.A1(n_1404),
.A2(n_1391),
.B1(n_1390),
.B2(n_1394),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1398),
.B(n_1384),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1398),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1392),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1392),
.Y(n_1414)
);

OA22x2_ASAP7_75t_L g1415 ( 
.A1(n_1393),
.A2(n_1357),
.B1(n_1383),
.B2(n_1384),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1389),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1397),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1415),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1410),
.A2(n_1415),
.B1(n_1353),
.B2(n_1378),
.Y(n_1419)
);

OA22x2_ASAP7_75t_L g1420 ( 
.A1(n_1413),
.A2(n_1397),
.B1(n_1389),
.B2(n_1403),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1407),
.Y(n_1421)
);

OA22x2_ASAP7_75t_L g1422 ( 
.A1(n_1413),
.A2(n_1403),
.B1(n_1392),
.B2(n_1388),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1417),
.Y(n_1423)
);

AOI22x1_ASAP7_75t_L g1424 ( 
.A1(n_1410),
.A2(n_1378),
.B1(n_1363),
.B2(n_1399),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1414),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1410),
.A2(n_1387),
.B1(n_1360),
.B2(n_1395),
.Y(n_1426)
);

OAI22x1_ASAP7_75t_SL g1427 ( 
.A1(n_1414),
.A2(n_1401),
.B1(n_1385),
.B2(n_1374),
.Y(n_1427)
);

XOR2x2_ASAP7_75t_L g1428 ( 
.A(n_1408),
.B(n_1405),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1409),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1406),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1416),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1423),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1425),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1424),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1421),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1430),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1430),
.Y(n_1437)
);

OAI322xp33_ASAP7_75t_L g1438 ( 
.A1(n_1418),
.A2(n_1396),
.A3(n_1412),
.B1(n_1363),
.B2(n_1358),
.C1(n_1411),
.C2(n_1361),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1420),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1434),
.A2(n_1419),
.B1(n_1426),
.B2(n_1422),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_1432),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1434),
.A2(n_1419),
.B1(n_1426),
.B2(n_1427),
.Y(n_1442)
);

NAND4xp25_ASAP7_75t_SL g1443 ( 
.A(n_1433),
.B(n_1428),
.C(n_1357),
.D(n_1431),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1435),
.Y(n_1444)
);

AOI221xp5_ASAP7_75t_L g1445 ( 
.A1(n_1438),
.A2(n_1427),
.B1(n_1429),
.B2(n_1396),
.C(n_1411),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1444),
.Y(n_1446)
);

AOI22x1_ASAP7_75t_L g1447 ( 
.A1(n_1441),
.A2(n_1439),
.B1(n_1437),
.B2(n_1436),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1440),
.Y(n_1448)
);

AO22x2_ASAP7_75t_L g1449 ( 
.A1(n_1442),
.A2(n_1438),
.B1(n_1400),
.B2(n_1383),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1443),
.A2(n_1445),
.B1(n_1385),
.B2(n_1368),
.C(n_1376),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1446),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1447),
.Y(n_1452)
);

NOR4xp25_ASAP7_75t_L g1453 ( 
.A(n_1448),
.B(n_1369),
.C(n_1359),
.D(n_1358),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1449),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1449),
.A2(n_1450),
.B1(n_1375),
.B2(n_1373),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1446),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1452),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1454),
.B(n_1371),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1451),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1455),
.A2(n_308),
.B1(n_310),
.B2(n_315),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1456),
.Y(n_1461)
);

NAND4xp25_ASAP7_75t_L g1462 ( 
.A(n_1458),
.B(n_1453),
.C(n_325),
.D(n_326),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1457),
.A2(n_1453),
.B1(n_327),
.B2(n_328),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1459),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1461),
.Y(n_1465)
);

NOR2xp67_ASAP7_75t_L g1466 ( 
.A(n_1460),
.B(n_383),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1464),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1465),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1466),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1462),
.Y(n_1470)
);

INVx1_ASAP7_75t_SL g1471 ( 
.A(n_1463),
.Y(n_1471)
);

OAI22x1_ASAP7_75t_L g1472 ( 
.A1(n_1469),
.A2(n_330),
.B1(n_331),
.B2(n_333),
.Y(n_1472)
);

AO22x2_ASAP7_75t_L g1473 ( 
.A1(n_1467),
.A2(n_381),
.B1(n_336),
.B2(n_337),
.Y(n_1473)
);

OAI22x1_ASAP7_75t_L g1474 ( 
.A1(n_1471),
.A2(n_335),
.B1(n_339),
.B2(n_341),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1470),
.Y(n_1475)
);

NOR2x1_ASAP7_75t_L g1476 ( 
.A(n_1468),
.B(n_344),
.Y(n_1476)
);

INVxp67_ASAP7_75t_SL g1477 ( 
.A(n_1476),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1475),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1473),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1472),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1478),
.A2(n_1474),
.B1(n_348),
.B2(n_349),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1481),
.Y(n_1482)
);

OAI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1482),
.A2(n_1479),
.B1(n_1480),
.B2(n_1477),
.Y(n_1483)
);

OR2x2_ASAP7_75t_SL g1484 ( 
.A(n_1483),
.B(n_379),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1484),
.A2(n_353),
.B1(n_356),
.B2(n_359),
.Y(n_1485)
);

AOI211xp5_ASAP7_75t_L g1486 ( 
.A1(n_1485),
.A2(n_362),
.B(n_363),
.C(n_367),
.Y(n_1486)
);


endmodule