module fake_jpeg_5034_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_29),
.Y(n_47)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_41),
.Y(n_50)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_29),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_14),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_46),
.B(n_68),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_52),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_23),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_61),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_21),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_64),
.Y(n_94)
);

CKINVDCx11_ASAP7_75t_R g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_31),
.B(n_24),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_22),
.Y(n_70)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_30),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_32),
.B(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_40),
.A2(n_17),
.B1(n_27),
.B2(n_16),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_17),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_73),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_17),
.B(n_16),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_46),
.B(n_51),
.Y(n_99)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_30),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_95),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_26),
.B1(n_27),
.B2(n_16),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_96),
.B1(n_74),
.B2(n_62),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_30),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_110),
.B1(n_92),
.B2(n_87),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_84),
.B(n_71),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_62),
.B1(n_59),
.B2(n_65),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_113),
.B1(n_93),
.B2(n_78),
.Y(n_127)
);

CKINVDCx12_ASAP7_75t_R g101 ( 
.A(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_112),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_50),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_107),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_91),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_76),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_96),
.B1(n_85),
.B2(n_75),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_94),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_58),
.B1(n_60),
.B2(n_66),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_121),
.C(n_124),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_82),
.C(n_90),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_128),
.C(n_121),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_127),
.Y(n_131)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_97),
.C(n_105),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_60),
.B1(n_67),
.B2(n_49),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_133),
.Y(n_140)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_104),
.A3(n_107),
.B1(n_97),
.B2(n_99),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_132),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_98),
.C(n_103),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_118),
.Y(n_146)
);

AOI322xp5_ASAP7_75t_SL g137 ( 
.A1(n_120),
.A2(n_103),
.A3(n_11),
.B1(n_6),
.B2(n_8),
.C1(n_9),
.C2(n_49),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_137),
.B(n_139),
.Y(n_143)
);

A2O1A1O1Ixp25_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_67),
.B(n_2),
.C(n_4),
.D(n_1),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_142),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_147),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_128),
.C(n_116),
.Y(n_152)
);

AOI21x1_ASAP7_75t_L g148 ( 
.A1(n_146),
.A2(n_138),
.B(n_137),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_148),
.A2(n_140),
.B(n_144),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_143),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_126),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_140),
.B(n_135),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_151),
.B(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_153),
.B(n_130),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_156),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_152),
.C(n_149),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_159),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_124),
.B1(n_114),
.B2(n_111),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_117),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_162),
.Y(n_164)
);


endmodule