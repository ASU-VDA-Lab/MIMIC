module fake_jpeg_5079_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx8_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_14),
.B1(n_9),
.B2(n_16),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_10),
.B1(n_15),
.B2(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

AND2x4_ASAP7_75t_SL g32 ( 
.A(n_23),
.B(n_12),
.Y(n_32)
);

NOR2x1_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_14),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_3),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_20),
.A2(n_15),
.B1(n_10),
.B2(n_8),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_30),
.B1(n_24),
.B2(n_32),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_L g29 ( 
.A1(n_17),
.A2(n_12),
.B(n_8),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_40),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_37),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_27),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_44),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_47),
.B(n_48),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_42),
.B(n_34),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_27),
.C(n_28),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_49),
.B(n_26),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_28),
.B(n_4),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_54),
.A2(n_7),
.B(n_37),
.Y(n_55)
);


endmodule