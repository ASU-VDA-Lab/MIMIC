module fake_jpeg_30305_n_92 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_92);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_92;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

CKINVDCx6p67_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_1),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_35),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_53),
.C(n_28),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_33),
.B1(n_36),
.B2(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_33),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_36),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

AND2x6_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_57),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_63),
.B1(n_4),
.B2(n_5),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_62),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_2),
.Y(n_66)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_48),
.B1(n_46),
.B2(n_44),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_47),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_3),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_3),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_54),
.B(n_5),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_4),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_17),
.B1(n_27),
.B2(n_8),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_16),
.C(n_25),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_79),
.C(n_75),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_15),
.C(n_24),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_83),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_69),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_81),
.A2(n_72),
.B(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_77),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_76),
.B1(n_84),
.B2(n_6),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_76),
.B(n_7),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_89),
.A2(n_10),
.B(n_12),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_13),
.C(n_14),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_19),
.Y(n_92)
);


endmodule