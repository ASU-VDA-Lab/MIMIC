module fake_jpeg_5512_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_32),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_0),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_2),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_56),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_24),
.B1(n_18),
.B2(n_15),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_63),
.B1(n_5),
.B2(n_6),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_29),
.B1(n_24),
.B2(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_65),
.B1(n_66),
.B2(n_72),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_52),
.B(n_62),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_53),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_32),
.B(n_23),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_70),
.Y(n_79)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_60),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_31),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_21),
.B1(n_25),
.B2(n_23),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_35),
.A2(n_17),
.B1(n_15),
.B2(n_20),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_15),
.B1(n_28),
.B2(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_28),
.Y(n_68)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_14),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_20),
.B1(n_28),
.B2(n_5),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_3),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_75),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_4),
.Y(n_75)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_82),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_14),
.B(n_6),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_85),
.B(n_86),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_55),
.B1(n_44),
.B2(n_46),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_5),
.B(n_13),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_89),
.Y(n_100)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_10),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_70),
.Y(n_112)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_46),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_95),
.B(n_58),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_107),
.Y(n_119)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_70),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_75),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_56),
.B1(n_62),
.B2(n_69),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_104),
.B1(n_81),
.B2(n_90),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_112),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_77),
.A2(n_61),
.B1(n_67),
.B2(n_47),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_58),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_79),
.Y(n_126)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_109),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_111),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_85),
.B1(n_110),
.B2(n_112),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_111),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_121),
.B(n_124),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_113),
.C(n_105),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_103),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_113),
.C(n_96),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_96),
.B(n_105),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_93),
.B1(n_79),
.B2(n_78),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_127),
.A2(n_102),
.B1(n_97),
.B2(n_98),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_93),
.B1(n_87),
.B2(n_74),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_127),
.B(n_124),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_132),
.C(n_133),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_126),
.C(n_123),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_136),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_109),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_138),
.B(n_116),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_145),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_127),
.B1(n_122),
.B2(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_143),
.B(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_146),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_88),
.C(n_115),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_135),
.B(n_119),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_116),
.B1(n_99),
.B2(n_100),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_82),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_150),
.A2(n_141),
.B(n_147),
.C(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_145),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_140),
.A2(n_107),
.B(n_91),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_152),
.B(n_153),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_53),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_156),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_157),
.B(n_142),
.Y(n_160)
);

NAND2x1p5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_148),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_159),
.B(n_149),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_89),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_158),
.Y(n_164)
);


endmodule