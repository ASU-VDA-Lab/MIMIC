module fake_jpeg_10797_n_379 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_379);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_379;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_55),
.B(n_56),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_9),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_57),
.B(n_61),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_34),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_68),
.B(n_80),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_33),
.B(n_0),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_78),
.Y(n_123)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_71),
.Y(n_125)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_24),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_74),
.B(n_79),
.Y(n_147)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_41),
.A2(n_45),
.B1(n_37),
.B2(n_39),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_76),
.A2(n_42),
.B1(n_49),
.B2(n_51),
.Y(n_149)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_77),
.Y(n_166)
);

INVx2_ASAP7_75t_R g78 ( 
.A(n_33),
.Y(n_78)
);

INVx2_ASAP7_75t_R g79 ( 
.A(n_33),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_25),
.B(n_11),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_84),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_27),
.B(n_19),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_85),
.B(n_1),
.C(n_79),
.Y(n_164)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_25),
.B(n_11),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_87),
.B(n_90),
.Y(n_174)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_32),
.B(n_6),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_18),
.B(n_6),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_93),
.Y(n_148)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_92),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_32),
.B(n_6),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_23),
.Y(n_94)
);

CKINVDCx6p67_ASAP7_75t_R g127 ( 
.A(n_94),
.Y(n_127)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_34),
.B(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_96),
.B(n_98),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_19),
.B(n_14),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_99),
.A2(n_71),
.B(n_95),
.C(n_85),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_26),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_100),
.B(n_106),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_101),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_19),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_37),
.B(n_15),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_39),
.Y(n_112)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_26),
.Y(n_110)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_112),
.B(n_68),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_91),
.A2(n_45),
.B1(n_29),
.B2(n_30),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_119),
.A2(n_151),
.B1(n_155),
.B2(n_158),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_38),
.B(n_53),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_120),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_47),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_128),
.B(n_132),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_65),
.A2(n_23),
.B1(n_30),
.B2(n_29),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g193 ( 
.A1(n_131),
.A2(n_137),
.B(n_144),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_47),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_66),
.A2(n_23),
.B1(n_54),
.B2(n_35),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_69),
.A2(n_31),
.B(n_53),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_164),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_69),
.B(n_49),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_145),
.B(n_154),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_149),
.A2(n_156),
.B1(n_157),
.B2(n_175),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_72),
.A2(n_35),
.B1(n_54),
.B2(n_31),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_60),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_152),
.B(n_125),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_78),
.B(n_51),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_83),
.A2(n_43),
.B1(n_48),
.B2(n_42),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_84),
.A2(n_43),
.B1(n_48),
.B2(n_26),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_85),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_97),
.A2(n_1),
.B1(n_102),
.B2(n_105),
.Y(n_158)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_81),
.Y(n_168)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

OR2x2_ASAP7_75t_SL g189 ( 
.A(n_173),
.B(n_106),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_109),
.A2(n_59),
.B1(n_111),
.B2(n_62),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_146),
.A2(n_94),
.B1(n_82),
.B2(n_75),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_177),
.Y(n_233)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

AO22x1_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_77),
.B1(n_89),
.B2(n_58),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_179),
.A2(n_187),
.B(n_189),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_159),
.A2(n_110),
.B1(n_108),
.B2(n_104),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_180),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_123),
.A2(n_77),
.B(n_103),
.C(n_101),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_181),
.B(n_197),
.Y(n_236)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_183),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_117),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_184),
.B(n_195),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_133),
.A2(n_103),
.B1(n_67),
.B2(n_63),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_123),
.A2(n_151),
.B1(n_174),
.B2(n_133),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_188),
.B(n_206),
.Y(n_231)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_192),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_193),
.A2(n_205),
.B1(n_207),
.B2(n_217),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_136),
.A2(n_140),
.B1(n_124),
.B2(n_170),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_144),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_148),
.A2(n_147),
.B(n_118),
.C(n_169),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_198),
.Y(n_247)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_199),
.Y(n_252)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_202),
.Y(n_241)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_131),
.A2(n_153),
.B1(n_163),
.B2(n_167),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_204),
.A2(n_181),
.B1(n_227),
.B2(n_205),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_138),
.B(n_171),
.Y(n_206)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_142),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_210),
.Y(n_250)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_115),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_211),
.B(n_212),
.Y(n_268)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_126),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_116),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_213),
.B(n_214),
.Y(n_237)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_116),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_215),
.B(n_216),
.Y(n_238)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_135),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_166),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_127),
.B(n_156),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_218),
.B(n_219),
.Y(n_270)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_139),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_220),
.A2(n_205),
.B1(n_200),
.B2(n_219),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_L g222 ( 
.A1(n_137),
.A2(n_162),
.B1(n_135),
.B2(n_122),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_224),
.B1(n_227),
.B2(n_217),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_122),
.A2(n_162),
.B1(n_142),
.B2(n_127),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_127),
.B(n_139),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_225),
.B(n_226),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_165),
.A2(n_141),
.B(n_139),
.C(n_134),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g227 ( 
.A1(n_134),
.A2(n_156),
.B1(n_131),
.B2(n_137),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_161),
.A2(n_158),
.B1(n_119),
.B2(n_75),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_228),
.A2(n_192),
.B1(n_199),
.B2(n_207),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_161),
.B(n_141),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_229),
.B(n_230),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_221),
.A2(n_187),
.B1(n_193),
.B2(n_204),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_242),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_221),
.A2(n_182),
.B1(n_189),
.B2(n_208),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_190),
.B(n_223),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_254),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_249),
.B(n_260),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_251),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_190),
.B(n_191),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_190),
.B(n_201),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_257),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_186),
.B(n_203),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_222),
.A2(n_179),
.B1(n_196),
.B2(n_183),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_262),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_197),
.B(n_224),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_261),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_178),
.B(n_226),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_211),
.A2(n_215),
.B1(n_209),
.B2(n_214),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_263),
.A2(n_249),
.B1(n_235),
.B2(n_238),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_205),
.B(n_220),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_265),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_190),
.B(n_145),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_231),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_289),
.Y(n_302)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_272),
.Y(n_309)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_239),
.Y(n_273)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_239),
.Y(n_274)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_274),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_240),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_277),
.Y(n_305)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_269),
.Y(n_277)
);

AND2x6_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_236),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_281),
.Y(n_306)
);

INVx11_ASAP7_75t_L g279 ( 
.A(n_251),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_239),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_258),
.A2(n_262),
.B(n_253),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_282),
.A2(n_294),
.B(n_244),
.Y(n_313)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_285),
.B(n_288),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_258),
.A2(n_236),
.B(n_242),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_286),
.A2(n_234),
.B(n_270),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_287),
.A2(n_261),
.B1(n_233),
.B2(n_248),
.Y(n_314)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_235),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_268),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_291),
.Y(n_310)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_247),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_267),
.B(n_254),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_292),
.Y(n_303)
);

OR2x2_ASAP7_75t_SL g294 ( 
.A(n_260),
.B(n_246),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_245),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_300),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_241),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_266),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_252),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_256),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_307),
.C(n_311),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_265),
.Y(n_307)
);

AOI21xp33_ASAP7_75t_L g326 ( 
.A1(n_308),
.A2(n_286),
.B(n_299),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_264),
.C(n_259),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_282),
.A2(n_233),
.B(n_244),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_312),
.A2(n_232),
.B(n_255),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_275),
.Y(n_327)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_314),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_298),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_315),
.B(n_284),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_317),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_272),
.B(n_237),
.Y(n_319)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_319),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_250),
.C(n_266),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_298),
.C(n_293),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_326),
.B(n_308),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_327),
.B(n_320),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_310),
.C(n_304),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_311),
.A2(n_283),
.B1(n_293),
.B2(n_275),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_329),
.A2(n_311),
.B1(n_320),
.B2(n_309),
.Y(n_341)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_330),
.Y(n_340)
);

NOR3xp33_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_278),
.C(n_279),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_331),
.B(n_337),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_321),
.A2(n_248),
.B(n_295),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_334),
.A2(n_335),
.B(n_338),
.Y(n_343)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_316),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_316),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_310),
.A2(n_287),
.B1(n_296),
.B2(n_255),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_334),
.A2(n_312),
.B(n_313),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_339),
.A2(n_338),
.B(n_324),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_341),
.A2(n_332),
.B1(n_315),
.B2(n_333),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_SL g354 ( 
.A(n_342),
.B(n_336),
.C(n_303),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_329),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_347),
.C(n_348),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_304),
.C(n_307),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_306),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_302),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_350),
.C(n_322),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_294),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_300),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_352),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_290),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_354),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_355),
.A2(n_343),
.B(n_339),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_356),
.B(n_359),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_341),
.A2(n_332),
.B1(n_303),
.B2(n_333),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_357),
.B(n_347),
.C(n_348),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_360),
.B(n_361),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_357),
.B(n_344),
.C(n_349),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_355),
.B(n_345),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_363),
.A2(n_364),
.B(n_350),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_366),
.B(n_360),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_367),
.B(n_362),
.Y(n_373)
);

NAND3xp33_ASAP7_75t_L g368 ( 
.A(n_361),
.B(n_305),
.C(n_354),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_370),
.Y(n_374)
);

AOI322xp5_ASAP7_75t_L g370 ( 
.A1(n_363),
.A2(n_358),
.A3(n_356),
.B1(n_318),
.B2(n_322),
.C1(n_353),
.C2(n_323),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_371),
.A2(n_365),
.B(n_359),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_372),
.B(n_373),
.Y(n_376)
);

OA21x2_ASAP7_75t_SL g375 ( 
.A1(n_374),
.A2(n_369),
.B(n_362),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_375),
.B(n_288),
.C(n_291),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_377),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_376),
.Y(n_379)
);


endmodule