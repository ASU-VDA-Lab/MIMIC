module fake_jpeg_4486_n_185 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_185);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

INVx11_ASAP7_75t_SL g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_25),
.Y(n_40)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_0),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_29),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_22),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2x1_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_14),
.Y(n_37)
);

NOR2xp67_ASAP7_75t_R g52 ( 
.A(n_37),
.B(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_29),
.B(n_27),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_44),
.B(n_21),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_25),
.B1(n_21),
.B2(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_49),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_52),
.B(n_41),
.C(n_36),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_27),
.B1(n_31),
.B2(n_15),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_17),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_27),
.B1(n_32),
.B2(n_31),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_12),
.B1(n_17),
.B2(n_18),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_33),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_59),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_53),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_69),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_46),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_75),
.B1(n_57),
.B2(n_64),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_43),
.C(n_56),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_84),
.C(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_83),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_60),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_43),
.C(n_54),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_83),
.B1(n_73),
.B2(n_63),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_97),
.B1(n_76),
.B2(n_78),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_74),
.A2(n_69),
.B(n_45),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_91),
.C(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_70),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_98),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_92),
.B(n_62),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_94),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_48),
.B1(n_34),
.B2(n_65),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_41),
.C(n_34),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_36),
.B(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_59),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_78),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_85),
.C(n_76),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_114),
.C(n_19),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_24),
.B1(n_18),
.B2(n_16),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_112),
.C(n_105),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_59),
.Y(n_108)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_42),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_97),
.B(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_111),
.B(n_113),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_33),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_12),
.C(n_19),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_91),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_122),
.B1(n_125),
.B2(n_109),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_99),
.B(n_86),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_113),
.B1(n_109),
.B2(n_106),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_123),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_16),
.B1(n_20),
.B2(n_22),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_33),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_128),
.C(n_124),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_102),
.C(n_105),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_131),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_101),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_20),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_136),
.C(n_141),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_20),
.B1(n_0),
.B2(n_1),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_127),
.C(n_117),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_28),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_142),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_140),
.B(n_1),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_119),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_30),
.C(n_23),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_133),
.A2(n_8),
.B(n_2),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_145),
.B(n_146),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_136),
.A2(n_8),
.B(n_2),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_150),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_30),
.B(n_1),
.Y(n_148)
);

OAI21x1_ASAP7_75t_SL g156 ( 
.A1(n_148),
.A2(n_9),
.B(n_3),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_141),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_153),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_139),
.A2(n_7),
.B(n_3),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_154),
.A2(n_156),
.B(n_161),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_142),
.B1(n_138),
.B2(n_39),
.Y(n_155)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_138),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_162),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_23),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_23),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_160),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_164),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_149),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_39),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_165),
.B(n_6),
.Y(n_172)
);

AOI31xp33_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_9),
.A3(n_4),
.B(n_5),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_170),
.Y(n_173)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_172),
.B(n_7),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_23),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_175),
.C(n_176),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_1),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_7),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_177),
.B(n_178),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_166),
.C(n_39),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_180),
.A2(n_10),
.B(n_11),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_166),
.B(n_10),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_183),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_181),
.Y(n_185)
);


endmodule