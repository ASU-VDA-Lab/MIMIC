module fake_jpeg_30860_n_140 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx8_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_19),
.Y(n_35)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_35),
.Y(n_50)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_8),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_22),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_53),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_21),
.B(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_52),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_25),
.B1(n_15),
.B2(n_17),
.Y(n_51)
);

NOR2xp67_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_35),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_61),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_23),
.B1(n_27),
.B2(n_16),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_24),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_35),
.A2(n_23),
.B1(n_24),
.B2(n_17),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_63),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_20),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_29),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_71),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_21),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_10),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_73),
.B(n_77),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_58),
.B1(n_52),
.B2(n_47),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_56),
.B1(n_54),
.B2(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_34),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_34),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_42),
.A3(n_38),
.B1(n_36),
.B2(n_9),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_50),
.Y(n_88)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_55),
.B1(n_56),
.B2(n_62),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_86),
.B1(n_90),
.B2(n_91),
.Y(n_106)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_67),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_44),
.B1(n_50),
.B2(n_42),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_44),
.B1(n_50),
.B2(n_42),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_38),
.B1(n_1),
.B2(n_2),
.Y(n_94)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_101),
.C(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_103),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_105),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_75),
.B(n_78),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_96),
.A2(n_64),
.B1(n_80),
.B2(n_65),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_104),
.B1(n_107),
.B2(n_101),
.Y(n_118)
);

NOR4xp25_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_75),
.C(n_81),
.D(n_11),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_86),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_80),
.Y(n_107)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_91),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_111),
.B(n_115),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_83),
.B1(n_92),
.B2(n_82),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_118),
.B1(n_102),
.B2(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

AO221x1_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_92),
.B1(n_77),
.B2(n_76),
.C(n_113),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_98),
.C(n_105),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_123),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_120),
.Y(n_126)
);

AO221x1_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_109),
.B1(n_93),
.B2(n_87),
.C(n_84),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_125),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_84),
.C(n_38),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_121),
.A2(n_111),
.B1(n_110),
.B2(n_4),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_130),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_110),
.B1(n_8),
.B2(n_11),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_125),
.C(n_119),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_132),
.B(n_133),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_0),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_12),
.C(n_3),
.Y(n_133)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_130),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_135),
.B(n_134),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_126),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g139 ( 
.A(n_137),
.B(n_138),
.C(n_0),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_4),
.Y(n_140)
);


endmodule