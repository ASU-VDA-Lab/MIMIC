module fake_netlist_6_3005_n_1951 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1951);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1951;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_62),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_48),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_59),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_122),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_166),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_73),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_27),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_86),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_71),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_136),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_6),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_61),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_27),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_117),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_83),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_100),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_109),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_64),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_101),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_91),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_41),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_50),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_9),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_61),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_76),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_60),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_73),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_108),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_70),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_24),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_8),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_185),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_65),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_156),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_139),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_138),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_44),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_113),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_103),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_2),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_158),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_130),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_4),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_81),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_97),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_10),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_34),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_167),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_114),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_6),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_92),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_37),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_22),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_133),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_186),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_169),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_94),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_28),
.Y(n_257)
);

BUFx8_ASAP7_75t_SL g258 ( 
.A(n_29),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_93),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_127),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_172),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_1),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_43),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_110),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_187),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_43),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_47),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_105),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_98),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_38),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_30),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_148),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_104),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_69),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_66),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_126),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_63),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_78),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_24),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_45),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_80),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_85),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_34),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_29),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_0),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_191),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_53),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_54),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_2),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_49),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_3),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_164),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_70),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_79),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_36),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_134),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_68),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_68),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_175),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_10),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_58),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_48),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_53),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_88),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_178),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_121),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_28),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_36),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_12),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_19),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_189),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_0),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_132),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_174),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_131),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_173),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_90),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_64),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_152),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_55),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_58),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_45),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_57),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_12),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_33),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_118),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_119),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_95),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_1),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_65),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_112),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_40),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_163),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_155),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_190),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_77),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_128),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_69),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_145),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_51),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_165),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_15),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_30),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_150),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_171),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_59),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_57),
.Y(n_347)
);

BUFx10_ASAP7_75t_L g348 ( 
.A(n_39),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_125),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_18),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_37),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_71),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_153),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_87),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_102),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_160),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_135),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_4),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_116),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_141),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_182),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_143),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_99),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_7),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_39),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_84),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_54),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_38),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_170),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_176),
.Y(n_370)
);

BUFx10_ASAP7_75t_L g371 ( 
.A(n_17),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_115),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_32),
.Y(n_373)
);

BUFx10_ASAP7_75t_L g374 ( 
.A(n_162),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_31),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_16),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_74),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_9),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_96),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_180),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_47),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_63),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_192),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_82),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_123),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_199),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_234),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_258),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_239),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_208),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_224),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_242),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_246),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_224),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_247),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_224),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_224),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_224),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_227),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_236),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_249),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_227),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_254),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_255),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_227),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_199),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_260),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_356),
.B(n_3),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_227),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_287),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_287),
.Y(n_411)
);

INVxp33_ASAP7_75t_L g412 ( 
.A(n_194),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_265),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_269),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_272),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_227),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_356),
.B(n_5),
.Y(n_417)
);

INVxp33_ASAP7_75t_SL g418 ( 
.A(n_193),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_273),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_250),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_250),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_217),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_250),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_281),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_282),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_372),
.B(n_5),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_250),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_250),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_218),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_209),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_278),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_286),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_330),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_193),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_210),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_330),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_236),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_330),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_330),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_304),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_305),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_311),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_330),
.Y(n_443)
);

INVxp33_ASAP7_75t_SL g444 ( 
.A(n_196),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_287),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_363),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_296),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_199),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_238),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_334),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_238),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_245),
.Y(n_452)
);

INVxp33_ASAP7_75t_SL g453 ( 
.A(n_196),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_245),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_284),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_316),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_349),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_348),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_360),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_384),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_284),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_288),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_244),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_252),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_257),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_197),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_288),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_334),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_277),
.B(n_7),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_323),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_323),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_325),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_197),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_198),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_198),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_325),
.Y(n_476)
);

NOR2xp67_ASAP7_75t_L g477 ( 
.A(n_364),
.B(n_8),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_209),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_262),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_216),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_267),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_372),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_391),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_430),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_202),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_417),
.B(n_380),
.Y(n_487)
);

AND3x2_ASAP7_75t_L g488 ( 
.A(n_408),
.B(n_370),
.C(n_315),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_394),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_434),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_394),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_430),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_426),
.B(n_387),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_430),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_396),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_468),
.B(n_202),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_396),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_386),
.B(n_315),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_SL g499 ( 
.A(n_412),
.B(n_280),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_397),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_430),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_397),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_406),
.B(n_205),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_430),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_450),
.B(n_205),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_478),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_478),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_478),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_478),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_398),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_478),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_448),
.B(n_370),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_418),
.B(n_203),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_398),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_448),
.B(n_280),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_399),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_399),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_402),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_402),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_405),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_405),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_409),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_409),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_400),
.B(n_290),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_437),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_416),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_416),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_420),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_457),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_420),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_421),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_421),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_435),
.A2(n_318),
.B1(n_300),
.B2(n_308),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_423),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_423),
.B(n_211),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_427),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_389),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_427),
.B(n_211),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_428),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_R g541 ( 
.A(n_444),
.B(n_201),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_428),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_433),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_433),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_455),
.Y(n_545)
);

AND3x2_ASAP7_75t_L g546 ( 
.A(n_410),
.B(n_445),
.C(n_411),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_436),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_436),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_437),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_438),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_438),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_439),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_453),
.B(n_463),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_439),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_443),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_443),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g557 ( 
.A(n_464),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_455),
.B(n_209),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_480),
.B(n_212),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_449),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_507),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_515),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_558),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_515),
.Y(n_564)
);

AND2x2_ASAP7_75t_SL g565 ( 
.A(n_487),
.B(n_209),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_515),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_515),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_517),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_558),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_487),
.B(n_498),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_517),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_514),
.B(n_392),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_514),
.B(n_393),
.Y(n_573)
);

OAI22xp33_ASAP7_75t_L g574 ( 
.A1(n_490),
.A2(n_541),
.B1(n_503),
.B2(n_303),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_558),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_494),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_503),
.B(n_395),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_538),
.B(n_387),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_505),
.B(n_401),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_494),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_493),
.B(n_469),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_553),
.B(n_403),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_517),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_494),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_498),
.A2(n_320),
.B1(n_290),
.B2(n_222),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_534),
.B(n_390),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_517),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_498),
.B(n_404),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_507),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_526),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_494),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_520),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_525),
.A2(n_320),
.B1(n_225),
.B2(n_231),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_558),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_505),
.B(n_407),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_558),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_520),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_520),
.Y(n_598)
);

AND2x6_ASAP7_75t_L g599 ( 
.A(n_513),
.B(n_209),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_520),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_494),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_526),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_494),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_558),
.Y(n_604)
);

AND2x2_ASAP7_75t_SL g605 ( 
.A(n_557),
.B(n_215),
.Y(n_605)
);

NAND3xp33_ASAP7_75t_L g606 ( 
.A(n_490),
.B(n_479),
.C(n_465),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_486),
.B(n_413),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_493),
.B(n_414),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_483),
.Y(n_609)
);

BUFx4f_ASAP7_75t_L g610 ( 
.A(n_513),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_494),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_494),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_525),
.A2(n_219),
.B1(n_263),
.B2(n_248),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_525),
.B(n_449),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_483),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_534),
.B(n_422),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_549),
.Y(n_617)
);

AND2x2_ASAP7_75t_SL g618 ( 
.A(n_557),
.B(n_215),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_L g619 ( 
.A1(n_541),
.A2(n_342),
.B1(n_347),
.B2(n_266),
.Y(n_619)
);

INVxp67_ASAP7_75t_SL g620 ( 
.A(n_549),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_486),
.B(n_415),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_553),
.B(n_419),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_496),
.B(n_424),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_483),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_494),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_501),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_501),
.Y(n_627)
);

AND2x6_ASAP7_75t_L g628 ( 
.A(n_513),
.B(n_215),
.Y(n_628)
);

INVxp67_ASAP7_75t_SL g629 ( 
.A(n_536),
.Y(n_629)
);

NAND3xp33_ASAP7_75t_L g630 ( 
.A(n_559),
.B(n_481),
.C(n_440),
.Y(n_630)
);

BUFx10_ASAP7_75t_L g631 ( 
.A(n_530),
.Y(n_631)
);

INVx5_ASAP7_75t_L g632 ( 
.A(n_501),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_485),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_516),
.A2(n_302),
.B1(n_338),
.B2(n_329),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_485),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_485),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_521),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_496),
.B(n_425),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_501),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_L g640 ( 
.A(n_559),
.B(n_456),
.C(n_442),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_489),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_521),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_489),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_489),
.Y(n_644)
);

AND3x2_ASAP7_75t_L g645 ( 
.A(n_557),
.B(n_458),
.C(n_200),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_516),
.A2(n_346),
.B1(n_381),
.B2(n_373),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_491),
.Y(n_647)
);

BUFx6f_ASAP7_75t_SL g648 ( 
.A(n_560),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_488),
.B(n_459),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_491),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_516),
.B(n_560),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_501),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_488),
.B(n_240),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_499),
.B(n_466),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_530),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_521),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_491),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_495),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_495),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_501),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_536),
.B(n_215),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_499),
.A2(n_475),
.B1(n_474),
.B2(n_473),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_495),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_539),
.B(n_253),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_497),
.Y(n_665)
);

AND2x6_ASAP7_75t_L g666 ( 
.A(n_482),
.B(n_215),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_539),
.B(n_447),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_482),
.B(n_477),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_521),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_528),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_497),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_501),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_501),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_545),
.B(n_264),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_528),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_545),
.B(n_294),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_497),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_545),
.B(n_460),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_528),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_528),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_545),
.B(n_388),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_560),
.B(n_377),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_546),
.A2(n_429),
.B1(n_446),
.B2(n_441),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_500),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_546),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_545),
.B(n_480),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_500),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_500),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_545),
.B(n_299),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_502),
.B(n_431),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_529),
.Y(n_691)
);

INVx4_ASAP7_75t_L g692 ( 
.A(n_501),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_502),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_502),
.A2(n_352),
.B1(n_382),
.B2(n_336),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_529),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_511),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_511),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_511),
.B(n_261),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_535),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_529),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_518),
.B(n_379),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_518),
.B(n_451),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_518),
.B(n_451),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_519),
.B(n_432),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_535),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_529),
.Y(n_706)
);

CKINVDCx16_ASAP7_75t_R g707 ( 
.A(n_519),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_535),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_535),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_519),
.B(n_452),
.Y(n_710)
);

AND2x6_ASAP7_75t_L g711 ( 
.A(n_522),
.B(n_336),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_522),
.A2(n_233),
.B1(n_230),
.B2(n_383),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_522),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_605),
.B(n_212),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_609),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_629),
.B(n_527),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_565),
.B(n_527),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_609),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_565),
.B(n_527),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_577),
.B(n_531),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_572),
.B(n_573),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_563),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_579),
.B(n_595),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_623),
.B(n_531),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_570),
.B(n_531),
.Y(n_725)
);

INVx8_ASAP7_75t_L g726 ( 
.A(n_648),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_561),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_608),
.B(n_230),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_615),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_605),
.B(n_233),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_615),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_624),
.Y(n_732)
);

NOR3xp33_ASAP7_75t_SL g733 ( 
.A(n_619),
.B(n_204),
.C(n_201),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_607),
.B(n_326),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_618),
.B(n_610),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_618),
.B(n_326),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_563),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_569),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_624),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_610),
.B(n_328),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_633),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_633),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_569),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_635),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_635),
.Y(n_745)
);

NAND2x1p5_ASAP7_75t_L g746 ( 
.A(n_610),
.B(n_195),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_664),
.B(n_533),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_621),
.B(n_328),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_636),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_575),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_575),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_707),
.B(n_331),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_707),
.B(n_331),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_617),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_588),
.B(n_533),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_594),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_638),
.A2(n_213),
.B1(n_214),
.B2(n_223),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_561),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_590),
.B(n_337),
.Y(n_759)
);

AND2x4_ASAP7_75t_SL g760 ( 
.A(n_631),
.B(n_261),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_651),
.A2(n_237),
.B1(n_232),
.B2(n_226),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_620),
.B(n_337),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_590),
.B(n_339),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_SL g764 ( 
.A(n_648),
.B(n_241),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_651),
.A2(n_251),
.B1(n_319),
.B2(n_333),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_589),
.Y(n_766)
);

NOR2xp67_ASAP7_75t_L g767 ( 
.A(n_606),
.B(n_339),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_602),
.B(n_341),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_636),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_614),
.B(n_533),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_696),
.B(n_540),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_696),
.B(n_540),
.Y(n_772)
);

NAND3xp33_ASAP7_75t_L g773 ( 
.A(n_690),
.B(n_271),
.C(n_270),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_614),
.B(n_540),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_589),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_581),
.A2(n_341),
.B1(n_344),
.B2(n_353),
.Y(n_776)
);

NAND2x1_ASAP7_75t_L g777 ( 
.A(n_591),
.B(n_523),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_602),
.B(n_344),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_581),
.A2(n_243),
.B1(n_256),
.B2(n_259),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_686),
.B(n_594),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_617),
.B(n_353),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_682),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_686),
.B(n_547),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_580),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_686),
.B(n_547),
.Y(n_785)
);

NOR2xp67_ASAP7_75t_L g786 ( 
.A(n_630),
.B(n_354),
.Y(n_786)
);

O2A1O1Ixp5_ASAP7_75t_L g787 ( 
.A1(n_596),
.A2(n_556),
.B(n_547),
.C(n_548),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_596),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_674),
.A2(n_492),
.B(n_484),
.Y(n_789)
);

OAI22xp33_ASAP7_75t_L g790 ( 
.A1(n_581),
.A2(n_327),
.B1(n_268),
.B2(n_292),
.Y(n_790)
);

NOR3xp33_ASAP7_75t_L g791 ( 
.A(n_574),
.B(n_275),
.C(n_274),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_641),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_604),
.A2(n_357),
.B1(n_276),
.B2(n_306),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_604),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_581),
.A2(n_366),
.B1(n_369),
.B2(n_361),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_655),
.Y(n_796)
);

OAI221xp5_ASAP7_75t_L g797 ( 
.A1(n_585),
.A2(n_335),
.B1(n_313),
.B2(n_314),
.C(n_317),
.Y(n_797)
);

BUFx12f_ASAP7_75t_SL g798 ( 
.A(n_668),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_687),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_641),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_643),
.A2(n_359),
.B1(n_355),
.B2(n_385),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_643),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_640),
.B(n_354),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_697),
.B(n_548),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_682),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_644),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_697),
.B(n_548),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_668),
.A2(n_369),
.B1(n_361),
.B2(n_362),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_644),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_704),
.B(n_362),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_599),
.B(n_336),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_668),
.A2(n_383),
.B1(n_366),
.B2(n_376),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_647),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_653),
.B(n_261),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_676),
.B(n_550),
.Y(n_815)
);

AOI221xp5_ASAP7_75t_L g816 ( 
.A1(n_634),
.A2(n_646),
.B1(n_343),
.B2(n_340),
.C(n_378),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_582),
.B(n_279),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_647),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_650),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_650),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_657),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_657),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_SL g823 ( 
.A(n_631),
.B(n_345),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_658),
.Y(n_824)
);

AND2x6_ASAP7_75t_SL g825 ( 
.A(n_649),
.B(n_452),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_655),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_681),
.B(n_701),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_622),
.B(n_283),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_667),
.B(n_204),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_685),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_658),
.A2(n_336),
.B1(n_556),
.B2(n_550),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_689),
.B(n_550),
.Y(n_832)
);

OAI22xp33_ASAP7_75t_L g833 ( 
.A1(n_668),
.A2(n_712),
.B1(n_662),
.B2(n_685),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_L g834 ( 
.A(n_599),
.B(n_336),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_631),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_648),
.A2(n_556),
.B1(n_551),
.B2(n_322),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_678),
.B(n_206),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_645),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_654),
.B(n_285),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_698),
.B(n_345),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_659),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_659),
.B(n_551),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_663),
.B(n_665),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_580),
.Y(n_844)
);

INVx4_ASAP7_75t_L g845 ( 
.A(n_580),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_578),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_663),
.B(n_289),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_665),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_671),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_702),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_703),
.B(n_551),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_671),
.B(n_523),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_677),
.B(n_523),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_677),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_684),
.B(n_523),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_684),
.B(n_523),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_688),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_702),
.B(n_454),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_613),
.B(n_345),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_688),
.B(n_523),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_693),
.B(n_713),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_661),
.A2(n_584),
.B(n_576),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_580),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_703),
.B(n_454),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_580),
.Y(n_865)
);

NAND2xp33_ASAP7_75t_L g866 ( 
.A(n_599),
.B(n_206),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_593),
.A2(n_321),
.B1(n_291),
.B2(n_293),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_693),
.B(n_524),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_627),
.Y(n_869)
);

NOR2x1p5_ASAP7_75t_L g870 ( 
.A(n_586),
.B(n_207),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_713),
.A2(n_555),
.B1(n_554),
.B2(n_552),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_702),
.B(n_374),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_599),
.A2(n_555),
.B1(n_554),
.B2(n_552),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_562),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_586),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_562),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_710),
.B(n_374),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_710),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_683),
.B(n_374),
.Y(n_879)
);

AND2x2_ASAP7_75t_SL g880 ( 
.A(n_661),
.B(n_461),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_616),
.B(n_295),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_564),
.Y(n_882)
);

INVx8_ASAP7_75t_L g883 ( 
.A(n_599),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_576),
.B(n_524),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_564),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_566),
.B(n_461),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_723),
.B(n_576),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_721),
.A2(n_584),
.B(n_601),
.C(n_603),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_782),
.B(n_616),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_717),
.A2(n_601),
.B(n_584),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_728),
.B(n_601),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_727),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_734),
.A2(n_652),
.B(n_603),
.C(n_625),
.Y(n_893)
);

AOI21x1_ASAP7_75t_L g894 ( 
.A1(n_777),
.A2(n_567),
.B(n_566),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_720),
.B(n_603),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_719),
.A2(n_652),
.B(n_625),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_845),
.A2(n_626),
.B(n_591),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_743),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_780),
.A2(n_652),
.B(n_625),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_735),
.A2(n_694),
.B1(n_660),
.B2(n_673),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_724),
.B(n_755),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_715),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_782),
.B(n_805),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_826),
.Y(n_904)
);

INVx11_ASAP7_75t_L g905 ( 
.A(n_835),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_748),
.B(n_660),
.Y(n_906)
);

OAI21xp33_ASAP7_75t_L g907 ( 
.A1(n_781),
.A2(n_220),
.B(n_207),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_747),
.B(n_660),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_845),
.A2(n_626),
.B(n_591),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_845),
.A2(n_692),
.B(n_626),
.Y(n_910)
);

O2A1O1Ixp33_ASAP7_75t_SL g911 ( 
.A1(n_714),
.A2(n_675),
.B(n_567),
.C(n_568),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_725),
.B(n_673),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_878),
.A2(n_673),
.B1(n_692),
.B2(n_627),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_878),
.B(n_692),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_784),
.A2(n_672),
.B(n_627),
.Y(n_915)
);

AO21x1_ASAP7_75t_L g916 ( 
.A1(n_746),
.A2(n_709),
.B(n_571),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_805),
.B(n_348),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_715),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_862),
.A2(n_571),
.B(n_568),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_727),
.B(n_462),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_830),
.Y(n_921)
);

AOI33xp33_ASAP7_75t_L g922 ( 
.A1(n_816),
.A2(n_470),
.A3(n_462),
.B1(n_467),
.B2(n_471),
.B3(n_472),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_754),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_750),
.A2(n_627),
.B1(n_672),
.B2(n_598),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_784),
.A2(n_672),
.B(n_627),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_784),
.A2(n_672),
.B(n_709),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_784),
.A2(n_672),
.B(n_709),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_827),
.A2(n_599),
.B1(n_628),
.B2(n_666),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_770),
.B(n_583),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_SL g930 ( 
.A(n_798),
.B(n_348),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_830),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_758),
.B(n_371),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_817),
.A2(n_669),
.B(n_597),
.C(n_706),
.Y(n_933)
);

NAND2x1_ASAP7_75t_L g934 ( 
.A(n_784),
.B(n_699),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_750),
.A2(n_669),
.B1(n_597),
.B2(n_706),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_844),
.A2(n_612),
.B(n_611),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_804),
.A2(n_637),
.B(n_700),
.C(n_695),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_844),
.A2(n_612),
.B(n_611),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_718),
.Y(n_939)
);

AO21x1_ASAP7_75t_L g940 ( 
.A1(n_746),
.A2(n_587),
.B(n_583),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_807),
.B(n_297),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_770),
.B(n_587),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_844),
.A2(n_611),
.B(n_612),
.Y(n_943)
);

BUFx4f_ASAP7_75t_L g944 ( 
.A(n_726),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_774),
.B(n_592),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_833),
.B(n_850),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_828),
.A2(n_598),
.B(n_600),
.C(n_592),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_844),
.A2(n_611),
.B(n_632),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_799),
.B(n_298),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_844),
.A2(n_611),
.B(n_632),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_865),
.A2(n_785),
.B(n_783),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_774),
.B(n_600),
.Y(n_952)
);

AOI22x1_ASAP7_75t_L g953 ( 
.A1(n_751),
.A2(n_679),
.B1(n_656),
.B2(n_642),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_839),
.A2(n_637),
.B(n_642),
.C(n_656),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_850),
.Y(n_955)
);

OAI22x1_ASAP7_75t_L g956 ( 
.A1(n_881),
.A2(n_235),
.B1(n_220),
.B2(n_221),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_716),
.B(n_670),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_722),
.A2(n_738),
.B1(n_756),
.B2(n_737),
.Y(n_958)
);

CKINVDCx10_ASAP7_75t_R g959 ( 
.A(n_826),
.Y(n_959)
);

OAI21xp33_ASAP7_75t_L g960 ( 
.A1(n_823),
.A2(n_235),
.B(n_221),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_758),
.B(n_699),
.Y(n_961)
);

AOI21xp33_ASAP7_75t_L g962 ( 
.A1(n_837),
.A2(n_301),
.B(n_307),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_766),
.B(n_699),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_851),
.A2(n_599),
.B1(n_628),
.B2(n_666),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_851),
.B(n_670),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_766),
.B(n_699),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_865),
.A2(n_632),
.B(n_612),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_852),
.A2(n_680),
.B(n_700),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_865),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_864),
.B(n_675),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_865),
.A2(n_612),
.B(n_632),
.Y(n_971)
);

AOI21x1_ASAP7_75t_L g972 ( 
.A1(n_777),
.A2(n_680),
.B(n_679),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_746),
.A2(n_691),
.B1(n_695),
.B2(n_309),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_865),
.A2(n_632),
.B(n_639),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_800),
.A2(n_324),
.B(n_229),
.C(n_332),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_864),
.B(n_691),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_853),
.A2(n_628),
.B(n_666),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_847),
.A2(n_312),
.B(n_310),
.C(n_542),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_759),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_800),
.A2(n_332),
.B(n_324),
.C(n_229),
.Y(n_980)
);

BUFx12f_ASAP7_75t_L g981 ( 
.A(n_825),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_775),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_729),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_815),
.A2(n_832),
.B(n_843),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_809),
.B(n_628),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_809),
.B(n_628),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_775),
.B(n_699),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_829),
.B(n_228),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_730),
.A2(n_524),
.B(n_542),
.C(n_544),
.Y(n_989)
);

NOR3xp33_ASAP7_75t_L g990 ( 
.A(n_875),
.B(n_343),
.C(n_228),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_731),
.B(n_705),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_861),
.A2(n_639),
.B(n_708),
.Y(n_992)
);

CKINVDCx6p67_ASAP7_75t_R g993 ( 
.A(n_835),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_846),
.B(n_340),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_813),
.B(n_628),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_855),
.A2(n_628),
.B(n_666),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_813),
.Y(n_997)
);

O2A1O1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_736),
.A2(n_542),
.B(n_524),
.C(n_544),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_856),
.A2(n_666),
.B(n_484),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_771),
.A2(n_639),
.B(n_708),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_732),
.B(n_705),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_739),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_739),
.B(n_705),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_858),
.Y(n_1004)
);

NAND2xp33_ASAP7_75t_L g1005 ( 
.A(n_726),
.B(n_666),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_837),
.B(n_350),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_726),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_741),
.B(n_705),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_772),
.A2(n_639),
.B(n_708),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_819),
.B(n_820),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_741),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_788),
.Y(n_1012)
);

AOI21x1_ASAP7_75t_L g1013 ( 
.A1(n_842),
.A2(n_492),
.B(n_504),
.Y(n_1013)
);

AOI21xp33_ASAP7_75t_L g1014 ( 
.A1(n_829),
.A2(n_350),
.B(n_351),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_810),
.B(n_351),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_819),
.B(n_705),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_884),
.A2(n_639),
.B(n_708),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_883),
.A2(n_708),
.B(n_508),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_794),
.A2(n_666),
.B1(n_711),
.B2(n_524),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_742),
.B(n_535),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_752),
.B(n_358),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_883),
.A2(n_789),
.B(n_863),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_820),
.B(n_524),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_824),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_883),
.A2(n_506),
.B(n_484),
.Y(n_1025)
);

INVx3_ASAP7_75t_SL g1026 ( 
.A(n_796),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_753),
.B(n_358),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_883),
.A2(n_506),
.B(n_484),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_863),
.A2(n_508),
.B(n_492),
.Y(n_1029)
);

OAI21xp33_ASAP7_75t_L g1030 ( 
.A1(n_762),
.A2(n_367),
.B(n_378),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_863),
.A2(n_508),
.B(n_492),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_824),
.B(n_542),
.Y(n_1032)
);

INVxp67_ASAP7_75t_L g1033 ( 
.A(n_763),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_SL g1034 ( 
.A(n_798),
.B(n_726),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_869),
.A2(n_740),
.B(n_860),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_744),
.B(n_535),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_841),
.A2(n_375),
.B(n_365),
.C(n_368),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_841),
.B(n_542),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_848),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_796),
.Y(n_1040)
);

CKINVDCx8_ASAP7_75t_R g1041 ( 
.A(n_838),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_848),
.B(n_857),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_857),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_858),
.B(n_467),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_869),
.A2(n_509),
.B(n_504),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_812),
.B(n_365),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_744),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_745),
.A2(n_367),
.B1(n_375),
.B2(n_368),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_869),
.A2(n_512),
.B(n_508),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_745),
.Y(n_1050)
);

NOR2xp67_ASAP7_75t_L g1051 ( 
.A(n_773),
.B(n_75),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_760),
.B(n_371),
.Y(n_1052)
);

OR2x6_ASAP7_75t_L g1053 ( 
.A(n_838),
.B(n_470),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_868),
.A2(n_506),
.B(n_509),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_858),
.B(n_471),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_776),
.B(n_11),
.Y(n_1056)
);

AOI21x1_ASAP7_75t_L g1057 ( 
.A1(n_885),
.A2(n_506),
.B(n_512),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_749),
.A2(n_509),
.B(n_504),
.Y(n_1058)
);

NOR2x1_ASAP7_75t_L g1059 ( 
.A(n_786),
.B(n_767),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_749),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_769),
.B(n_792),
.Y(n_1061)
);

AOI21x1_ASAP7_75t_L g1062 ( 
.A1(n_885),
.A2(n_504),
.B(n_510),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_769),
.A2(n_510),
.B(n_512),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_792),
.A2(n_822),
.B(n_821),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_802),
.A2(n_510),
.B(n_512),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_802),
.B(n_542),
.Y(n_1066)
);

O2A1O1Ixp5_ASAP7_75t_L g1067 ( 
.A1(n_806),
.A2(n_510),
.B(n_509),
.C(n_544),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_806),
.B(n_544),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_818),
.B(n_821),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_818),
.A2(n_544),
.B1(n_555),
.B2(n_554),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_822),
.B(n_544),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_849),
.B(n_532),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_849),
.B(n_535),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_SL g1074 ( 
.A1(n_946),
.A2(n_803),
.B(n_814),
.C(n_757),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_898),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_901),
.A2(n_854),
.B1(n_761),
.B2(n_765),
.Y(n_1076)
);

A2O1A1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_1015),
.A2(n_795),
.B(n_779),
.C(n_733),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_946),
.A2(n_872),
.B1(n_764),
.B2(n_877),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1006),
.B(n_870),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_978),
.A2(n_854),
.B(n_790),
.C(n_787),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_931),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_993),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_983),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_941),
.B(n_921),
.Y(n_1084)
);

BUFx4f_ASAP7_75t_L g1085 ( 
.A(n_1026),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_1004),
.B(n_764),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_1007),
.B(n_840),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_984),
.A2(n_882),
.B(n_880),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_1056),
.A2(n_791),
.B1(n_797),
.B2(n_886),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_1010),
.A2(n_836),
.B(n_866),
.C(n_886),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_1040),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_941),
.B(n_768),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1014),
.B(n_778),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1042),
.A2(n_866),
.B(n_859),
.C(n_876),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_1015),
.A2(n_760),
.B(n_880),
.C(n_879),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_969),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1056),
.A2(n_867),
.B1(n_834),
.B2(n_811),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_891),
.A2(n_834),
.B(n_811),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1006),
.B(n_889),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_983),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1012),
.B(n_874),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_923),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_917),
.B(n_808),
.Y(n_1103)
);

AO32x2_ASAP7_75t_L g1104 ( 
.A1(n_924),
.A2(n_935),
.A3(n_900),
.B1(n_973),
.B2(n_913),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_1021),
.A2(n_876),
.B(n_874),
.C(n_793),
.Y(n_1105)
);

INVxp67_ASAP7_75t_L g1106 ( 
.A(n_923),
.Y(n_1106)
);

NOR2x1_ASAP7_75t_L g1107 ( 
.A(n_1007),
.B(n_472),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_906),
.A2(n_873),
.B(n_831),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_912),
.A2(n_951),
.B(n_909),
.Y(n_1109)
);

CKINVDCx14_ASAP7_75t_R g1110 ( 
.A(n_904),
.Y(n_1110)
);

NOR2x1_ASAP7_75t_L g1111 ( 
.A(n_1059),
.B(n_955),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1012),
.B(n_801),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_903),
.B(n_371),
.Y(n_1113)
);

BUFx10_ASAP7_75t_L g1114 ( 
.A(n_1021),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_887),
.B(n_871),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_897),
.A2(n_555),
.B(n_554),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_1026),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_910),
.A2(n_552),
.B(n_537),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_969),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_1027),
.A2(n_476),
.B(n_537),
.C(n_532),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_982),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_969),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_958),
.A2(n_552),
.B1(n_537),
.B2(n_532),
.Y(n_1123)
);

CKINVDCx8_ASAP7_75t_R g1124 ( 
.A(n_959),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_SL g1125 ( 
.A1(n_1046),
.A2(n_476),
.B1(n_13),
.B2(n_14),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_1053),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_1041),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1011),
.Y(n_1128)
);

AOI21xp33_ASAP7_75t_L g1129 ( 
.A1(n_1046),
.A2(n_11),
.B(n_13),
.Y(n_1129)
);

AOI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1061),
.A2(n_537),
.B(n_532),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_920),
.B(n_997),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_905),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_920),
.B(n_711),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_888),
.A2(n_711),
.B(n_543),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1024),
.A2(n_535),
.B1(n_543),
.B2(n_144),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_903),
.B(n_14),
.Y(n_1136)
);

O2A1O1Ixp5_ASAP7_75t_L g1137 ( 
.A1(n_940),
.A2(n_711),
.B(n_188),
.C(n_183),
.Y(n_1137)
);

OAI21xp33_ASAP7_75t_SL g1138 ( 
.A1(n_1039),
.A2(n_15),
.B(n_16),
.Y(n_1138)
);

NAND2x1p5_ASAP7_75t_L g1139 ( 
.A(n_944),
.B(n_535),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_SL g1140 ( 
.A1(n_981),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_979),
.B(n_20),
.Y(n_1141)
);

NAND2xp33_ASAP7_75t_L g1142 ( 
.A(n_1043),
.B(n_711),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_929),
.A2(n_942),
.B1(n_945),
.B2(n_952),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_892),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_982),
.B(n_711),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1047),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_902),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_932),
.B(n_20),
.Y(n_1148)
);

NOR2x1_ASAP7_75t_R g1149 ( 
.A(n_1052),
.B(n_543),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1050),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_892),
.B(n_543),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_918),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_994),
.B(n_949),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1060),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_894),
.A2(n_140),
.B(n_168),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_965),
.A2(n_543),
.B1(n_161),
.B2(n_159),
.Y(n_1156)
);

INVxp67_ASAP7_75t_SL g1157 ( 
.A(n_970),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_939),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_976),
.A2(n_543),
.B1(n_157),
.B2(n_151),
.Y(n_1159)
);

O2A1O1Ixp5_ASAP7_75t_SL g1160 ( 
.A1(n_962),
.A2(n_1061),
.B(n_1069),
.C(n_966),
.Y(n_1160)
);

INVx3_ASAP7_75t_SL g1161 ( 
.A(n_1053),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_975),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_955),
.Y(n_1163)
);

OAI22x1_ASAP7_75t_L g1164 ( 
.A1(n_1027),
.A2(n_21),
.B1(n_23),
.B2(n_25),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1044),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1022),
.A2(n_895),
.B(n_957),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_899),
.A2(n_543),
.B(n_147),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_908),
.B(n_543),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_944),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_1053),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1033),
.B(n_25),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_926),
.A2(n_543),
.B(n_142),
.Y(n_1172)
);

AND2x2_ASAP7_75t_SL g1173 ( 
.A(n_1005),
.B(n_137),
.Y(n_1173)
);

NOR2x1_ASAP7_75t_L g1174 ( 
.A(n_1051),
.B(n_129),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_SL g1175 ( 
.A1(n_994),
.A2(n_124),
.B(n_120),
.C(n_111),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1002),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_1176)
);

OAI22x1_ASAP7_75t_L g1177 ( 
.A1(n_988),
.A2(n_26),
.B1(n_33),
.B2(n_35),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_927),
.A2(n_107),
.B(n_106),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_914),
.A2(n_89),
.B1(n_40),
.B2(n_41),
.Y(n_1179)
);

BUFx5_ASAP7_75t_L g1180 ( 
.A(n_1044),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_890),
.A2(n_35),
.B(n_42),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1055),
.B(n_42),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1055),
.B(n_44),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_922),
.B(n_46),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_975),
.B(n_46),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_907),
.B(n_1030),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_896),
.A2(n_49),
.B(n_50),
.Y(n_1187)
);

INVx5_ASAP7_75t_L g1188 ( 
.A(n_916),
.Y(n_1188)
);

BUFx8_ASAP7_75t_L g1189 ( 
.A(n_1034),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_953),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_930),
.B(n_51),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_949),
.B(n_52),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1069),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_960),
.B(n_52),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1064),
.A2(n_1035),
.B(n_998),
.C(n_989),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1072),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_956),
.B(n_55),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_990),
.A2(n_74),
.B1(n_60),
.B2(n_62),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_980),
.B(n_56),
.Y(n_1199)
);

INVx4_ASAP7_75t_L g1200 ( 
.A(n_934),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_915),
.A2(n_56),
.B(n_66),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_980),
.B(n_67),
.Y(n_1202)
);

NOR2x1_ASAP7_75t_L g1203 ( 
.A(n_961),
.B(n_67),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_925),
.A2(n_72),
.B(n_1016),
.Y(n_1204)
);

CKINVDCx16_ASAP7_75t_R g1205 ( 
.A(n_1048),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_919),
.A2(n_72),
.B(n_987),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_972),
.Y(n_1207)
);

AOI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1013),
.A2(n_1001),
.B(n_991),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1023),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1037),
.B(n_961),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1037),
.B(n_963),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_928),
.B(n_964),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1066),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_963),
.B(n_987),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_911),
.A2(n_893),
.B(n_933),
.C(n_947),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_966),
.B(n_1032),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_964),
.B(n_985),
.Y(n_1217)
);

AND2x4_ASAP7_75t_SL g1218 ( 
.A(n_1019),
.B(n_911),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_986),
.A2(n_995),
.B(n_937),
.C(n_996),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_992),
.A2(n_1018),
.B(n_1000),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1068),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_991),
.A2(n_1001),
.B1(n_1008),
.B2(n_1003),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1038),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1003),
.B(n_1008),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1009),
.A2(n_1017),
.B(n_968),
.Y(n_1225)
);

INVxp67_ASAP7_75t_L g1226 ( 
.A(n_1020),
.Y(n_1226)
);

AOI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1057),
.A2(n_1062),
.B(n_1073),
.Y(n_1227)
);

AO22x1_ASAP7_75t_L g1228 ( 
.A1(n_977),
.A2(n_999),
.B1(n_1071),
.B2(n_1070),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_954),
.B(n_1073),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1153),
.B(n_1020),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1124),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_SL g1232 ( 
.A1(n_1095),
.A2(n_1036),
.B(n_1028),
.C(n_1025),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1091),
.Y(n_1233)
);

NAND3xp33_ASAP7_75t_L g1234 ( 
.A(n_1092),
.B(n_1054),
.C(n_1065),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1092),
.A2(n_1063),
.B(n_1058),
.C(n_1029),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1166),
.A2(n_936),
.B(n_938),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1075),
.Y(n_1237)
);

INVxp67_ASAP7_75t_SL g1238 ( 
.A(n_1102),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1084),
.B(n_1036),
.Y(n_1239)
);

OA21x2_ASAP7_75t_L g1240 ( 
.A1(n_1206),
.A2(n_1067),
.B(n_1049),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_SL g1241 ( 
.A1(n_1077),
.A2(n_1045),
.B(n_1031),
.C(n_950),
.Y(n_1241)
);

INVx5_ASAP7_75t_L g1242 ( 
.A(n_1096),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1160),
.A2(n_943),
.B(n_948),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_1195),
.A2(n_967),
.A3(n_971),
.B(n_974),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1084),
.B(n_1099),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1225),
.A2(n_1167),
.A3(n_1219),
.B(n_1109),
.Y(n_1246)
);

NOR2xp67_ASAP7_75t_L g1247 ( 
.A(n_1078),
.B(n_1131),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1144),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1205),
.B(n_1093),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1088),
.A2(n_1157),
.B(n_1098),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1157),
.A2(n_1220),
.B(n_1108),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1103),
.B(n_1093),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1076),
.A2(n_1115),
.B(n_1228),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1192),
.B(n_1186),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1130),
.A2(n_1227),
.B(n_1208),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1186),
.A2(n_1136),
.B(n_1097),
.C(n_1113),
.Y(n_1256)
);

NAND3xp33_ASAP7_75t_L g1257 ( 
.A(n_1194),
.B(n_1113),
.C(n_1089),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1085),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1223),
.B(n_1136),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1094),
.A2(n_1215),
.B(n_1090),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1094),
.A2(n_1215),
.B(n_1090),
.Y(n_1261)
);

AO31x2_ASAP7_75t_L g1262 ( 
.A1(n_1222),
.A2(n_1181),
.A3(n_1187),
.B(n_1190),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1229),
.A2(n_1168),
.B(n_1216),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1079),
.B(n_1165),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1143),
.A2(n_1212),
.B(n_1105),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1210),
.A2(n_1204),
.A3(n_1135),
.B(n_1120),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1165),
.B(n_1148),
.Y(n_1267)
);

NOR2xp67_ASAP7_75t_L g1268 ( 
.A(n_1163),
.B(n_1112),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1116),
.A2(n_1118),
.B(n_1155),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1074),
.A2(n_1217),
.B(n_1080),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1169),
.B(n_1087),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1096),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1143),
.A2(n_1173),
.B(n_1214),
.Y(n_1273)
);

NAND2x1_ASAP7_75t_L g1274 ( 
.A(n_1200),
.B(n_1163),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1081),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1159),
.A2(n_1156),
.A3(n_1123),
.B(n_1172),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1173),
.A2(n_1080),
.B(n_1196),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1097),
.A2(n_1194),
.B(n_1089),
.C(n_1202),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1202),
.A2(n_1211),
.B(n_1129),
.C(n_1171),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1134),
.A2(n_1151),
.B(n_1193),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1142),
.A2(n_1221),
.B(n_1188),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1188),
.A2(n_1207),
.B(n_1218),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1179),
.A2(n_1201),
.A3(n_1164),
.B(n_1178),
.Y(n_1283)
);

AO21x1_ASAP7_75t_L g1284 ( 
.A1(n_1211),
.A2(n_1162),
.B(n_1224),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1137),
.A2(n_1213),
.B(n_1139),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1137),
.A2(n_1139),
.B(n_1150),
.Y(n_1286)
);

AOI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1209),
.A2(n_1086),
.B(n_1224),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1226),
.A2(n_1146),
.B(n_1154),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1081),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1114),
.B(n_1171),
.Y(n_1290)
);

INVx4_ASAP7_75t_L g1291 ( 
.A(n_1144),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1188),
.A2(n_1207),
.B(n_1209),
.Y(n_1292)
);

AOI31xp67_ASAP7_75t_L g1293 ( 
.A1(n_1147),
.A2(n_1152),
.A3(n_1158),
.B(n_1184),
.Y(n_1293)
);

O2A1O1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1191),
.A2(n_1162),
.B(n_1141),
.C(n_1199),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1096),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1144),
.Y(n_1296)
);

AO21x1_ASAP7_75t_L g1297 ( 
.A1(n_1185),
.A2(n_1145),
.B(n_1141),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1114),
.B(n_1106),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1087),
.B(n_1111),
.Y(n_1299)
);

INVx8_ASAP7_75t_L g1300 ( 
.A(n_1096),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1125),
.A2(n_1198),
.B1(n_1177),
.B2(n_1197),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1101),
.B(n_1180),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1226),
.A2(n_1188),
.B(n_1203),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1121),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1121),
.B(n_1126),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1083),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1207),
.A2(n_1149),
.B(n_1174),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1100),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1138),
.A2(n_1182),
.B(n_1183),
.C(n_1133),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1128),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1200),
.A2(n_1104),
.A3(n_1175),
.B(n_1207),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1180),
.B(n_1144),
.Y(n_1312)
);

AOI31xp67_ASAP7_75t_L g1313 ( 
.A1(n_1104),
.A2(n_1107),
.A3(n_1122),
.B(n_1119),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1104),
.A2(n_1176),
.B(n_1180),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1104),
.A2(n_1176),
.B(n_1180),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1180),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1180),
.Y(n_1317)
);

AOI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1189),
.A2(n_1161),
.B(n_1170),
.Y(n_1318)
);

AOI221xp5_ASAP7_75t_L g1319 ( 
.A1(n_1140),
.A2(n_1161),
.B1(n_1110),
.B2(n_1117),
.C(n_1127),
.Y(n_1319)
);

BUFx10_ASAP7_75t_L g1320 ( 
.A(n_1132),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1085),
.A2(n_1189),
.B(n_1082),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1092),
.A2(n_723),
.B(n_721),
.C(n_1093),
.Y(n_1322)
);

AND2x6_ASAP7_75t_L g1323 ( 
.A(n_1211),
.B(n_1096),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1084),
.B(n_723),
.Y(n_1324)
);

AOI221xp5_ASAP7_75t_L g1325 ( 
.A1(n_1153),
.A2(n_721),
.B1(n_1014),
.B2(n_723),
.C(n_1006),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_SL g1326 ( 
.A1(n_1095),
.A2(n_1077),
.B(n_735),
.C(n_1210),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1130),
.A2(n_1220),
.B(n_1109),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1130),
.A2(n_1220),
.B(n_1109),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_1124),
.Y(n_1329)
);

O2A1O1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1092),
.A2(n_721),
.B(n_723),
.C(n_728),
.Y(n_1330)
);

AO31x2_ASAP7_75t_L g1331 ( 
.A1(n_1195),
.A2(n_916),
.A3(n_940),
.B(n_1225),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1091),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1166),
.A2(n_723),
.B(n_610),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1153),
.B(n_721),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1195),
.A2(n_916),
.A3(n_940),
.B(n_1225),
.Y(n_1335)
);

O2A1O1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1092),
.A2(n_721),
.B(n_723),
.C(n_728),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1130),
.A2(n_1220),
.B(n_1109),
.Y(n_1337)
);

AOI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1228),
.A2(n_1225),
.B(n_1206),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1099),
.B(n_1153),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1099),
.B(n_1153),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1130),
.A2(n_1220),
.B(n_1109),
.Y(n_1341)
);

AO31x2_ASAP7_75t_L g1342 ( 
.A1(n_1195),
.A2(n_916),
.A3(n_940),
.B(n_1225),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1166),
.A2(n_723),
.B(n_610),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1130),
.A2(n_1220),
.B(n_1109),
.Y(n_1344)
);

AO31x2_ASAP7_75t_L g1345 ( 
.A1(n_1195),
.A2(n_916),
.A3(n_940),
.B(n_1225),
.Y(n_1345)
);

INVx5_ASAP7_75t_L g1346 ( 
.A(n_1096),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1153),
.B(n_721),
.Y(n_1347)
);

INVxp67_ASAP7_75t_SL g1348 ( 
.A(n_1102),
.Y(n_1348)
);

AOI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1153),
.A2(n_723),
.B1(n_721),
.B2(n_1092),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1124),
.Y(n_1350)
);

AOI21x1_ASAP7_75t_SL g1351 ( 
.A1(n_1185),
.A2(n_1199),
.B(n_1192),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1153),
.A2(n_723),
.B1(n_721),
.B2(n_1092),
.Y(n_1352)
);

O2A1O1Ixp5_ASAP7_75t_SL g1353 ( 
.A1(n_1129),
.A2(n_493),
.B(n_810),
.C(n_827),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1163),
.B(n_1169),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_SL g1355 ( 
.A1(n_1095),
.A2(n_1077),
.B(n_735),
.C(n_1210),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1130),
.A2(n_1220),
.B(n_1109),
.Y(n_1356)
);

AO31x2_ASAP7_75t_L g1357 ( 
.A1(n_1195),
.A2(n_916),
.A3(n_940),
.B(n_1225),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_SL g1358 ( 
.A(n_1124),
.B(n_835),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1075),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1092),
.A2(n_723),
.B(n_721),
.C(n_1093),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1091),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1166),
.A2(n_723),
.B(n_610),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1099),
.B(n_782),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1075),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1169),
.B(n_1007),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1153),
.B(n_721),
.Y(n_1366)
);

AO31x2_ASAP7_75t_L g1367 ( 
.A1(n_1195),
.A2(n_916),
.A3(n_940),
.B(n_1225),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1206),
.A2(n_1088),
.B(n_1166),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1166),
.A2(n_723),
.B(n_610),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1153),
.B(n_721),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1153),
.B(n_721),
.Y(n_1371)
);

O2A1O1Ixp5_ASAP7_75t_L g1372 ( 
.A1(n_1092),
.A2(n_723),
.B(n_721),
.C(n_728),
.Y(n_1372)
);

AOI221xp5_ASAP7_75t_L g1373 ( 
.A1(n_1153),
.A2(n_721),
.B1(n_1014),
.B2(n_723),
.C(n_1006),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1099),
.B(n_1153),
.Y(n_1374)
);

AO32x2_ASAP7_75t_L g1375 ( 
.A1(n_1125),
.A2(n_1179),
.A3(n_1076),
.B1(n_1222),
.B2(n_1156),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1166),
.A2(n_723),
.B(n_610),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1153),
.B(n_721),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1130),
.A2(n_1220),
.B(n_1109),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1153),
.B(n_721),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1166),
.A2(n_723),
.B(n_610),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1130),
.A2(n_1220),
.B(n_1109),
.Y(n_1381)
);

A2O1A1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1092),
.A2(n_723),
.B(n_721),
.C(n_1093),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1153),
.B(n_721),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_1110),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1075),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1092),
.A2(n_723),
.B1(n_721),
.B2(n_728),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1166),
.A2(n_723),
.B(n_610),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1166),
.A2(n_723),
.B(n_610),
.Y(n_1388)
);

NAND3xp33_ASAP7_75t_L g1389 ( 
.A(n_1092),
.B(n_721),
.C(n_723),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1092),
.A2(n_723),
.B1(n_721),
.B2(n_728),
.Y(n_1390)
);

BUFx4f_ASAP7_75t_SL g1391 ( 
.A(n_1329),
.Y(n_1391)
);

BUFx4_ASAP7_75t_SL g1392 ( 
.A(n_1231),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1386),
.A2(n_1390),
.B1(n_1249),
.B2(n_1257),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1257),
.A2(n_1389),
.B1(n_1325),
.B2(n_1373),
.Y(n_1394)
);

BUFx10_ASAP7_75t_L g1395 ( 
.A(n_1350),
.Y(n_1395)
);

CKINVDCx14_ASAP7_75t_R g1396 ( 
.A(n_1332),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1384),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1364),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1389),
.A2(n_1349),
.B1(n_1352),
.B2(n_1324),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1349),
.A2(n_1352),
.B1(n_1383),
.B2(n_1301),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1245),
.A2(n_1290),
.B1(n_1254),
.B2(n_1252),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1301),
.A2(n_1366),
.B1(n_1347),
.B2(n_1370),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1334),
.A2(n_1371),
.B1(n_1379),
.B2(n_1377),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1242),
.Y(n_1404)
);

OAI21xp33_ASAP7_75t_L g1405 ( 
.A1(n_1322),
.A2(n_1382),
.B(n_1360),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1233),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1297),
.A2(n_1284),
.B1(n_1340),
.B2(n_1339),
.Y(n_1407)
);

BUFx4f_ASAP7_75t_SL g1408 ( 
.A(n_1258),
.Y(n_1408)
);

BUFx12f_ASAP7_75t_L g1409 ( 
.A(n_1320),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1374),
.A2(n_1265),
.B1(n_1259),
.B2(n_1239),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1247),
.A2(n_1314),
.B1(n_1315),
.B2(n_1273),
.Y(n_1411)
);

INVx6_ASAP7_75t_L g1412 ( 
.A(n_1320),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1278),
.A2(n_1264),
.B1(n_1330),
.B2(n_1336),
.Y(n_1413)
);

CKINVDCx11_ASAP7_75t_R g1414 ( 
.A(n_1361),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1288),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1359),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1247),
.A2(n_1319),
.B1(n_1253),
.B2(n_1260),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1363),
.A2(n_1230),
.B1(n_1304),
.B2(n_1385),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1267),
.A2(n_1299),
.B1(n_1298),
.B2(n_1303),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1268),
.A2(n_1303),
.B1(n_1277),
.B2(n_1299),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1256),
.A2(n_1279),
.B1(n_1268),
.B2(n_1238),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_1348),
.Y(n_1422)
);

CKINVDCx11_ASAP7_75t_R g1423 ( 
.A(n_1271),
.Y(n_1423)
);

OAI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1304),
.A2(n_1289),
.B1(n_1275),
.B2(n_1261),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1242),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1271),
.A2(n_1358),
.B1(n_1305),
.B2(n_1323),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1270),
.A2(n_1372),
.B1(n_1250),
.B2(n_1368),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1270),
.A2(n_1368),
.B1(n_1263),
.B2(n_1310),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1287),
.Y(n_1429)
);

CKINVDCx10_ASAP7_75t_R g1430 ( 
.A(n_1318),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1306),
.B(n_1308),
.Y(n_1431)
);

BUFx4f_ASAP7_75t_L g1432 ( 
.A(n_1365),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1365),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1321),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_SL g1435 ( 
.A(n_1248),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1294),
.B(n_1302),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1309),
.A2(n_1282),
.B1(n_1354),
.B2(n_1292),
.Y(n_1437)
);

CKINVDCx6p67_ASAP7_75t_R g1438 ( 
.A(n_1346),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1248),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1326),
.B(n_1355),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1296),
.Y(n_1441)
);

INVx6_ASAP7_75t_L g1442 ( 
.A(n_1291),
.Y(n_1442)
);

BUFx8_ASAP7_75t_L g1443 ( 
.A(n_1296),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1293),
.Y(n_1444)
);

INVx6_ASAP7_75t_L g1445 ( 
.A(n_1291),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_SL g1446 ( 
.A1(n_1323),
.A2(n_1375),
.B1(n_1343),
.B2(n_1387),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1300),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1323),
.A2(n_1234),
.B1(n_1362),
.B2(n_1380),
.Y(n_1448)
);

BUFx2_ASAP7_75t_SL g1449 ( 
.A(n_1272),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1323),
.A2(n_1234),
.B1(n_1369),
.B2(n_1333),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1376),
.A2(n_1388),
.B1(n_1375),
.B2(n_1251),
.Y(n_1451)
);

BUFx10_ASAP7_75t_L g1452 ( 
.A(n_1316),
.Y(n_1452)
);

INVx6_ASAP7_75t_L g1453 ( 
.A(n_1300),
.Y(n_1453)
);

INVx4_ASAP7_75t_L g1454 ( 
.A(n_1295),
.Y(n_1454)
);

CKINVDCx11_ASAP7_75t_R g1455 ( 
.A(n_1317),
.Y(n_1455)
);

CKINVDCx11_ASAP7_75t_R g1456 ( 
.A(n_1351),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1375),
.A2(n_1280),
.B1(n_1307),
.B2(n_1312),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_SL g1458 ( 
.A1(n_1353),
.A2(n_1286),
.B1(n_1281),
.B2(n_1285),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1240),
.A2(n_1243),
.B1(n_1236),
.B2(n_1378),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1313),
.Y(n_1460)
);

INVx6_ASAP7_75t_L g1461 ( 
.A(n_1274),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1283),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1262),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1235),
.A2(n_1338),
.B(n_1232),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1240),
.A2(n_1328),
.B1(n_1356),
.B2(n_1344),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1283),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1311),
.Y(n_1467)
);

CKINVDCx14_ASAP7_75t_R g1468 ( 
.A(n_1241),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1262),
.A2(n_1276),
.B1(n_1266),
.B2(n_1311),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1327),
.A2(n_1381),
.B1(n_1341),
.B2(n_1337),
.Y(n_1470)
);

CKINVDCx11_ASAP7_75t_R g1471 ( 
.A(n_1266),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1262),
.A2(n_1311),
.B1(n_1276),
.B2(n_1266),
.Y(n_1472)
);

INVx6_ASAP7_75t_L g1473 ( 
.A(n_1244),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_1331),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1331),
.Y(n_1475)
);

OAI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1255),
.A2(n_1269),
.B(n_1276),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1246),
.A2(n_1335),
.B1(n_1342),
.B2(n_1345),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1335),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1246),
.A2(n_1342),
.B1(n_1345),
.B2(n_1357),
.Y(n_1479)
);

OAI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1246),
.A2(n_1342),
.B1(n_1345),
.B2(n_1357),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1367),
.A2(n_1257),
.B1(n_723),
.B2(n_1386),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1244),
.Y(n_1482)
);

BUFx12f_ASAP7_75t_L g1483 ( 
.A(n_1244),
.Y(n_1483)
);

OAI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1367),
.A2(n_1352),
.B1(n_1349),
.B2(n_1386),
.Y(n_1484)
);

INVx2_ASAP7_75t_SL g1485 ( 
.A(n_1320),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1248),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1389),
.A2(n_721),
.B1(n_723),
.B2(n_1386),
.Y(n_1487)
);

CKINVDCx8_ASAP7_75t_R g1488 ( 
.A(n_1384),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1386),
.A2(n_723),
.B1(n_721),
.B2(n_1390),
.Y(n_1489)
);

CKINVDCx11_ASAP7_75t_R g1490 ( 
.A(n_1329),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1329),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1257),
.A2(n_723),
.B1(n_1390),
.B2(n_1386),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1257),
.A2(n_723),
.B1(n_1390),
.B2(n_1386),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1237),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1257),
.A2(n_723),
.B1(n_1390),
.B2(n_1386),
.Y(n_1495)
);

CKINVDCx11_ASAP7_75t_R g1496 ( 
.A(n_1329),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1389),
.A2(n_721),
.B1(n_723),
.B2(n_1386),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1237),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1389),
.A2(n_721),
.B1(n_723),
.B2(n_1386),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1339),
.B(n_1340),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1242),
.Y(n_1501)
);

OAI21xp33_ASAP7_75t_L g1502 ( 
.A1(n_1325),
.A2(n_721),
.B(n_723),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1237),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1237),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1257),
.A2(n_723),
.B1(n_1390),
.B2(n_1386),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1242),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1242),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1237),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1389),
.A2(n_721),
.B1(n_723),
.B2(n_1386),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1233),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1332),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1242),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1333),
.A2(n_723),
.B(n_1387),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1332),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_SL g1515 ( 
.A1(n_1386),
.A2(n_723),
.B1(n_721),
.B2(n_1390),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_SL g1516 ( 
.A1(n_1386),
.A2(n_723),
.B1(n_721),
.B2(n_1390),
.Y(n_1516)
);

INVx5_ASAP7_75t_L g1517 ( 
.A(n_1300),
.Y(n_1517)
);

CKINVDCx11_ASAP7_75t_R g1518 ( 
.A(n_1329),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1257),
.A2(n_723),
.B1(n_1390),
.B2(n_1386),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1389),
.A2(n_721),
.B1(n_723),
.B2(n_1386),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1257),
.A2(n_723),
.B1(n_1390),
.B2(n_1386),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1231),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1392),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1403),
.B(n_1402),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1476),
.A2(n_1464),
.B(n_1470),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_SL g1526 ( 
.A(n_1488),
.Y(n_1526)
);

NOR2xp67_ASAP7_75t_R g1527 ( 
.A(n_1409),
.B(n_1412),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1415),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1415),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1463),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1481),
.B(n_1462),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1470),
.A2(n_1465),
.B(n_1459),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1483),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1475),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1481),
.B(n_1466),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1465),
.A2(n_1459),
.B(n_1513),
.Y(n_1536)
);

AOI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1444),
.A2(n_1437),
.B(n_1429),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1478),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1472),
.B(n_1429),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1502),
.A2(n_1489),
.B1(n_1515),
.B2(n_1516),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1460),
.Y(n_1541)
);

CKINVDCx8_ASAP7_75t_R g1542 ( 
.A(n_1430),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1403),
.B(n_1402),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1416),
.Y(n_1544)
);

INVxp67_ASAP7_75t_SL g1545 ( 
.A(n_1422),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1479),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1473),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1487),
.A2(n_1497),
.B(n_1509),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1467),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1473),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1474),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1412),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1482),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1392),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1482),
.Y(n_1555)
);

AOI22x1_ASAP7_75t_L g1556 ( 
.A1(n_1499),
.A2(n_1520),
.B1(n_1495),
.B2(n_1492),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1448),
.A2(n_1450),
.B(n_1451),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1500),
.B(n_1391),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1401),
.B(n_1394),
.Y(n_1559)
);

INVxp67_ASAP7_75t_SL g1560 ( 
.A(n_1436),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1480),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1480),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1511),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1448),
.A2(n_1450),
.B(n_1451),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1471),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1469),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1469),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1477),
.Y(n_1568)
);

CKINVDCx12_ASAP7_75t_R g1569 ( 
.A(n_1391),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1477),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1440),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1443),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1456),
.Y(n_1573)
);

NAND2x1p5_ASAP7_75t_L g1574 ( 
.A(n_1517),
.B(n_1404),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1398),
.Y(n_1575)
);

OAI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1427),
.A2(n_1428),
.B(n_1411),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1494),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1427),
.A2(n_1428),
.B(n_1411),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1410),
.B(n_1484),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1399),
.B(n_1413),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1498),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1503),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1504),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1399),
.B(n_1410),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1394),
.B(n_1393),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1508),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1424),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1492),
.A2(n_1505),
.B1(n_1493),
.B2(n_1521),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1443),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1407),
.B(n_1400),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1484),
.B(n_1407),
.Y(n_1591)
);

AO21x2_ASAP7_75t_L g1592 ( 
.A1(n_1424),
.A2(n_1421),
.B(n_1405),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1420),
.B(n_1457),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1514),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1452),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1457),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1468),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1418),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1490),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1431),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1418),
.B(n_1400),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1426),
.B(n_1417),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_SL g1603 ( 
.A1(n_1425),
.A2(n_1506),
.B(n_1501),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1446),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1458),
.Y(n_1605)
);

OAI21x1_ASAP7_75t_L g1606 ( 
.A1(n_1417),
.A2(n_1493),
.B(n_1505),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1461),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1495),
.A2(n_1521),
.B1(n_1519),
.B2(n_1419),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1519),
.Y(n_1609)
);

NOR2x1_ASAP7_75t_SL g1610 ( 
.A(n_1425),
.B(n_1506),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1461),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1486),
.B(n_1441),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1461),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1449),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1454),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1439),
.A2(n_1433),
.B(n_1485),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1406),
.B(n_1510),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1432),
.B(n_1455),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1506),
.Y(n_1619)
);

OA21x2_ASAP7_75t_L g1620 ( 
.A1(n_1397),
.A2(n_1435),
.B(n_1404),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1434),
.A2(n_1414),
.B1(n_1423),
.B2(n_1396),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1551),
.B(n_1395),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1536),
.A2(n_1435),
.B(n_1438),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1585),
.B(n_1560),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1551),
.B(n_1395),
.Y(n_1625)
);

O2A1O1Ixp33_ASAP7_75t_SL g1626 ( 
.A1(n_1588),
.A2(n_1512),
.B(n_1507),
.C(n_1517),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1548),
.B(n_1442),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1523),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_SL g1629 ( 
.A(n_1542),
.B(n_1408),
.Y(n_1629)
);

A2O1A1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_1540),
.A2(n_1507),
.B(n_1512),
.C(n_1517),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1556),
.A2(n_1580),
.B1(n_1608),
.B2(n_1584),
.Y(n_1631)
);

OAI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1556),
.A2(n_1491),
.B(n_1517),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1559),
.B(n_1442),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1601),
.A2(n_1573),
.B1(n_1597),
.B2(n_1524),
.Y(n_1634)
);

OA21x2_ASAP7_75t_L g1635 ( 
.A1(n_1525),
.A2(n_1512),
.B(n_1445),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1528),
.Y(n_1636)
);

BUFx4f_ASAP7_75t_SL g1637 ( 
.A(n_1572),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1565),
.B(n_1447),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1606),
.A2(n_1522),
.B(n_1408),
.Y(n_1639)
);

O2A1O1Ixp33_ASAP7_75t_SL g1640 ( 
.A1(n_1543),
.A2(n_1453),
.B(n_1496),
.C(n_1518),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1565),
.B(n_1453),
.Y(n_1641)
);

OAI21x1_ASAP7_75t_L g1642 ( 
.A1(n_1536),
.A2(n_1532),
.B(n_1537),
.Y(n_1642)
);

AOI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1609),
.A2(n_1584),
.B1(n_1590),
.B2(n_1587),
.C(n_1604),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1600),
.B(n_1612),
.Y(n_1644)
);

CKINVDCx20_ASAP7_75t_R g1645 ( 
.A(n_1599),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1533),
.B(n_1547),
.Y(n_1646)
);

A2O1A1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1602),
.A2(n_1579),
.B(n_1590),
.C(n_1601),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1546),
.B(n_1545),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1533),
.B(n_1547),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1602),
.A2(n_1592),
.B1(n_1609),
.B2(n_1573),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1579),
.A2(n_1602),
.B(n_1564),
.Y(n_1651)
);

NAND2xp33_ASAP7_75t_L g1652 ( 
.A(n_1573),
.B(n_1618),
.Y(n_1652)
);

A2O1A1Ixp33_ASAP7_75t_L g1653 ( 
.A1(n_1602),
.A2(n_1591),
.B(n_1587),
.C(n_1593),
.Y(n_1653)
);

AOI221xp5_ASAP7_75t_L g1654 ( 
.A1(n_1546),
.A2(n_1592),
.B1(n_1598),
.B2(n_1605),
.C(n_1593),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1554),
.Y(n_1655)
);

INVx5_ASAP7_75t_SL g1656 ( 
.A(n_1573),
.Y(n_1656)
);

NAND2x1p5_ASAP7_75t_L g1657 ( 
.A(n_1616),
.B(n_1620),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1529),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1531),
.B(n_1535),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1592),
.B(n_1598),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1544),
.B(n_1575),
.Y(n_1661)
);

OR2x6_ASAP7_75t_L g1662 ( 
.A(n_1533),
.B(n_1557),
.Y(n_1662)
);

OAI21xp33_ASAP7_75t_SL g1663 ( 
.A1(n_1603),
.A2(n_1591),
.B(n_1614),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1535),
.B(n_1616),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1573),
.A2(n_1558),
.B1(n_1593),
.B2(n_1618),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1557),
.A2(n_1564),
.B(n_1578),
.Y(n_1666)
);

AO32x2_ASAP7_75t_L g1667 ( 
.A1(n_1539),
.A2(n_1561),
.A3(n_1562),
.B1(n_1567),
.B2(n_1566),
.Y(n_1667)
);

NAND3xp33_ASAP7_75t_L g1668 ( 
.A(n_1573),
.B(n_1563),
.C(n_1614),
.Y(n_1668)
);

AO21x2_ASAP7_75t_L g1669 ( 
.A1(n_1537),
.A2(n_1532),
.B(n_1525),
.Y(n_1669)
);

AOI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1593),
.A2(n_1596),
.B1(n_1562),
.B2(n_1561),
.C(n_1594),
.Y(n_1670)
);

OA21x2_ASAP7_75t_L g1671 ( 
.A1(n_1576),
.A2(n_1578),
.B(n_1541),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1603),
.A2(n_1610),
.B(n_1616),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1575),
.B(n_1581),
.Y(n_1673)
);

AO32x2_ASAP7_75t_L g1674 ( 
.A1(n_1539),
.A2(n_1596),
.A3(n_1570),
.B1(n_1568),
.B2(n_1549),
.Y(n_1674)
);

OA21x2_ASAP7_75t_L g1675 ( 
.A1(n_1534),
.A2(n_1538),
.B(n_1530),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1581),
.B(n_1582),
.Y(n_1676)
);

AO21x1_ASAP7_75t_L g1677 ( 
.A1(n_1615),
.A2(n_1549),
.B(n_1586),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1582),
.B(n_1583),
.Y(n_1678)
);

A2O1A1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1597),
.A2(n_1568),
.B(n_1570),
.C(n_1571),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1675),
.Y(n_1680)
);

BUFx3_ASAP7_75t_L g1681 ( 
.A(n_1657),
.Y(n_1681)
);

OAI221xp5_ASAP7_75t_L g1682 ( 
.A1(n_1631),
.A2(n_1542),
.B1(n_1621),
.B2(n_1617),
.C(n_1552),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1675),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1631),
.A2(n_1611),
.B1(n_1607),
.B2(n_1613),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1624),
.B(n_1583),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1636),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1664),
.B(n_1530),
.Y(n_1687)
);

NOR2xp67_ASAP7_75t_L g1688 ( 
.A(n_1672),
.B(n_1595),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1659),
.B(n_1553),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1644),
.B(n_1538),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1653),
.A2(n_1526),
.B1(n_1571),
.B2(n_1572),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1636),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1658),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1633),
.B(n_1617),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1653),
.A2(n_1571),
.B1(n_1572),
.B2(n_1589),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1645),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1635),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1673),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1674),
.B(n_1555),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1676),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1674),
.B(n_1667),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1660),
.B(n_1650),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1660),
.B(n_1577),
.Y(n_1703)
);

AND2x2_ASAP7_75t_SL g1704 ( 
.A(n_1652),
.B(n_1620),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1674),
.B(n_1555),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1633),
.B(n_1569),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1678),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1622),
.B(n_1569),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1677),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1662),
.B(n_1550),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1661),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1639),
.B(n_1552),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1699),
.B(n_1666),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1699),
.B(n_1662),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1683),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1683),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1680),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1705),
.B(n_1662),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1705),
.B(n_1671),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1696),
.Y(n_1720)
);

OAI21xp33_ASAP7_75t_L g1721 ( 
.A1(n_1702),
.A2(n_1647),
.B(n_1643),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1697),
.B(n_1710),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1697),
.B(n_1623),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1701),
.B(n_1671),
.Y(n_1724)
);

INVx4_ASAP7_75t_L g1725 ( 
.A(n_1704),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1697),
.B(n_1623),
.Y(n_1726)
);

AO21x2_ASAP7_75t_L g1727 ( 
.A1(n_1709),
.A2(n_1642),
.B(n_1669),
.Y(n_1727)
);

INVxp67_ASAP7_75t_L g1728 ( 
.A(n_1709),
.Y(n_1728)
);

OAI31xp33_ASAP7_75t_L g1729 ( 
.A1(n_1691),
.A2(n_1682),
.A3(n_1647),
.B(n_1695),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1684),
.A2(n_1630),
.B1(n_1654),
.B2(n_1679),
.Y(n_1730)
);

NAND3xp33_ASAP7_75t_L g1731 ( 
.A(n_1691),
.B(n_1670),
.C(n_1679),
.Y(n_1731)
);

NOR2x1_ASAP7_75t_L g1732 ( 
.A(n_1688),
.B(n_1668),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1695),
.A2(n_1630),
.B1(n_1634),
.B2(n_1651),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_1686),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1703),
.B(n_1711),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1700),
.B(n_1667),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1687),
.B(n_1648),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1700),
.B(n_1667),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1697),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1697),
.B(n_1667),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1698),
.B(n_1646),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1698),
.B(n_1649),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1728),
.B(n_1685),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1728),
.B(n_1707),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1719),
.B(n_1681),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1740),
.B(n_1692),
.Y(n_1746)
);

INVx1_ASAP7_75t_SL g1747 ( 
.A(n_1734),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1715),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1715),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1719),
.B(n_1704),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1735),
.B(n_1707),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1717),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1719),
.B(n_1704),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1740),
.B(n_1710),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1717),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1725),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1735),
.B(n_1690),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1722),
.B(n_1710),
.Y(n_1758)
);

BUFx2_ASAP7_75t_L g1759 ( 
.A(n_1725),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1724),
.B(n_1710),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1724),
.B(n_1689),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1736),
.B(n_1690),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1716),
.Y(n_1763)
);

INVx3_ASAP7_75t_L g1764 ( 
.A(n_1722),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1736),
.B(n_1693),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1716),
.Y(n_1766)
);

BUFx2_ASAP7_75t_L g1767 ( 
.A(n_1725),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1736),
.B(n_1693),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1716),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1738),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1762),
.B(n_1734),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1750),
.B(n_1713),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1750),
.B(n_1713),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1748),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1750),
.B(n_1713),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1747),
.B(n_1721),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1762),
.B(n_1737),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1756),
.B(n_1725),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1748),
.Y(n_1779)
);

NAND2xp33_ASAP7_75t_L g1780 ( 
.A(n_1747),
.B(n_1721),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1750),
.B(n_1725),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1757),
.B(n_1741),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1757),
.B(n_1741),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1746),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1753),
.B(n_1725),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1746),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1743),
.B(n_1741),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1753),
.B(n_1756),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1748),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1749),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1749),
.Y(n_1791)
);

INVxp67_ASAP7_75t_L g1792 ( 
.A(n_1743),
.Y(n_1792)
);

NAND2x1_ASAP7_75t_L g1793 ( 
.A(n_1756),
.B(n_1732),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1759),
.B(n_1723),
.Y(n_1794)
);

NAND2x1p5_ASAP7_75t_L g1795 ( 
.A(n_1759),
.B(n_1732),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1749),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1763),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1763),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1763),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1765),
.B(n_1737),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1751),
.B(n_1720),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1753),
.B(n_1714),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1766),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1766),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1751),
.B(n_1742),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1758),
.B(n_1720),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1746),
.Y(n_1807)
);

NOR2xp67_ASAP7_75t_L g1808 ( 
.A(n_1764),
.B(n_1714),
.Y(n_1808)
);

OAI31xp33_ASAP7_75t_L g1809 ( 
.A1(n_1759),
.A2(n_1731),
.A3(n_1729),
.B(n_1733),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1766),
.Y(n_1810)
);

INVxp67_ASAP7_75t_L g1811 ( 
.A(n_1744),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1744),
.B(n_1742),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1753),
.B(n_1742),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1767),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1769),
.Y(n_1815)
);

NOR3xp33_ASAP7_75t_L g1816 ( 
.A(n_1780),
.B(n_1731),
.C(n_1733),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1779),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1809),
.B(n_1694),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1788),
.B(n_1754),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1788),
.B(n_1754),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1771),
.B(n_1765),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1795),
.Y(n_1822)
);

NOR3xp33_ASAP7_75t_SL g1823 ( 
.A(n_1776),
.B(n_1655),
.C(n_1628),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1802),
.B(n_1754),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1779),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1797),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1780),
.B(n_1754),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1771),
.B(n_1768),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1792),
.B(n_1714),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1801),
.B(n_1811),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1787),
.B(n_1768),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1802),
.B(n_1772),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1777),
.B(n_1746),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1814),
.B(n_1718),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1772),
.B(n_1767),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1773),
.B(n_1767),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1806),
.B(n_1718),
.Y(n_1837)
);

NOR3xp33_ASAP7_75t_L g1838 ( 
.A(n_1793),
.B(n_1730),
.C(n_1632),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1777),
.B(n_1800),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1797),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1798),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1773),
.B(n_1758),
.Y(n_1842)
);

INVxp67_ASAP7_75t_SL g1843 ( 
.A(n_1793),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_L g1844 ( 
.A(n_1812),
.B(n_1645),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1798),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1782),
.B(n_1628),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1810),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1810),
.Y(n_1848)
);

BUFx2_ASAP7_75t_SL g1849 ( 
.A(n_1778),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1775),
.B(n_1758),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1784),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1815),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1817),
.Y(n_1853)
);

AOI21xp33_ASAP7_75t_L g1854 ( 
.A1(n_1830),
.A2(n_1795),
.B(n_1729),
.Y(n_1854)
);

OAI21xp33_ASAP7_75t_SL g1855 ( 
.A1(n_1843),
.A2(n_1818),
.B(n_1827),
.Y(n_1855)
);

AOI211xp5_ASAP7_75t_L g1856 ( 
.A1(n_1816),
.A2(n_1730),
.B(n_1640),
.C(n_1778),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1832),
.B(n_1775),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1838),
.A2(n_1795),
.B1(n_1808),
.B2(n_1813),
.Y(n_1858)
);

OAI21xp33_ASAP7_75t_L g1859 ( 
.A1(n_1832),
.A2(n_1785),
.B(n_1781),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1835),
.B(n_1836),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1817),
.Y(n_1861)
);

AOI222xp33_ASAP7_75t_L g1862 ( 
.A1(n_1844),
.A2(n_1778),
.B1(n_1781),
.B2(n_1785),
.C1(n_1712),
.C2(n_1794),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1823),
.B(n_1794),
.Y(n_1863)
);

NAND3xp33_ASAP7_75t_L g1864 ( 
.A(n_1822),
.B(n_1627),
.C(n_1774),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1835),
.B(n_1805),
.Y(n_1865)
);

OAI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1837),
.A2(n_1732),
.B1(n_1656),
.B2(n_1665),
.Y(n_1866)
);

INVxp67_ASAP7_75t_L g1867 ( 
.A(n_1849),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1836),
.B(n_1758),
.Y(n_1868)
);

NAND4xp25_ASAP7_75t_L g1869 ( 
.A(n_1846),
.B(n_1640),
.C(n_1629),
.D(n_1706),
.Y(n_1869)
);

AOI322xp5_ASAP7_75t_L g1870 ( 
.A1(n_1819),
.A2(n_1770),
.A3(n_1718),
.B1(n_1783),
.B2(n_1745),
.C1(n_1794),
.C2(n_1761),
.Y(n_1870)
);

INVxp67_ASAP7_75t_SL g1871 ( 
.A(n_1851),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_SL g1872 ( 
.A1(n_1819),
.A2(n_1625),
.B(n_1708),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1849),
.A2(n_1652),
.B1(n_1663),
.B2(n_1723),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1820),
.B(n_1800),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1822),
.Y(n_1875)
);

INVx1_ASAP7_75t_SL g1876 ( 
.A(n_1839),
.Y(n_1876)
);

OAI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1829),
.A2(n_1656),
.B1(n_1758),
.B2(n_1764),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1820),
.A2(n_1727),
.B1(n_1723),
.B2(n_1726),
.Y(n_1878)
);

INVxp67_ASAP7_75t_L g1879 ( 
.A(n_1871),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1876),
.B(n_1824),
.Y(n_1880)
);

A2O1A1Ixp33_ASAP7_75t_L g1881 ( 
.A1(n_1855),
.A2(n_1839),
.B(n_1834),
.C(n_1828),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1871),
.Y(n_1882)
);

AOI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1863),
.A2(n_1824),
.B1(n_1842),
.B2(n_1850),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1860),
.B(n_1842),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1867),
.B(n_1850),
.Y(n_1885)
);

OAI21xp33_ASAP7_75t_L g1886 ( 
.A1(n_1854),
.A2(n_1828),
.B(n_1821),
.Y(n_1886)
);

INVxp33_ASAP7_75t_L g1887 ( 
.A(n_1869),
.Y(n_1887)
);

A2O1A1Ixp33_ASAP7_75t_L g1888 ( 
.A1(n_1856),
.A2(n_1821),
.B(n_1833),
.C(n_1723),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_SL g1889 ( 
.A1(n_1858),
.A2(n_1637),
.B1(n_1833),
.B2(n_1770),
.Y(n_1889)
);

OAI21xp5_ASAP7_75t_SL g1890 ( 
.A1(n_1862),
.A2(n_1764),
.B(n_1831),
.Y(n_1890)
);

OAI21xp5_ASAP7_75t_SL g1891 ( 
.A1(n_1863),
.A2(n_1764),
.B(n_1831),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1853),
.Y(n_1892)
);

AOI21xp33_ASAP7_75t_SL g1893 ( 
.A1(n_1866),
.A2(n_1655),
.B(n_1851),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1859),
.A2(n_1726),
.B1(n_1723),
.B2(n_1764),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1864),
.A2(n_1851),
.B(n_1826),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1868),
.B(n_1758),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1861),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1857),
.Y(n_1898)
);

INVx1_ASAP7_75t_SL g1899 ( 
.A(n_1882),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1887),
.B(n_1872),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1898),
.B(n_1865),
.Y(n_1901)
);

INVxp67_ASAP7_75t_L g1902 ( 
.A(n_1885),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1884),
.B(n_1875),
.Y(n_1903)
);

INVxp67_ASAP7_75t_L g1904 ( 
.A(n_1880),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1879),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1881),
.B(n_1874),
.Y(n_1906)
);

INVx2_ASAP7_75t_SL g1907 ( 
.A(n_1896),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1879),
.B(n_1870),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1892),
.B(n_1873),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1883),
.B(n_1877),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1903),
.B(n_1889),
.Y(n_1911)
);

OAI32xp33_ASAP7_75t_L g1912 ( 
.A1(n_1908),
.A2(n_1886),
.A3(n_1895),
.B1(n_1897),
.B2(n_1878),
.Y(n_1912)
);

NOR2xp33_ASAP7_75t_L g1913 ( 
.A(n_1904),
.B(n_1891),
.Y(n_1913)
);

NOR3xp33_ASAP7_75t_L g1914 ( 
.A(n_1902),
.B(n_1893),
.C(n_1889),
.Y(n_1914)
);

NOR3xp33_ASAP7_75t_L g1915 ( 
.A(n_1900),
.B(n_1888),
.C(n_1890),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1907),
.Y(n_1916)
);

NOR3x1_ASAP7_75t_L g1917 ( 
.A(n_1908),
.B(n_1826),
.C(n_1825),
.Y(n_1917)
);

NOR2x1_ASAP7_75t_L g1918 ( 
.A(n_1905),
.B(n_1825),
.Y(n_1918)
);

OAI322xp33_ASAP7_75t_L g1919 ( 
.A1(n_1906),
.A2(n_1894),
.A3(n_1845),
.B1(n_1852),
.B2(n_1848),
.C1(n_1847),
.C2(n_1840),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1899),
.B(n_1784),
.Y(n_1920)
);

AOI322xp5_ASAP7_75t_L g1921 ( 
.A1(n_1915),
.A2(n_1901),
.A3(n_1899),
.B1(n_1909),
.B2(n_1910),
.C1(n_1878),
.C2(n_1852),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1920),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1911),
.B(n_1909),
.Y(n_1923)
);

AOI221xp5_ASAP7_75t_L g1924 ( 
.A1(n_1912),
.A2(n_1848),
.B1(n_1847),
.B2(n_1845),
.C(n_1841),
.Y(n_1924)
);

NOR2xp67_ASAP7_75t_L g1925 ( 
.A(n_1916),
.B(n_1840),
.Y(n_1925)
);

NOR2x1_ASAP7_75t_L g1926 ( 
.A(n_1923),
.B(n_1918),
.Y(n_1926)
);

NAND2x1p5_ASAP7_75t_L g1927 ( 
.A(n_1922),
.B(n_1925),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1924),
.Y(n_1928)
);

O2A1O1Ixp33_ASAP7_75t_SL g1929 ( 
.A1(n_1921),
.A2(n_1913),
.B(n_1917),
.C(n_1841),
.Y(n_1929)
);

AOI221xp5_ASAP7_75t_L g1930 ( 
.A1(n_1923),
.A2(n_1914),
.B1(n_1919),
.B2(n_1807),
.C(n_1786),
.Y(n_1930)
);

NAND4xp25_ASAP7_75t_L g1931 ( 
.A(n_1923),
.B(n_1589),
.C(n_1638),
.D(n_1641),
.Y(n_1931)
);

AND2x4_ASAP7_75t_L g1932 ( 
.A(n_1926),
.B(n_1786),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1930),
.B(n_1807),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1927),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1931),
.B(n_1637),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1928),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1932),
.Y(n_1937)
);

AOI322xp5_ASAP7_75t_L g1938 ( 
.A1(n_1936),
.A2(n_1929),
.A3(n_1764),
.B1(n_1745),
.B2(n_1815),
.C1(n_1799),
.C2(n_1796),
.Y(n_1938)
);

OAI32xp33_ASAP7_75t_L g1939 ( 
.A1(n_1934),
.A2(n_1589),
.A3(n_1803),
.B1(n_1791),
.B2(n_1790),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1937),
.Y(n_1940)
);

BUFx2_ASAP7_75t_L g1941 ( 
.A(n_1940),
.Y(n_1941)
);

AO22x2_ASAP7_75t_L g1942 ( 
.A1(n_1941),
.A2(n_1932),
.B1(n_1933),
.B2(n_1938),
.Y(n_1942)
);

NOR2xp67_ASAP7_75t_L g1943 ( 
.A(n_1941),
.B(n_1935),
.Y(n_1943)
);

OAI22x1_ASAP7_75t_L g1944 ( 
.A1(n_1942),
.A2(n_1939),
.B1(n_1804),
.B2(n_1789),
.Y(n_1944)
);

AND3x1_ASAP7_75t_L g1945 ( 
.A(n_1943),
.B(n_1527),
.C(n_1739),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1945),
.B(n_1760),
.Y(n_1946)
);

OAI22xp5_ASAP7_75t_SL g1947 ( 
.A1(n_1946),
.A2(n_1944),
.B1(n_1620),
.B2(n_1574),
.Y(n_1947)
);

AOI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1947),
.A2(n_1755),
.B(n_1752),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1948),
.Y(n_1949)
);

AOI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1949),
.A2(n_1739),
.B1(n_1726),
.B2(n_1723),
.Y(n_1950)
);

AOI211xp5_ASAP7_75t_L g1951 ( 
.A1(n_1950),
.A2(n_1626),
.B(n_1739),
.C(n_1619),
.Y(n_1951)
);


endmodule