module fake_jpeg_17905_n_39 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_39);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_17;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

AND2x2_ASAP7_75t_L g15 ( 
.A(n_14),
.B(n_1),
.Y(n_15)
);

INVxp67_ASAP7_75t_SL g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_5),
.A2(n_7),
.B1(n_1),
.B2(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_18),
.A2(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_25),
.B(n_30),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_9),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_15),
.B(n_2),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_27),
.B(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_3),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_15),
.A2(n_8),
.B1(n_20),
.B2(n_21),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_25),
.C(n_31),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_35),
.Y(n_37)
);

AOI322xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_33),
.A3(n_28),
.B1(n_16),
.B2(n_17),
.C1(n_27),
.C2(n_24),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_17),
.B(n_24),
.Y(n_39)
);


endmodule