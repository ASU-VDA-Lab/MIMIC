module fake_jpeg_209_n_265 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_0),
.B(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_39),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_42),
.B(n_55),
.Y(n_118)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_64),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_1),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_68),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_17),
.B(n_3),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_6),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_73),
.Y(n_95)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_72),
.Y(n_88)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_77),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_34),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_21),
.Y(n_104)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_76),
.A2(n_31),
.B1(n_35),
.B2(n_38),
.Y(n_94)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_79),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_81),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_13),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_23),
.B1(n_30),
.B2(n_40),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_99),
.B1(n_108),
.B2(n_117),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_46),
.A2(n_21),
.B1(n_33),
.B2(n_29),
.Y(n_99)
);

NAND2x1_ASAP7_75t_SL g154 ( 
.A(n_104),
.B(n_115),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_42),
.B(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_112),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_68),
.A2(n_18),
.B1(n_33),
.B2(n_29),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_30),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_41),
.B(n_38),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_122),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_50),
.A2(n_28),
.B1(n_24),
.B2(n_18),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_28),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_52),
.B(n_6),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_9),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_63),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_125)
);

OAI22x1_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_67),
.B1(n_9),
.B2(n_11),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_126),
.A2(n_127),
.B1(n_140),
.B2(n_148),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_99),
.A2(n_102),
.B1(n_83),
.B2(n_97),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_128),
.B(n_135),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_62),
.C(n_69),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_147),
.Y(n_164)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_131),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_95),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_136),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_91),
.B(n_8),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_146),
.Y(n_182)
);

BUFx8_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_94),
.A2(n_66),
.B1(n_78),
.B2(n_79),
.Y(n_140)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_11),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_98),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_154),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_88),
.B(n_58),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_86),
.A2(n_89),
.B1(n_87),
.B2(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_82),
.B(n_13),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_13),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_106),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_152),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_111),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_105),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_155),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_89),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_158),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

NOR2x1_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_100),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_84),
.B(n_116),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_114),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_161),
.Y(n_172)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_100),
.B(n_119),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_96),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_127),
.B(n_147),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_130),
.A2(n_110),
.B1(n_92),
.B2(n_119),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_183),
.B1(n_131),
.B2(n_153),
.Y(n_193)
);

NAND2xp33_ASAP7_75t_SL g179 ( 
.A(n_129),
.B(n_140),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_187),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_137),
.A2(n_92),
.B1(n_148),
.B2(n_126),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_141),
.B(n_145),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_144),
.B(n_150),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_194),
.Y(n_221)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_132),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_195),
.B(n_202),
.Y(n_219)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_139),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_206),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_144),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_164),
.C(n_175),
.Y(n_211)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_201),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_162),
.B1(n_143),
.B2(n_160),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_199),
.A2(n_200),
.B(n_179),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_172),
.A2(n_178),
.B1(n_181),
.B2(n_186),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_203),
.B(n_204),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_139),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_157),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_157),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_175),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_136),
.B1(n_170),
.B2(n_183),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_208),
.A2(n_199),
.B(n_205),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_213),
.C(n_218),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_192),
.C(n_191),
.Y(n_213)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_175),
.B(n_185),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_224),
.B(n_200),
.Y(n_227)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_209),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_187),
.C(n_180),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_222),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_177),
.C(n_165),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_205),
.A2(n_166),
.B(n_168),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_227),
.A2(n_215),
.B(n_224),
.Y(n_241)
);

AOI21xp33_ASAP7_75t_SL g228 ( 
.A1(n_213),
.A2(n_207),
.B(n_168),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_226),
.C(n_232),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_223),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_231),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_221),
.Y(n_230)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_190),
.B1(n_196),
.B2(n_201),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_182),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_190),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_243),
.Y(n_248)
);

A2O1A1O1Ixp25_ASAP7_75t_L g240 ( 
.A1(n_226),
.A2(n_211),
.B(n_220),
.C(n_222),
.D(n_218),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_241),
.B(n_238),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_232),
.C(n_225),
.Y(n_246)
);

OAI321xp33_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_177),
.A3(n_203),
.B1(n_176),
.B2(n_198),
.C(n_194),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_246),
.C(n_234),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_244),
.A2(n_234),
.B1(n_233),
.B2(n_230),
.Y(n_247)
);

AO21x1_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_227),
.B(n_174),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_231),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_249),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_225),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_241),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_253),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_254),
.A2(n_248),
.B1(n_247),
.B2(n_174),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_169),
.B(n_189),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_251),
.B(n_188),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_258),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_188),
.C(n_189),
.Y(n_258)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_256),
.B(n_166),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_260),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_258),
.C(n_165),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_263),
.B(n_259),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_262),
.Y(n_265)
);


endmodule