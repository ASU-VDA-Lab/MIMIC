module real_aes_13905_n_9 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_1, n_9);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_1;
output n_9;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_23;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_10;
OAI221xp5_ASAP7_75t_L g20 ( .A1(n_0), .A2(n_4), .B1(n_14), .B2(n_21), .C(n_25), .Y(n_20) );
INVx1_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
AOI321xp33_ASAP7_75t_L g9 ( .A1(n_2), .A2(n_8), .A3(n_10), .B1(n_13), .B2(n_15), .C(n_19), .Y(n_9) );
INVx1_ASAP7_75t_L g17 ( .A(n_3), .Y(n_17) );
INVx3_ASAP7_75t_L g24 ( .A(n_5), .Y(n_24) );
OAI21xp33_ASAP7_75t_L g15 ( .A1(n_6), .A2(n_16), .B(n_18), .Y(n_15) );
INVx1_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_10), .B(n_20), .Y(n_19) );
INVx1_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_11), .B(n_13), .Y(n_18) );
INVx1_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
INVx1_ASAP7_75t_L g13 ( .A(n_14), .Y(n_13) );
INVx1_ASAP7_75t_L g16 ( .A(n_17), .Y(n_16) );
BUFx3_ASAP7_75t_L g21 ( .A(n_22), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
INVx2_ASAP7_75t_L g23 ( .A(n_24), .Y(n_23) );
INVx1_ASAP7_75t_L g25 ( .A(n_26), .Y(n_25) );
endmodule