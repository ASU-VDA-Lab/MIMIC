module real_jpeg_430_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_1),
.A2(n_67),
.B1(n_68),
.B2(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_75),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_1),
.A2(n_34),
.B1(n_36),
.B2(n_75),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_2),
.A2(n_82),
.B1(n_83),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_2),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_2),
.A2(n_67),
.B1(n_68),
.B2(n_109),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_109),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_2),
.A2(n_34),
.B1(n_36),
.B2(n_109),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_4),
.A2(n_82),
.B1(n_83),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_4),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_4),
.A2(n_67),
.B1(n_68),
.B2(n_94),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_94),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_4),
.A2(n_34),
.B1(n_36),
.B2(n_94),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_5),
.A2(n_67),
.B(n_71),
.C(n_72),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_5),
.B(n_67),
.Y(n_71)
);

AO22x2_ASAP7_75t_L g72 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_73),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_5),
.A2(n_11),
.B(n_67),
.C(n_158),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_6),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_8),
.A2(n_34),
.B1(n_36),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_10),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_10),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_10),
.A2(n_67),
.B1(n_68),
.B2(n_81),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_81),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_10),
.A2(n_34),
.B1(n_36),
.B2(n_81),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_11),
.B(n_83),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_11),
.B(n_110),
.Y(n_146)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_11),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_11),
.B(n_72),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_11),
.A2(n_67),
.B1(n_68),
.B2(n_159),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_11),
.B(n_31),
.C(n_34),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_159),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_11),
.B(n_46),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_11),
.B(n_61),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_12),
.A2(n_34),
.B1(n_36),
.B2(n_41),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_13),
.A2(n_34),
.B1(n_36),
.B2(n_39),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_14),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_15),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_15),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_15),
.A2(n_34),
.B1(n_36),
.B2(n_60),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_135),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_111),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_21),
.B(n_111),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_96),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_25),
.A2(n_33),
.B1(n_152),
.B2(n_186),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_25),
.A2(n_154),
.B(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_26),
.A2(n_38),
.B1(n_59),
.B2(n_61),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_26),
.A2(n_59),
.B1(n_61),
.B2(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_26),
.A2(n_151),
.B(n_153),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_26),
.B(n_155),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_28),
.A2(n_73),
.B(n_159),
.Y(n_158)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_29),
.B(n_204),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_33),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_33),
.A2(n_175),
.B(n_186),
.Y(n_185)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_34),
.B(n_215),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_46),
.B(n_47),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_43),
.A2(n_46),
.B1(n_56),
.B2(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_43),
.A2(n_159),
.B(n_192),
.Y(n_216)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_44),
.A2(n_45),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_44),
.A2(n_45),
.B1(n_133),
.B2(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_44),
.B(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_44),
.A2(n_190),
.B(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_44),
.A2(n_45),
.B1(n_190),
.B2(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_45),
.A2(n_149),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_45),
.B(n_163),
.Y(n_192)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_46),
.A2(n_162),
.B(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_62),
.B1(n_63),
.B2(n_95),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_54),
.A2(n_57),
.B1(n_58),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_61),
.B(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_78),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_65),
.A2(n_124),
.B(n_126),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_65),
.A2(n_126),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_66),
.A2(n_72),
.B1(n_125),
.B2(n_143),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_68),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

AOI32xp33_ASAP7_75t_L g128 ( 
.A1(n_67),
.A2(n_82),
.A3(n_87),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g130 ( 
.A(n_68),
.B(n_88),
.Y(n_130)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_106),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_76),
.B(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_76),
.A2(n_105),
.B(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_84),
.B(n_91),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_85),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_83),
.B1(n_87),
.B2(n_88),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_82),
.A2(n_84),
.B(n_159),
.C(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_92),
.B(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_103),
.C(n_107),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_98),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_99),
.B(n_101),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_100),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_102),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_104),
.B1(n_107),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_118),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_112),
.B(n_116),
.Y(n_239)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_118),
.B(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.C(n_127),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_119),
.B(n_123),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_127),
.B(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_131),
.B1(n_132),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI31xp33_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_236),
.A3(n_246),
.B(n_251),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_180),
.B(n_235),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_164),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_139),
.B(n_164),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_150),
.C(n_156),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_140),
.B(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_145),
.C(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_150),
.B(n_156),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_160),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_176),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_165),
.B(n_177),
.C(n_179),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_166),
.B(n_171),
.C(n_172),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_230),
.B(n_234),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_199),
.B(n_229),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_193),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_193),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_188),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_189),
.B1(n_208),
.B2(n_210),
.Y(n_207)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_197),
.C(n_198),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_211),
.B(n_228),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_207),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_208),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_222),
.B(n_227),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_217),
.B(n_221),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_220),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_219),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_225),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_233),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_240),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.C(n_244),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_243),
.Y(n_249)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_250),
.Y(n_252)
);


endmodule