module fake_jpeg_9576_n_38 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_5),
.B(n_0),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVxp67_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx8_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

AND2x2_ASAP7_75t_SL g14 ( 
.A(n_13),
.B(n_0),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_14),
.A2(n_18),
.B(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_1),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_17),
.B(n_19),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_10),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_3),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_20),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

OA21x2_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_13),
.B(n_7),
.Y(n_30)
);

BUFx24_ASAP7_75t_SL g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_14),
.C(n_17),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_21),
.C(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_25),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_34),
.B(n_28),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_33),
.B(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_36),
.B(n_34),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_6),
.B1(n_12),
.B2(n_22),
.Y(n_38)
);


endmodule