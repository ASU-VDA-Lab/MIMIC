module fake_jpeg_1843_n_536 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_536);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_536;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_7),
.B(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_49),
.Y(n_133)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_51),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_53),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_14),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_54),
.B(n_82),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_59),
.B(n_81),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_60),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_62),
.Y(n_118)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_64),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_72),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_76),
.B(n_78),
.Y(n_149)
);

HAxp5_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_0),
.CON(n_77),
.SN(n_77)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_77),
.A2(n_30),
.B(n_33),
.Y(n_123)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_15),
.B(n_14),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_17),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_84),
.Y(n_128)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_17),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_90),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_13),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_89),
.B(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_45),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

CKINVDCx6p67_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_18),
.B(n_13),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_32),
.B1(n_37),
.B2(n_19),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_106),
.A2(n_116),
.B1(n_30),
.B2(n_37),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx11_ASAP7_75t_L g207 ( 
.A(n_109),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_77),
.B(n_39),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_114),
.B(n_144),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_46),
.A2(n_37),
.B1(n_32),
.B2(n_38),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_123),
.B(n_125),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_39),
.Y(n_125)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_130),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

BUFx2_ASAP7_75t_R g134 ( 
.A(n_55),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_134),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_74),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_62),
.B(n_38),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_148),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_63),
.B(n_18),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_156),
.Y(n_187)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_56),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_92),
.A2(n_37),
.B1(n_32),
.B2(n_19),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_35),
.B1(n_65),
.B2(n_73),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_78),
.B(n_45),
.C(n_29),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_0),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_95),
.B(n_31),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_96),
.B(n_31),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_57),
.Y(n_191)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_162),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_L g163 ( 
.A1(n_106),
.A2(n_97),
.B1(n_67),
.B2(n_80),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_163),
.A2(n_170),
.B1(n_182),
.B2(n_137),
.Y(n_222)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_99),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_164),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_167),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

O2A1O1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_30),
.B(n_85),
.C(n_29),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_33),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_185),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_L g233 ( 
.A1(n_172),
.A2(n_196),
.B1(n_204),
.B2(n_117),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_119),
.A2(n_60),
.B1(n_52),
.B2(n_53),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_173),
.A2(n_189),
.B1(n_161),
.B2(n_111),
.Y(n_226)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_175),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_121),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_193),
.Y(n_223)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_102),
.Y(n_177)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

INVx13_ASAP7_75t_L g244 ( 
.A(n_179),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_184),
.B(n_191),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_140),
.B(n_98),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_110),
.B(n_69),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_198),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_71),
.B1(n_75),
.B2(n_79),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_118),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_192),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_135),
.B(n_57),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_139),
.B(n_157),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_200),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_108),
.A2(n_35),
.B1(n_56),
.B2(n_79),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_103),
.B(n_133),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_138),
.B(n_159),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_0),
.Y(n_245)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_201),
.Y(n_221)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_99),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_203),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_8),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_108),
.A2(n_35),
.B1(n_27),
.B2(n_26),
.Y(n_204)
);

NAND2x1_ASAP7_75t_SL g205 ( 
.A(n_130),
.B(n_27),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_205),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_SL g206 ( 
.A1(n_101),
.A2(n_27),
.B(n_26),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_206),
.B(n_102),
.Y(n_220)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_118),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_122),
.B1(n_132),
.B2(n_127),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_215),
.A2(n_226),
.B1(n_228),
.B2(n_214),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_222),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_172),
.A2(n_142),
.B1(n_111),
.B2(n_155),
.Y(n_224)
);

AO22x1_ASAP7_75t_SL g248 ( 
.A1(n_224),
.A2(n_239),
.B1(n_192),
.B2(n_181),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_189),
.A2(n_136),
.B1(n_158),
.B2(n_129),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_190),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_241),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_163),
.A2(n_197),
.B1(n_184),
.B2(n_198),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_232),
.A2(n_240),
.B1(n_192),
.B2(n_176),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_166),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_184),
.A2(n_161),
.B1(n_155),
.B2(n_158),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_199),
.A2(n_137),
.B1(n_141),
.B2(n_146),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_190),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_180),
.B(n_102),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_242),
.B(n_168),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_245),
.B(n_175),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_274),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_223),
.Y(n_249)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_252),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_187),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_220),
.A2(n_206),
.B(n_205),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_254),
.A2(n_217),
.B(n_239),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_171),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_259),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_218),
.Y(n_257)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_257),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_258),
.A2(n_269),
.B1(n_221),
.B2(n_214),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_213),
.B(n_195),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_213),
.B(n_185),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_262),
.Y(n_295)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_227),
.Y(n_262)
);

OAI32xp33_ASAP7_75t_L g263 ( 
.A1(n_211),
.A2(n_195),
.A3(n_170),
.B1(n_188),
.B2(n_209),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_264),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_205),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_166),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_265),
.B(n_266),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_174),
.Y(n_266)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_236),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_268),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_232),
.A2(n_170),
.B1(n_115),
.B2(n_146),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_211),
.B(n_186),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_271),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_223),
.B(n_208),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_227),
.Y(n_272)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_272),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_273),
.A2(n_246),
.B1(n_178),
.B2(n_177),
.Y(n_302)
);

INVx3_ASAP7_75t_SL g274 ( 
.A(n_219),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_200),
.Y(n_275)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

INVx11_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_276),
.A2(n_214),
.B1(n_229),
.B2(n_241),
.Y(n_282)
);

AND2x6_ASAP7_75t_L g277 ( 
.A(n_218),
.B(n_162),
.Y(n_277)
);

AOI32xp33_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_242),
.A3(n_217),
.B1(n_225),
.B2(n_246),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_235),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_278),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_225),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_296),
.C(n_264),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_283),
.A2(n_302),
.B(n_305),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_253),
.A2(n_270),
.B1(n_222),
.B2(n_249),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_286),
.A2(n_294),
.B1(n_300),
.B2(n_304),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_253),
.A2(n_226),
.B1(n_240),
.B2(n_224),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_259),
.B(n_238),
.C(n_216),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_261),
.Y(n_303)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_253),
.A2(n_221),
.B1(n_167),
.B2(n_201),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_254),
.A2(n_178),
.B(n_216),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_253),
.A2(n_247),
.B1(n_219),
.B2(n_181),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_306),
.A2(n_278),
.B1(n_274),
.B2(n_276),
.Y(n_334)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_275),
.Y(n_307)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_307),
.Y(n_315)
);

AND2x2_ASAP7_75t_SL g310 ( 
.A(n_257),
.B(n_264),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_310),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_277),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_311),
.A2(n_323),
.B(n_325),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_283),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_289),
.B(n_255),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_316),
.B(n_319),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_309),
.Y(n_318)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_318),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_293),
.Y(n_319)
);

NOR3xp33_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_254),
.C(n_273),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_322),
.B(n_324),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_305),
.A2(n_273),
.B(n_277),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_291),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_285),
.A2(n_273),
.B(n_263),
.Y(n_325)
);

OAI32xp33_ASAP7_75t_L g326 ( 
.A1(n_295),
.A2(n_270),
.A3(n_262),
.B1(n_252),
.B2(n_263),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_326),
.A2(n_309),
.B(n_288),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_300),
.A2(n_267),
.B1(n_268),
.B2(n_248),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_328),
.A2(n_329),
.B1(n_286),
.B2(n_290),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_285),
.A2(n_248),
.B1(n_251),
.B2(n_258),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_297),
.B(n_271),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_330),
.B(n_331),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_266),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_281),
.Y(n_332)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_332),
.Y(n_356)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_333),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_334),
.A2(n_285),
.B1(n_308),
.B2(n_284),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_279),
.B(n_266),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_335),
.B(n_336),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_279),
.B(n_256),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_285),
.A2(n_250),
.B(n_275),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_337),
.A2(n_307),
.B(n_288),
.Y(n_364)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_299),
.Y(n_338)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_338),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_290),
.Y(n_339)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_339),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_289),
.B(n_250),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_341),
.B(n_342),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_298),
.B(n_265),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_258),
.Y(n_343)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_343),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_316),
.B(n_287),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_346),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_296),
.C(n_280),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_348),
.C(n_355),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_330),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_350),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_319),
.B(n_287),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_337),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_351),
.B(n_363),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_312),
.B(n_310),
.C(n_295),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_360),
.A2(n_376),
.B1(n_329),
.B2(n_337),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_361),
.A2(n_368),
.B1(n_372),
.B2(n_315),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_298),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_364),
.A2(n_317),
.B(n_325),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_318),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_338),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_310),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_366),
.B(n_335),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_310),
.C(n_303),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_374),
.C(n_317),
.Y(n_387)
);

AOI21xp33_ASAP7_75t_L g370 ( 
.A1(n_321),
.A2(n_304),
.B(n_306),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_370),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_328),
.A2(n_294),
.B1(n_284),
.B2(n_269),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_333),
.Y(n_373)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_373),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_308),
.C(n_302),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_313),
.Y(n_375)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_375),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_340),
.A2(n_248),
.B1(n_269),
.B2(n_274),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_348),
.B(n_326),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_377),
.B(n_393),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_361),
.A2(n_340),
.B1(n_343),
.B2(n_325),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_378),
.A2(n_375),
.B1(n_356),
.B2(n_247),
.Y(n_429)
);

BUFx5_ASAP7_75t_L g379 ( 
.A(n_354),
.Y(n_379)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_379),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_381),
.A2(n_389),
.B1(n_398),
.B2(n_405),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_384),
.A2(n_373),
.B(n_357),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_349),
.B(n_342),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_385),
.B(n_396),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_387),
.B(n_374),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_376),
.A2(n_323),
.B1(n_315),
.B2(n_322),
.Y(n_389)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_390),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_362),
.B(n_331),
.Y(n_391)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_391),
.Y(n_409)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_345),
.Y(n_392)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_392),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_347),
.B(n_311),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_404),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_345),
.B(n_238),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_367),
.A2(n_320),
.B1(n_311),
.B2(n_332),
.Y(n_398)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_399),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_352),
.B(n_314),
.Y(n_400)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_400),
.Y(n_417)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_357),
.Y(n_401)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_401),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_355),
.B(n_369),
.C(n_351),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_344),
.C(n_364),
.Y(n_418)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_352),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_403),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_368),
.B(n_314),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_371),
.A2(n_313),
.B1(n_334),
.B2(n_274),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_362),
.B(n_248),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_366),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_407),
.B(n_424),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_381),
.A2(n_367),
.B1(n_372),
.B2(n_344),
.Y(n_411)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_411),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_388),
.B(n_371),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_414),
.Y(n_445)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_416),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_418),
.B(n_423),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_398),
.A2(n_353),
.B1(n_358),
.B2(n_359),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_422),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_380),
.A2(n_353),
.B1(n_358),
.B2(n_359),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_391),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_382),
.B(n_360),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_404),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_231),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_428),
.A2(n_378),
.B(n_393),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_429),
.A2(n_405),
.B1(n_383),
.B2(n_389),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_387),
.B(n_356),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_430),
.B(n_402),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_382),
.B(n_235),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_432),
.B(n_433),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_395),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_394),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_436),
.B(n_446),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_441),
.Y(n_459)
);

O2A1O1Ixp33_ASAP7_75t_L g438 ( 
.A1(n_408),
.A2(n_397),
.B(n_384),
.C(n_406),
.Y(n_438)
);

O2A1O1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_438),
.A2(n_100),
.B(n_165),
.C(n_169),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_424),
.B(n_377),
.Y(n_441)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_444),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_410),
.A2(n_379),
.B1(n_386),
.B2(n_401),
.Y(n_446)
);

OAI21xp33_ASAP7_75t_L g467 ( 
.A1(n_447),
.A2(n_448),
.B(n_455),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_422),
.A2(n_212),
.B(n_276),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_212),
.C(n_235),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_449),
.B(n_452),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_417),
.A2(n_247),
.B1(n_237),
.B2(n_183),
.Y(n_450)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_450),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_419),
.B(n_237),
.Y(n_451)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_451),
.Y(n_474)
);

OAI21xp33_ASAP7_75t_L g452 ( 
.A1(n_421),
.A2(n_164),
.B(n_244),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_231),
.C(n_202),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_453),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_190),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_454),
.B(n_457),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_428),
.A2(n_237),
.B(n_244),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_456),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_429),
.B(n_141),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_419),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_461),
.B(n_463),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_418),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_440),
.A2(n_413),
.B1(n_431),
.B2(n_409),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_464),
.B(n_468),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_431),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_466),
.B(n_469),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_440),
.A2(n_416),
.B1(n_427),
.B2(n_411),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_443),
.A2(n_420),
.B1(n_415),
.B2(n_425),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_435),
.B(n_407),
.C(n_425),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_476),
.Y(n_488)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_475),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_435),
.B(n_447),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_434),
.B(n_210),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_477),
.B(n_449),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_470),
.B(n_443),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_478),
.B(n_480),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_476),
.B(n_454),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_482),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_474),
.B(n_439),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_463),
.B(n_453),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_481),
.B(n_131),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_459),
.B(n_439),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_459),
.B(n_441),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_483),
.B(n_490),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_465),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_487),
.B(n_489),
.Y(n_497)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_460),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_SL g490 ( 
.A1(n_472),
.A2(n_457),
.B1(n_448),
.B2(n_438),
.Y(n_490)
);

OAI21x1_ASAP7_75t_SL g491 ( 
.A1(n_473),
.A2(n_457),
.B(n_456),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_491),
.A2(n_455),
.B(n_467),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_493),
.B(n_494),
.Y(n_499)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_475),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_471),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_498),
.B(n_508),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_500),
.A2(n_501),
.B1(n_131),
.B2(n_109),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_486),
.A2(n_467),
.B1(n_462),
.B2(n_120),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_487),
.B(n_462),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_502),
.A2(n_503),
.B1(n_505),
.B2(n_34),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_484),
.A2(n_107),
.B(n_210),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_100),
.C(n_115),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_504),
.B(n_179),
.C(n_109),
.Y(n_514)
);

AOI321xp33_ASAP7_75t_L g507 ( 
.A1(n_485),
.A2(n_483),
.A3(n_492),
.B1(n_490),
.B2(n_479),
.C(n_207),
.Y(n_507)
);

AOI31xp67_ASAP7_75t_L g517 ( 
.A1(n_507),
.A2(n_504),
.A3(n_12),
.B(n_8),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_488),
.B(n_207),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_496),
.B(n_112),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_509),
.B(n_512),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_502),
.Y(n_510)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_510),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_112),
.Y(n_511)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_511),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_499),
.A2(n_497),
.B1(n_506),
.B2(n_495),
.Y(n_512)
);

XNOR2x1_ASAP7_75t_L g525 ( 
.A(n_513),
.B(n_514),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_515),
.A2(n_517),
.B(n_519),
.Y(n_526)
);

AOI322xp5_ASAP7_75t_L g516 ( 
.A1(n_506),
.A2(n_34),
.A3(n_26),
.B1(n_12),
.B2(n_11),
.C1(n_10),
.C2(n_8),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_516),
.B(n_12),
.C(n_1),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_499),
.A2(n_34),
.B1(n_12),
.B2(n_2),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_521),
.A2(n_523),
.B(n_514),
.Y(n_527)
);

NOR3xp33_ASAP7_75t_SL g523 ( 
.A(n_510),
.B(n_518),
.C(n_511),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_527),
.A2(n_530),
.B1(n_524),
.B2(n_525),
.Y(n_532)
);

AO21x1_ASAP7_75t_L g528 ( 
.A1(n_522),
.A2(n_0),
.B(n_1),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_528),
.A2(n_529),
.B(n_526),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_520),
.A2(n_1),
.B(n_2),
.Y(n_529)
);

AOI322xp5_ASAP7_75t_L g530 ( 
.A1(n_523),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_530)
);

AO21x1_ASAP7_75t_L g533 ( 
.A1(n_531),
.A2(n_532),
.B(n_7),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_533),
.A2(n_1),
.B(n_2),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_3),
.B(n_4),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_6),
.Y(n_536)
);


endmodule