module fake_jpeg_6436_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_42),
.B1(n_29),
.B2(n_27),
.Y(n_56)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_47),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_53),
.Y(n_93)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx2_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_54),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_29),
.B1(n_20),
.B2(n_21),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_19),
.B1(n_23),
.B2(n_20),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_33),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_71),
.Y(n_86)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_42),
.B1(n_47),
.B2(n_44),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_33),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_40),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_72),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_29),
.B1(n_31),
.B2(n_26),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_20),
.B1(n_19),
.B2(n_23),
.Y(n_89)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_80),
.Y(n_105)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_89),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_42),
.B1(n_47),
.B2(n_30),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_41),
.B1(n_46),
.B2(n_47),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_100),
.B1(n_21),
.B2(n_19),
.Y(n_125)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_70),
.A2(n_30),
.B1(n_46),
.B2(n_44),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_33),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_23),
.Y(n_116)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_102),
.Y(n_131)
);

BUFx10_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_55),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_128),
.Y(n_148)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_109),
.B(n_114),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_52),
.B(n_71),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_98),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_93),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_111),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_61),
.B1(n_44),
.B2(n_46),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_118),
.B1(n_30),
.B2(n_22),
.Y(n_149)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_82),
.B(n_65),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_57),
.B(n_21),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_75),
.A2(n_40),
.B1(n_44),
.B2(n_41),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_43),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_82),
.B(n_31),
.Y(n_124)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_125),
.A2(n_90),
.B1(n_80),
.B2(n_22),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_79),
.B(n_45),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_126),
.B(n_37),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_127),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_98),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_75),
.B(n_53),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_92),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_88),
.B1(n_41),
.B2(n_79),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_134),
.A2(n_135),
.B1(n_143),
.B2(n_147),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_41),
.B1(n_77),
.B2(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_137),
.B(n_139),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_138),
.B(n_48),
.Y(n_183)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g168 ( 
.A(n_140),
.B(n_156),
.CI(n_129),
.CON(n_168),
.SN(n_168)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_77),
.B1(n_99),
.B2(n_76),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_152),
.B1(n_155),
.B2(n_101),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_142),
.B(n_145),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_91),
.B1(n_83),
.B2(n_84),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_84),
.B1(n_51),
.B2(n_50),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_130),
.B1(n_123),
.B2(n_107),
.Y(n_177)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_151),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_106),
.A2(n_43),
.B1(n_60),
.B2(n_49),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_68),
.C(n_45),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_154),
.C(n_126),
.Y(n_163)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_48),
.C(n_43),
.Y(n_154)
);

AO22x1_ASAP7_75t_SL g155 ( 
.A1(n_119),
.A2(n_43),
.B1(n_60),
.B2(n_49),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_164),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_161),
.B(n_176),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_162),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_169),
.C(n_175),
.Y(n_195)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_171),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_155),
.A2(n_119),
.B1(n_128),
.B2(n_108),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_187),
.B(n_146),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_110),
.B1(n_111),
.B2(n_126),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_172),
.B1(n_140),
.B2(n_137),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_182),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_122),
.C(n_114),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_158),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_106),
.B1(n_124),
.B2(n_123),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_181),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_26),
.B(n_113),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_183),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_68),
.C(n_45),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_157),
.B1(n_104),
.B2(n_102),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_48),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_146),
.C(n_150),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_136),
.B(n_130),
.Y(n_181)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_148),
.B(n_45),
.CI(n_48),
.CON(n_182),
.SN(n_182)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_186),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_144),
.A2(n_63),
.A3(n_17),
.B1(n_28),
.B2(n_34),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_102),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_134),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_25),
.B(n_45),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_191),
.Y(n_219)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_193),
.A2(n_196),
.B(n_204),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_133),
.C(n_154),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_194),
.B(n_203),
.Y(n_236)
);

HAxp5_ASAP7_75t_SL g196 ( 
.A(n_165),
.B(n_145),
.CON(n_196),
.SN(n_196)
);

OA22x2_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_135),
.B1(n_141),
.B2(n_152),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_197),
.A2(n_214),
.B1(n_169),
.B2(n_175),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_208),
.C(n_212),
.Y(n_225)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_166),
.A2(n_136),
.B(n_25),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_206),
.Y(n_241)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_68),
.C(n_45),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_172),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_209),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_163),
.B(n_68),
.C(n_45),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_182),
.B(n_0),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_179),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_162),
.A2(n_176),
.B1(n_184),
.B2(n_182),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_215),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_216),
.B(n_217),
.Y(n_265)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_223),
.Y(n_245)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_168),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_231),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_205),
.B1(n_206),
.B2(n_199),
.Y(n_243)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_188),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_232),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_210),
.A2(n_168),
.B(n_161),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_229),
.B(n_236),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_183),
.C(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_235),
.A2(n_242),
.B(n_209),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_189),
.B(n_159),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_238),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_102),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_102),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_201),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_197),
.Y(n_240)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_243),
.A2(n_17),
.B1(n_34),
.B2(n_28),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_246),
.A2(n_255),
.B(n_261),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_215),
.B1(n_197),
.B2(n_190),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_248),
.A2(n_251),
.B1(n_231),
.B2(n_225),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_233),
.A2(n_191),
.B1(n_213),
.B2(n_203),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_218),
.A2(n_193),
.B1(n_204),
.B2(n_212),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_257),
.Y(n_268)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_219),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_258),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_211),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_230),
.A2(n_208),
.B(n_2),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_220),
.A2(n_226),
.B1(n_221),
.B2(n_228),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_240),
.A2(n_157),
.B1(n_104),
.B2(n_115),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_229),
.A2(n_115),
.B1(n_17),
.B2(n_28),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_266),
.B(n_269),
.Y(n_295)
);

XNOR2x1_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_227),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_225),
.C(n_238),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_272),
.C(n_281),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_239),
.C(n_217),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_216),
.Y(n_273)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_245),
.B(n_223),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_280),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_222),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_276),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_278),
.B(n_279),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_247),
.A2(n_115),
.B1(n_34),
.B2(n_28),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_25),
.C(n_18),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_243),
.B(n_25),
.C(n_18),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_284),
.C(n_281),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_252),
.A2(n_18),
.B1(n_2),
.B2(n_3),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_250),
.B1(n_261),
.B2(n_255),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_25),
.C(n_18),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_287),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_257),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_292),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_253),
.Y(n_289)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_289),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_248),
.Y(n_292)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_293),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g297 ( 
.A(n_266),
.B(n_251),
.CI(n_264),
.CON(n_297),
.SN(n_297)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_297),
.B(n_299),
.Y(n_304)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_298),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_267),
.B(n_8),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_277),
.A2(n_274),
.B1(n_273),
.B2(n_282),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_300),
.A2(n_283),
.B1(n_284),
.B2(n_272),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_302),
.A2(n_303),
.B(n_306),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_296),
.A2(n_271),
.B(n_9),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_16),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_311),
.C(n_295),
.Y(n_315)
);

AND2x4_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_1),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_307),
.A2(n_310),
.B1(n_313),
.B2(n_8),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_298),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_315),
.A2(n_13),
.B(n_16),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_285),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_320),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_SL g318 ( 
.A(n_306),
.B(n_297),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_306),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_290),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_319),
.A2(n_321),
.B(n_322),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_290),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_303),
.A2(n_288),
.B(n_10),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_10),
.C(n_15),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_10),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_8),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_324),
.A2(n_312),
.B1(n_314),
.B2(n_305),
.Y(n_328)
);

AO21x1_ASAP7_75t_L g335 ( 
.A1(n_326),
.A2(n_4),
.B(n_5),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_316),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_329),
.B(n_331),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_320),
.A2(n_11),
.B(n_15),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_332),
.C(n_5),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_13),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_333),
.A2(n_334),
.B(n_325),
.Y(n_339)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_325),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_337),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_327),
.B(n_336),
.Y(n_340)
);

AOI321xp33_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_6),
.A3(n_7),
.B1(n_326),
.B2(n_338),
.C(n_333),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_341),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_6),
.B(n_7),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_6),
.Y(n_344)
);


endmodule