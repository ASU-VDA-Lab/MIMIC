module fake_netlist_1_5158_n_554 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_554);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_554;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_22), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_50), .Y(n_80) );
BUFx5_ASAP7_75t_L g81 ( .A(n_5), .Y(n_81) );
OR2x2_ASAP7_75t_L g82 ( .A(n_69), .B(n_42), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_44), .Y(n_83) );
INVx1_ASAP7_75t_SL g84 ( .A(n_39), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_13), .Y(n_85) );
BUFx2_ASAP7_75t_SL g86 ( .A(n_21), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_67), .Y(n_87) );
BUFx2_ASAP7_75t_L g88 ( .A(n_73), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_58), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_18), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_6), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_19), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_53), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_63), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_1), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_77), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_41), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_0), .Y(n_98) );
BUFx6f_ASAP7_75t_L g99 ( .A(n_65), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_1), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_60), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_61), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_34), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_54), .Y(n_104) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_10), .Y(n_105) );
BUFx10_ASAP7_75t_L g106 ( .A(n_32), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_38), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_49), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_23), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_31), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_62), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_72), .Y(n_113) );
INVxp33_ASAP7_75t_L g114 ( .A(n_64), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_16), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_74), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_98), .Y(n_117) );
OAI21x1_ASAP7_75t_L g118 ( .A1(n_97), .A2(n_30), .B(n_76), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_114), .B(n_0), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_81), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_106), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_81), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_81), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_99), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_81), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_88), .B(n_2), .Y(n_126) );
NOR2x1_ASAP7_75t_L g127 ( .A(n_79), .B(n_3), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_97), .B(n_3), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_81), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_99), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_104), .B(n_4), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_80), .B(n_4), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_98), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_114), .B(n_7), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_81), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_81), .Y(n_136) );
BUFx8_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_99), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_87), .Y(n_139) );
BUFx10_ASAP7_75t_L g140 ( .A(n_126), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_121), .B(n_83), .Y(n_141) );
INVx5_ASAP7_75t_L g142 ( .A(n_124), .Y(n_142) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_117), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_120), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_120), .Y(n_145) );
NAND2xp33_ASAP7_75t_L g146 ( .A(n_121), .B(n_90), .Y(n_146) );
INVx4_ASAP7_75t_L g147 ( .A(n_128), .Y(n_147) );
NOR2x1p5_ASAP7_75t_L g148 ( .A(n_121), .B(n_100), .Y(n_148) );
NAND2xp33_ASAP7_75t_L g149 ( .A(n_121), .B(n_108), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_122), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_124), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_126), .B(n_106), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_122), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_119), .B(n_106), .Y(n_154) );
NOR2x1p5_ASAP7_75t_L g155 ( .A(n_132), .B(n_100), .Y(n_155) );
NAND2x1_ASAP7_75t_L g156 ( .A(n_128), .B(n_104), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_125), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_125), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_124), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_128), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_126), .B(n_85), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_128), .A2(n_95), .B1(n_112), .B2(n_91), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_131), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g164 ( .A1(n_133), .A2(n_115), .B1(n_92), .B2(n_101), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_126), .B(n_94), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_160), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_140), .B(n_137), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_154), .B(n_119), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_141), .B(n_137), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_154), .B(n_134), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_144), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_161), .B(n_134), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_155), .A2(n_137), .B1(n_131), .B2(n_101), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_160), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_161), .B(n_137), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_160), .A2(n_139), .B(n_131), .C(n_123), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_160), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_140), .B(n_131), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_161), .B(n_139), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_148), .B(n_127), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_161), .B(n_94), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_156), .Y(n_183) );
BUFx2_ASAP7_75t_L g184 ( .A(n_143), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_155), .A2(n_92), .B1(n_133), .B2(n_127), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_147), .A2(n_135), .B1(n_123), .B2(n_129), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_148), .B(n_118), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_147), .B(n_135), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_147), .A2(n_136), .B1(n_129), .B2(n_105), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_140), .B(n_136), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_163), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_152), .B(n_107), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_140), .B(n_84), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_165), .B(n_109), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_146), .B(n_86), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_163), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_162), .A2(n_115), .B1(n_89), .B2(n_111), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_163), .A2(n_105), .B1(n_93), .B2(n_103), .Y(n_198) );
NAND2x1p5_ASAP7_75t_L g199 ( .A(n_156), .B(n_163), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_196), .Y(n_200) );
BUFx4f_ASAP7_75t_L g201 ( .A(n_184), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_196), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_170), .B(n_149), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_168), .B(n_150), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_184), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_168), .A2(n_164), .B1(n_144), .B2(n_158), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_185), .A2(n_164), .B1(n_145), .B2(n_158), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_183), .B(n_157), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_176), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_172), .B(n_150), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_176), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_197), .B(n_8), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_196), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_188), .A2(n_145), .B(n_157), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_177), .A2(n_153), .B(n_118), .C(n_96), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_181), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_183), .B(n_153), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_166), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_179), .A2(n_116), .B(n_102), .Y(n_219) );
NOR3xp33_ASAP7_75t_SL g220 ( .A(n_169), .B(n_110), .C(n_113), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_166), .Y(n_221) );
NOR3xp33_ASAP7_75t_SL g222 ( .A(n_167), .B(n_193), .C(n_175), .Y(n_222) );
INVx4_ASAP7_75t_L g223 ( .A(n_176), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_171), .Y(n_224) );
NAND2xp33_ASAP7_75t_SL g225 ( .A(n_183), .B(n_105), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_183), .B(n_99), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_180), .A2(n_159), .B(n_151), .C(n_105), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_174), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_173), .A2(n_138), .B1(n_130), .B2(n_124), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_174), .A2(n_159), .B(n_151), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_183), .B(n_142), .Y(n_231) );
NOR2xp33_ASAP7_75t_SL g232 ( .A(n_187), .B(n_138), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_205), .B(n_181), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_212), .A2(n_181), .B1(n_178), .B2(n_191), .Y(n_234) );
AO32x2_ASAP7_75t_L g235 ( .A1(n_229), .A2(n_198), .A3(n_215), .B1(n_220), .B2(n_223), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_224), .Y(n_236) );
BUFx3_ASAP7_75t_L g237 ( .A(n_201), .Y(n_237) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_214), .A2(n_187), .B(n_191), .Y(n_238) );
AO31x2_ASAP7_75t_L g239 ( .A1(n_203), .A2(n_171), .A3(n_178), .B(n_195), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_208), .A2(n_187), .B(n_199), .Y(n_240) );
AOI22x1_ASAP7_75t_L g241 ( .A1(n_219), .A2(n_199), .B1(n_190), .B2(n_124), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_205), .B(n_182), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_203), .A2(n_194), .B1(n_199), .B2(n_190), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_204), .A2(n_192), .B1(n_189), .B2(n_186), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_218), .Y(n_245) );
INVxp67_ASAP7_75t_SL g246 ( .A(n_201), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_206), .A2(n_124), .B1(n_130), .B2(n_138), .Y(n_247) );
AO31x2_ASAP7_75t_L g248 ( .A1(n_221), .A2(n_159), .A3(n_151), .B(n_138), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_207), .A2(n_138), .B1(n_130), .B2(n_142), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_SL g250 ( .A1(n_226), .A2(n_40), .B(n_78), .C(n_75), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_208), .A2(n_142), .B(n_138), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_216), .B(n_8), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_228), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_210), .A2(n_142), .B(n_130), .Y(n_254) );
AOI221xp5_ASAP7_75t_L g255 ( .A1(n_220), .A2(n_130), .B1(n_10), .B2(n_11), .C(n_12), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_SL g256 ( .A1(n_226), .A2(n_37), .B(n_71), .C(n_70), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_211), .A2(n_130), .B1(n_142), .B2(n_12), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_222), .A2(n_142), .B(n_11), .C(n_13), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_217), .A2(n_142), .B(n_36), .Y(n_259) );
NAND2xp33_ASAP7_75t_L g260 ( .A(n_222), .B(n_35), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_234), .B(n_211), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_237), .Y(n_262) );
OA21x2_ASAP7_75t_L g263 ( .A1(n_238), .A2(n_217), .B(n_230), .Y(n_263) );
INVx2_ASAP7_75t_SL g264 ( .A(n_237), .Y(n_264) );
NOR2xp67_ASAP7_75t_L g265 ( .A(n_240), .B(n_223), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_260), .A2(n_232), .B(n_227), .Y(n_266) );
OA21x2_ASAP7_75t_L g267 ( .A1(n_254), .A2(n_200), .B(n_231), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_253), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_234), .B(n_213), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_242), .B(n_202), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_245), .B(n_209), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_236), .B(n_209), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_241), .A2(n_231), .B(n_225), .Y(n_273) );
OAI21x1_ASAP7_75t_SL g274 ( .A1(n_257), .A2(n_9), .B(n_14), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_239), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_239), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_233), .B(n_9), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_243), .B(n_14), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_243), .A2(n_45), .B(n_66), .Y(n_279) );
OA21x2_ASAP7_75t_L g280 ( .A1(n_258), .A2(n_43), .B(n_59), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_255), .A2(n_15), .B(n_16), .C(n_17), .Y(n_281) );
AOI21xp33_ASAP7_75t_L g282 ( .A1(n_252), .A2(n_15), .B(n_17), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_246), .A2(n_20), .B1(n_24), .B2(n_25), .C(n_26), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_275), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_271), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_275), .Y(n_286) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_276), .A2(n_274), .B(n_266), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_268), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_268), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_276), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_262), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_267), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_267), .B(n_235), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_265), .B(n_239), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_267), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_267), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_263), .B(n_271), .Y(n_297) );
AO21x1_ASAP7_75t_SL g298 ( .A1(n_261), .A2(n_257), .B(n_249), .Y(n_298) );
INVx2_ASAP7_75t_SL g299 ( .A(n_262), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_263), .Y(n_300) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_265), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_263), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_263), .B(n_235), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_278), .B(n_239), .Y(n_304) );
OAI221xp5_ASAP7_75t_L g305 ( .A1(n_281), .A2(n_244), .B1(n_247), .B2(n_259), .C(n_251), .Y(n_305) );
BUFx3_ASAP7_75t_L g306 ( .A(n_262), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_300), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_294), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_286), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_303), .B(n_235), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_303), .B(n_235), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_303), .B(n_280), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_306), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_297), .B(n_280), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_294), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_294), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_297), .B(n_248), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_286), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_300), .Y(n_319) );
NOR2x1_ASAP7_75t_SL g320 ( .A(n_306), .B(n_269), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_284), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_290), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_300), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_297), .B(n_280), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_290), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_294), .Y(n_326) );
INVx5_ASAP7_75t_L g327 ( .A(n_299), .Y(n_327) );
INVx5_ASAP7_75t_SL g328 ( .A(n_294), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_284), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_284), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_288), .B(n_277), .Y(n_331) );
AOI33xp33_ASAP7_75t_L g332 ( .A1(n_288), .A2(n_264), .A3(n_244), .B1(n_271), .B2(n_272), .B3(n_283), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_293), .B(n_280), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_301), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_301), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_293), .B(n_248), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_308), .B(n_302), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_310), .B(n_293), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_322), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_309), .B(n_304), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_322), .B(n_289), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_325), .B(n_289), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_325), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_328), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_307), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_309), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_327), .B(n_291), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_310), .B(n_311), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_310), .B(n_302), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_307), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_311), .B(n_295), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_311), .B(n_295), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_336), .B(n_292), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_307), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_328), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_331), .B(n_299), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_308), .B(n_287), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_336), .B(n_292), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_319), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_331), .B(n_299), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_336), .B(n_296), .Y(n_361) );
NOR2x1_ASAP7_75t_L g362 ( .A(n_313), .B(n_306), .Y(n_362) );
INVx2_ASAP7_75t_SL g363 ( .A(n_327), .Y(n_363) );
NAND4xp25_ASAP7_75t_L g364 ( .A(n_332), .B(n_282), .C(n_304), .D(n_285), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_319), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_318), .B(n_285), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_319), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_308), .B(n_287), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_317), .B(n_296), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_318), .B(n_285), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_330), .B(n_285), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_317), .B(n_287), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_323), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_323), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_317), .B(n_287), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_335), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_330), .B(n_285), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_323), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_334), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_308), .B(n_287), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_340), .B(n_329), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_369), .B(n_317), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_369), .B(n_317), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_339), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_340), .B(n_329), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_355), .B(n_326), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_348), .B(n_264), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_339), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_362), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_355), .B(n_326), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_363), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_348), .B(n_314), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_362), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_343), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_338), .B(n_314), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_338), .B(n_314), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_353), .B(n_324), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_349), .B(n_321), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_353), .B(n_324), .Y(n_399) );
NOR3x1_ASAP7_75t_L g400 ( .A(n_347), .B(n_305), .C(n_304), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_358), .B(n_324), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_351), .B(n_335), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_343), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_356), .B(n_313), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_341), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_349), .B(n_321), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_351), .B(n_334), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_346), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_352), .B(n_333), .Y(n_409) );
BUFx2_ASAP7_75t_L g410 ( .A(n_376), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_379), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_350), .Y(n_412) );
INVx3_ASAP7_75t_SL g413 ( .A(n_363), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_379), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_342), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_352), .B(n_333), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_360), .B(n_333), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_358), .B(n_312), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_361), .B(n_308), .Y(n_419) );
NOR2xp67_ASAP7_75t_SL g420 ( .A(n_355), .B(n_327), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_345), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_361), .B(n_312), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_345), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_372), .B(n_315), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_366), .B(n_315), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_370), .B(n_312), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_371), .B(n_313), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_372), .B(n_326), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_350), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_375), .B(n_326), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_375), .B(n_326), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_378), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_337), .B(n_316), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_413), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_414), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_408), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_405), .B(n_359), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_411), .Y(n_438) );
O2A1O1Ixp33_ASAP7_75t_SL g439 ( .A1(n_393), .A2(n_355), .B(n_344), .C(n_354), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_402), .B(n_377), .Y(n_440) );
INVx1_ASAP7_75t_SL g441 ( .A(n_413), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_410), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_410), .Y(n_443) );
OAI221xp5_ASAP7_75t_SL g444 ( .A1(n_381), .A2(n_385), .B1(n_402), .B2(n_425), .C(n_407), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_394), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_389), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_382), .B(n_315), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_381), .Y(n_448) );
AOI21xp33_ASAP7_75t_SL g449 ( .A1(n_391), .A2(n_344), .B(n_380), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_389), .A2(n_320), .B(n_327), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_391), .Y(n_451) );
NAND2x1p5_ASAP7_75t_L g452 ( .A(n_420), .B(n_327), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_382), .B(n_315), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_418), .B(n_365), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_386), .B(n_327), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_394), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_403), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_383), .B(n_315), .Y(n_458) );
INVxp67_ASAP7_75t_L g459 ( .A(n_387), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_383), .B(n_316), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_385), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_405), .B(n_367), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_403), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_415), .B(n_367), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_384), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_422), .B(n_365), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_409), .B(n_354), .Y(n_467) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_412), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_388), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_392), .B(n_359), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_398), .B(n_364), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_416), .B(n_374), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_426), .B(n_374), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_406), .Y(n_474) );
INVx2_ASAP7_75t_SL g475 ( .A(n_419), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_417), .B(n_373), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_392), .B(n_373), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_419), .B(n_316), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_395), .B(n_396), .Y(n_479) );
NAND4xp25_ASAP7_75t_L g480 ( .A(n_471), .B(n_400), .C(n_404), .D(n_390), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_443), .Y(n_481) );
OAI211xp5_ASAP7_75t_L g482 ( .A1(n_441), .A2(n_344), .B(n_427), .C(n_433), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_441), .Y(n_483) );
OAI21xp33_ASAP7_75t_L g484 ( .A1(n_444), .A2(n_428), .B(n_431), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_470), .B(n_397), .Y(n_485) );
INVxp33_ASAP7_75t_L g486 ( .A(n_452), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_474), .A2(n_431), .B1(n_430), .B2(n_428), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_448), .Y(n_488) );
AOI322xp5_ASAP7_75t_L g489 ( .A1(n_479), .A2(n_396), .A3(n_395), .B1(n_397), .B2(n_401), .C1(n_399), .C2(n_430), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_464), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_464), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_437), .Y(n_492) );
OAI221xp5_ASAP7_75t_L g493 ( .A1(n_434), .A2(n_425), .B1(n_420), .B2(n_433), .C(n_423), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_437), .Y(n_494) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_452), .A2(n_327), .B1(n_316), .B2(n_386), .Y(n_495) );
OAI21xp5_ASAP7_75t_SL g496 ( .A1(n_449), .A2(n_386), .B(n_390), .Y(n_496) );
XNOR2xp5_ASAP7_75t_L g497 ( .A(n_461), .B(n_401), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_462), .Y(n_498) );
AOI221xp5_ASAP7_75t_SL g499 ( .A1(n_459), .A2(n_424), .B1(n_399), .B2(n_421), .C(n_423), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_451), .Y(n_500) );
AOI21xp33_ASAP7_75t_L g501 ( .A1(n_436), .A2(n_274), .B(n_421), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_442), .A2(n_327), .B1(n_328), .B2(n_424), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_470), .B(n_390), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_451), .Y(n_504) );
INVx1_ASAP7_75t_SL g505 ( .A(n_477), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_462), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_435), .B(n_432), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_438), .Y(n_508) );
INVxp67_ASAP7_75t_L g509 ( .A(n_446), .Y(n_509) );
AOI222xp33_ASAP7_75t_L g510 ( .A1(n_446), .A2(n_357), .B1(n_368), .B2(n_380), .C1(n_337), .C2(n_432), .Y(n_510) );
AOI211xp5_ASAP7_75t_L g511 ( .A1(n_486), .A2(n_439), .B(n_450), .C(n_455), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g512 ( .A1(n_499), .A2(n_477), .B1(n_475), .B2(n_469), .C(n_465), .Y(n_512) );
OA22x2_ASAP7_75t_L g513 ( .A1(n_496), .A2(n_453), .B1(n_447), .B2(n_458), .Y(n_513) );
AO21x1_ASAP7_75t_L g514 ( .A1(n_495), .A2(n_450), .B(n_468), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_481), .Y(n_515) );
OAI221xp5_ASAP7_75t_L g516 ( .A1(n_480), .A2(n_476), .B1(n_473), .B2(n_440), .C(n_466), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_489), .B(n_445), .Y(n_517) );
NAND2x1_ASAP7_75t_L g518 ( .A(n_502), .B(n_460), .Y(n_518) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_484), .A2(n_463), .B1(n_457), .B2(n_456), .C(n_478), .Y(n_519) );
NOR2xp67_ASAP7_75t_SL g520 ( .A(n_482), .B(n_306), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_497), .A2(n_454), .B1(n_472), .B2(n_467), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_504), .Y(n_522) );
OAI211xp5_ASAP7_75t_L g523 ( .A1(n_483), .A2(n_316), .B(n_412), .C(n_429), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_490), .Y(n_524) );
OAI221xp5_ASAP7_75t_L g525 ( .A1(n_493), .A2(n_429), .B1(n_305), .B2(n_378), .C(n_279), .Y(n_525) );
AO21x1_ASAP7_75t_L g526 ( .A1(n_502), .A2(n_380), .B(n_368), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_509), .A2(n_380), .B(n_368), .C(n_357), .Y(n_527) );
OAI211xp5_ASAP7_75t_L g528 ( .A1(n_510), .A2(n_273), .B(n_270), .C(n_256), .Y(n_528) );
OAI22xp33_ASAP7_75t_L g529 ( .A1(n_513), .A2(n_487), .B1(n_505), .B2(n_485), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g530 ( .A1(n_511), .A2(n_488), .B1(n_500), .B2(n_491), .C(n_492), .Y(n_530) );
AOI32xp33_ASAP7_75t_L g531 ( .A1(n_511), .A2(n_503), .A3(n_494), .B1(n_506), .B2(n_498), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_517), .B(n_508), .Y(n_532) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_512), .A2(n_501), .B(n_507), .Y(n_533) );
AOI221xp5_ASAP7_75t_L g534 ( .A1(n_519), .A2(n_501), .B1(n_507), .B2(n_368), .C(n_357), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_522), .B(n_357), .Y(n_535) );
OAI211xp5_ASAP7_75t_SL g536 ( .A1(n_527), .A2(n_250), .B(n_320), .C(n_298), .Y(n_536) );
AOI222xp33_ASAP7_75t_L g537 ( .A1(n_521), .A2(n_337), .B1(n_328), .B2(n_271), .C1(n_272), .C2(n_298), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_L g538 ( .A1(n_514), .A2(n_337), .B(n_298), .C(n_328), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_532), .Y(n_539) );
OAI322xp33_ASAP7_75t_L g540 ( .A1(n_529), .A2(n_518), .A3(n_516), .B1(n_524), .B2(n_525), .C1(n_515), .C2(n_526), .Y(n_540) );
NAND3xp33_ASAP7_75t_L g541 ( .A(n_531), .B(n_528), .C(n_523), .Y(n_541) );
BUFx3_ASAP7_75t_L g542 ( .A(n_535), .Y(n_542) );
OAI221xp5_ASAP7_75t_L g543 ( .A1(n_530), .A2(n_520), .B1(n_328), .B2(n_29), .C(n_33), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_539), .B(n_533), .Y(n_544) );
NAND4xp25_ASAP7_75t_SL g545 ( .A(n_541), .B(n_538), .C(n_534), .D(n_537), .Y(n_545) );
NOR5xp2_ASAP7_75t_L g546 ( .A(n_540), .B(n_536), .C(n_28), .D(n_46), .E(n_47), .Y(n_546) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_544), .A2(n_543), .B(n_542), .Y(n_547) );
BUFx2_ASAP7_75t_L g548 ( .A(n_546), .Y(n_548) );
INVx3_ASAP7_75t_SL g549 ( .A(n_548), .Y(n_549) );
AOI22x1_ASAP7_75t_L g550 ( .A1(n_549), .A2(n_545), .B1(n_547), .B2(n_51), .Y(n_550) );
OAI22xp5_ASAP7_75t_SL g551 ( .A1(n_550), .A2(n_547), .B1(n_48), .B2(n_52), .Y(n_551) );
OAI21xp5_ASAP7_75t_SL g552 ( .A1(n_551), .A2(n_27), .B(n_55), .Y(n_552) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_552), .A2(n_56), .B(n_57), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_553), .A2(n_68), .B1(n_248), .B2(n_545), .Y(n_554) );
endmodule