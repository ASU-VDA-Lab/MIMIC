module fake_netlist_6_2258_n_2258 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2258);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2258;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1317;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2209;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_SL g230 ( 
.A(n_194),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_17),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_86),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_12),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_133),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_189),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_134),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_25),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_138),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_9),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_65),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_178),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_128),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_114),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_131),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_129),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_161),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_136),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_110),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_65),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_15),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_163),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_119),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_198),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_193),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_122),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_199),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_174),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_191),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_204),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_202),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_38),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_26),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_34),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_39),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_92),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_79),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_73),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_58),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_69),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_19),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_160),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_23),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_166),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_92),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_1),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_108),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_42),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_48),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_16),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_90),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_95),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_8),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_87),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_45),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_20),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_190),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_221),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_99),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_159),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_186),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_69),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_97),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_54),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_126),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_14),
.Y(n_299)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_187),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_85),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_16),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_40),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_68),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_172),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_225),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_39),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_73),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_142),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_88),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_137),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_11),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_185),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_196),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_71),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_207),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_70),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_75),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_200),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_27),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_31),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_6),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_24),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_28),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_64),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_41),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_24),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_68),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_26),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_100),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_10),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_123),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_61),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_27),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_124),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_169),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_76),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_102),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_145),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_15),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_44),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_51),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_60),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_121),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_55),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_220),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_157),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_175),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_85),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_38),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_150),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_164),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_30),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_152),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_203),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_77),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_227),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_60),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_28),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_107),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_79),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_70),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_153),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_208),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_89),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_33),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_84),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_40),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_95),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_170),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_11),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_12),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_72),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_226),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_149),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_206),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_42),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_120),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_34),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_14),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_72),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_62),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_66),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_213),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_101),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_80),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_52),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_31),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_23),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_57),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_9),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_195),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_94),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_84),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_171),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_61),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_105),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_4),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_74),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_109),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_80),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_21),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_104),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_155),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_168),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_49),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_75),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_43),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_32),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_51),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_141),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_177),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_115),
.Y(n_413)
);

BUFx8_ASAP7_75t_SL g414 ( 
.A(n_112),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_130),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_54),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_93),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_46),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_83),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_4),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_25),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_224),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_81),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_35),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_67),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_6),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_184),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_219),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_94),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_90),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_173),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_89),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_17),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_19),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_211),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_20),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_77),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_44),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_229),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_96),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_53),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_0),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_55),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_1),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_63),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_88),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_63),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_0),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_58),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_151),
.Y(n_450)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_154),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_234),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_377),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_326),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_414),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_326),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_326),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_240),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_243),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_326),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_326),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_250),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_347),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_293),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_326),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_244),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_356),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_431),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_327),
.B(n_2),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_253),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_356),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_344),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_356),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_255),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_356),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_356),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_378),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_356),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_378),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_417),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_417),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_417),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_258),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_259),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_417),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_417),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_417),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_260),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_304),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_319),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_451),
.Y(n_491)
);

INVxp33_ASAP7_75t_SL g492 ( 
.A(n_445),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_304),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_232),
.B(n_2),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_304),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_437),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_263),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_264),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_234),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_235),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_235),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_275),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_277),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_231),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_231),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_L g506 ( 
.A(n_405),
.B(n_3),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_271),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_232),
.B(n_3),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_271),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_283),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_283),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_280),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_290),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_308),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_232),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_236),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_292),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_236),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_294),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_332),
.B(n_5),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_296),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_298),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_309),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_238),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_314),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_238),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_330),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_335),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_308),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_368),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_368),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_344),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_380),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_332),
.B(n_428),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_338),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_380),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

INVxp33_ASAP7_75t_L g538 ( 
.A(n_233),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_339),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_346),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_344),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_438),
.Y(n_542)
);

NOR2xp67_ASAP7_75t_L g543 ( 
.A(n_405),
.B(n_5),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_281),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_351),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_300),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_352),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_281),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_355),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_281),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_310),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_405),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_R g553 ( 
.A(n_405),
.B(n_7),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_428),
.B(n_7),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_357),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_310),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_310),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_323),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_323),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_323),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_386),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_336),
.B(n_8),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_386),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_336),
.B(n_10),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_360),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_374),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_400),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_404),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_386),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_434),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_434),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_411),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_434),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_456),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_456),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_534),
.B(n_412),
.Y(n_576)
);

NOR2x1_ASAP7_75t_L g577 ( 
.A(n_506),
.B(n_239),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_477),
.A2(n_377),
.B1(n_321),
.B2(n_252),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_471),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_471),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_472),
.B(n_266),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_494),
.B(n_370),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_471),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_552),
.B(n_415),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_454),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_453),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_454),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_479),
.A2(n_433),
.B1(n_410),
.B2(n_324),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_457),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_457),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_460),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_460),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_461),
.Y(n_593)
);

INVx6_ASAP7_75t_L g594 ( 
.A(n_541),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_515),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_461),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_494),
.B(n_239),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_465),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_465),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_467),
.Y(n_600)
);

NOR2x1_ASAP7_75t_L g601 ( 
.A(n_543),
.B(n_245),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_467),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_473),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_508),
.B(n_370),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_473),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_475),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_SL g607 ( 
.A(n_469),
.B(n_341),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_490),
.B(n_300),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_475),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_550),
.B(n_422),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_550),
.B(n_427),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_476),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_476),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_496),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_478),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_458),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_492),
.A2(n_362),
.B1(n_302),
.B2(n_233),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_478),
.Y(n_618)
);

AND2x6_ASAP7_75t_L g619 ( 
.A(n_508),
.B(n_370),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_550),
.B(n_532),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_SL g621 ( 
.A(n_491),
.B(n_341),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_480),
.Y(n_622)
);

AND2x6_ASAP7_75t_L g623 ( 
.A(n_480),
.B(n_370),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_481),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_548),
.B(n_439),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_481),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_548),
.B(n_230),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_482),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_482),
.Y(n_629)
);

AND2x2_ASAP7_75t_SL g630 ( 
.A(n_562),
.B(n_370),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_462),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_515),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_485),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_485),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_486),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_486),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_459),
.B(n_247),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_487),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_573),
.B(n_520),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_487),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_464),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_504),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_489),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_573),
.B(n_254),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_504),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_466),
.B(n_470),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_489),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_452),
.B(n_245),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_493),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_493),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_495),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_495),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_505),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_505),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_507),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_468),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_499),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_554),
.B(n_348),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_500),
.B(n_246),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_501),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_507),
.Y(n_661)
);

INVx5_ASAP7_75t_L g662 ( 
.A(n_541),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_509),
.Y(n_663)
);

CKINVDCx8_ASAP7_75t_R g664 ( 
.A(n_455),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_509),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_544),
.B(n_266),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_544),
.B(n_325),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_510),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_607),
.B(n_474),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_658),
.B(n_483),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_616),
.B(n_325),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_658),
.B(n_484),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_637),
.B(n_488),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_580),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_574),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_585),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_585),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_632),
.B(n_546),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_574),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_574),
.Y(n_680)
);

BUFx10_ASAP7_75t_L g681 ( 
.A(n_646),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_594),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_597),
.B(n_551),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_607),
.B(n_498),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_631),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_584),
.B(n_502),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_595),
.B(n_512),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_645),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_645),
.Y(n_689)
);

BUFx2_ASAP7_75t_L g690 ( 
.A(n_632),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_645),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_589),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_584),
.B(n_513),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_L g694 ( 
.A(n_620),
.B(n_553),
.C(n_463),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_645),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_589),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_SL g697 ( 
.A(n_617),
.B(n_497),
.Y(n_697)
);

AO21x2_ASAP7_75t_L g698 ( 
.A1(n_620),
.A2(n_611),
.B(n_610),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_576),
.B(n_517),
.Y(n_699)
);

INVx4_ASAP7_75t_L g700 ( 
.A(n_662),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_610),
.B(n_523),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_611),
.B(n_576),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_639),
.B(n_527),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_645),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_591),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_645),
.Y(n_706)
);

AND2x6_ASAP7_75t_L g707 ( 
.A(n_597),
.B(n_370),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_630),
.A2(n_564),
.B1(n_518),
.B2(n_524),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_650),
.Y(n_709)
);

CKINVDCx16_ASAP7_75t_R g710 ( 
.A(n_621),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_591),
.Y(n_711)
);

OR2x6_ASAP7_75t_L g712 ( 
.A(n_608),
.B(n_546),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_639),
.B(n_535),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_631),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_598),
.Y(n_715)
);

INVx5_ASAP7_75t_L g716 ( 
.A(n_582),
.Y(n_716)
);

BUFx10_ASAP7_75t_L g717 ( 
.A(n_586),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_625),
.B(n_545),
.Y(n_718)
);

NAND3xp33_ASAP7_75t_L g719 ( 
.A(n_627),
.B(n_566),
.C(n_549),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_594),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_650),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_598),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_594),
.B(n_503),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_630),
.A2(n_526),
.B1(n_516),
.B2(n_242),
.Y(n_724)
);

AND3x2_ASAP7_75t_L g725 ( 
.A(n_621),
.B(n_441),
.C(n_248),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_581),
.B(n_551),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_650),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_625),
.B(n_556),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_650),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_599),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_627),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_580),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_594),
.B(n_519),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_599),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_594),
.B(n_556),
.Y(n_735)
);

AND2x2_ASAP7_75t_SL g736 ( 
.A(n_630),
.B(n_246),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_597),
.B(n_581),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_600),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_600),
.Y(n_739)
);

OAI21xp33_ASAP7_75t_SL g740 ( 
.A1(n_577),
.A2(n_249),
.B(n_248),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_644),
.B(n_521),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_602),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_650),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_602),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_644),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_650),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_587),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_580),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_587),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_597),
.B(n_572),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_587),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_582),
.A2(n_242),
.B1(n_265),
.B2(n_237),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_641),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_582),
.A2(n_265),
.B1(n_268),
.B2(n_237),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_580),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_582),
.B(n_557),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_590),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_580),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_609),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_656),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_590),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_609),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_582),
.A2(n_273),
.B1(n_276),
.B2(n_268),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_662),
.B(n_522),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_662),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_582),
.B(n_557),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_615),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_615),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_578),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_580),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_662),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_666),
.B(n_525),
.Y(n_772)
);

INVx5_ASAP7_75t_L g773 ( 
.A(n_582),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_662),
.B(n_528),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_622),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_662),
.B(n_539),
.Y(n_776)
);

INVx5_ASAP7_75t_L g777 ( 
.A(n_582),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_662),
.B(n_540),
.Y(n_778)
);

INVx5_ASAP7_75t_L g779 ( 
.A(n_604),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_622),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_SL g781 ( 
.A(n_664),
.B(n_547),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_583),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_590),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_628),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_583),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_614),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_666),
.B(n_571),
.Y(n_787)
);

AND3x2_ASAP7_75t_L g788 ( 
.A(n_614),
.B(n_256),
.C(n_249),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_628),
.Y(n_789)
);

AND2x6_ASAP7_75t_L g790 ( 
.A(n_577),
.B(n_375),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_633),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_604),
.B(n_558),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_664),
.B(n_555),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_604),
.B(n_558),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_667),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_667),
.B(n_565),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_617),
.A2(n_568),
.B1(n_567),
.B2(n_251),
.Y(n_797)
);

NAND3xp33_ASAP7_75t_L g798 ( 
.A(n_601),
.B(n_560),
.C(n_559),
.Y(n_798)
);

INVxp33_ASAP7_75t_SL g799 ( 
.A(n_588),
.Y(n_799)
);

NAND3xp33_ASAP7_75t_L g800 ( 
.A(n_601),
.B(n_659),
.C(n_648),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_633),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_592),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_648),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_634),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_648),
.B(n_559),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_634),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_635),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_656),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_604),
.B(n_560),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_635),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_657),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_648),
.B(n_538),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_657),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_657),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_659),
.B(n_571),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_592),
.Y(n_816)
);

AND3x1_ASAP7_75t_L g817 ( 
.A(n_588),
.B(n_276),
.C(n_273),
.Y(n_817)
);

INVxp67_ASAP7_75t_SL g818 ( 
.A(n_583),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_659),
.B(n_561),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_664),
.B(n_300),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_578),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_592),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_606),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_659),
.B(n_300),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_604),
.B(n_561),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_654),
.B(n_563),
.Y(n_826)
);

AND2x6_ASAP7_75t_L g827 ( 
.A(n_593),
.B(n_375),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_657),
.B(n_563),
.Y(n_828)
);

AND2x2_ASAP7_75t_SL g829 ( 
.A(n_583),
.B(n_375),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_826),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_676),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_736),
.B(n_375),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_826),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_736),
.B(n_375),
.Y(n_834)
);

BUFx8_ASAP7_75t_L g835 ( 
.A(n_786),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_702),
.B(n_375),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_670),
.A2(n_619),
.B1(n_604),
.B2(n_256),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_735),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_703),
.B(n_604),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_713),
.B(n_604),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_803),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_672),
.B(n_619),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_673),
.B(n_619),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_803),
.Y(n_844)
);

NAND3xp33_ASAP7_75t_L g845 ( 
.A(n_694),
.B(n_267),
.C(n_241),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_731),
.B(n_569),
.Y(n_846)
);

AOI221xp5_ASAP7_75t_L g847 ( 
.A1(n_817),
.A2(n_350),
.B1(n_343),
.B2(n_342),
.C(n_337),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_731),
.B(n_619),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_683),
.Y(n_849)
);

BUFx6f_ASAP7_75t_SL g850 ( 
.A(n_717),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_745),
.B(n_619),
.Y(n_851)
);

BUFx6f_ASAP7_75t_SL g852 ( 
.A(n_717),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_675),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_745),
.B(n_619),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_683),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_737),
.B(n_619),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_741),
.B(n_657),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_795),
.A2(n_619),
.B1(n_261),
.B2(n_262),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_724),
.B(n_657),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_683),
.B(n_569),
.Y(n_860)
);

BUFx10_ASAP7_75t_L g861 ( 
.A(n_725),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_678),
.Y(n_862)
);

CKINVDCx11_ASAP7_75t_R g863 ( 
.A(n_760),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_674),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_674),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_716),
.B(n_660),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_676),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_678),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_690),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_686),
.B(n_660),
.Y(n_870)
);

NAND2xp33_ASAP7_75t_SL g871 ( 
.A(n_820),
.B(n_269),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_674),
.Y(n_872)
);

INVxp67_ASAP7_75t_SL g873 ( 
.A(n_674),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_693),
.B(n_660),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_675),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_795),
.B(n_570),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_679),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_677),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_728),
.B(n_660),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_679),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_690),
.B(n_570),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_680),
.Y(n_882)
);

OR2x6_ASAP7_75t_L g883 ( 
.A(n_786),
.B(n_279),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_718),
.B(n_660),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_701),
.B(n_660),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_772),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_719),
.B(n_270),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_680),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_698),
.A2(n_282),
.B1(n_288),
.B2(n_279),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_685),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_698),
.A2(n_288),
.B1(n_295),
.B2(n_282),
.Y(n_891)
);

NAND3xp33_ASAP7_75t_L g892 ( 
.A(n_796),
.B(n_274),
.C(n_272),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_812),
.B(n_583),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_677),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_732),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_747),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_716),
.B(n_773),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_708),
.B(n_583),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_698),
.B(n_593),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_819),
.B(n_593),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_716),
.B(n_257),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_805),
.B(n_593),
.Y(n_902)
);

NAND3xp33_ASAP7_75t_L g903 ( 
.A(n_769),
.B(n_684),
.C(n_669),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_800),
.A2(n_261),
.B1(n_262),
.B2(n_257),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_805),
.B(n_596),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_699),
.B(n_687),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_787),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_692),
.Y(n_908)
);

NOR2xp67_ASAP7_75t_L g909 ( 
.A(n_798),
.B(n_651),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_750),
.B(n_278),
.Y(n_910)
);

INVx8_ASAP7_75t_L g911 ( 
.A(n_671),
.Y(n_911)
);

NAND3xp33_ASAP7_75t_SL g912 ( 
.A(n_797),
.B(n_821),
.C(n_808),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_716),
.B(n_291),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_818),
.A2(n_579),
.B(n_606),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_815),
.B(n_596),
.Y(n_915)
);

NAND3xp33_ASAP7_75t_L g916 ( 
.A(n_726),
.B(n_285),
.C(n_284),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_815),
.B(n_596),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_674),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_723),
.B(n_286),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_726),
.A2(n_305),
.B1(n_306),
.B2(n_291),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_716),
.B(n_305),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_692),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_696),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_696),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_753),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_717),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_733),
.B(n_287),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_714),
.B(n_289),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_824),
.A2(n_311),
.B1(n_313),
.B2(n_306),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_829),
.A2(n_313),
.B1(n_316),
.B2(n_311),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_716),
.B(n_316),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_773),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_787),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_705),
.B(n_297),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_705),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_711),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_711),
.B(n_299),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_788),
.Y(n_938)
);

NAND3xp33_ASAP7_75t_L g939 ( 
.A(n_697),
.B(n_315),
.C(n_303),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_773),
.B(n_354),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_773),
.B(n_354),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_773),
.B(n_777),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_682),
.B(n_654),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_747),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_715),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_715),
.B(n_317),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_SL g947 ( 
.A(n_781),
.B(n_363),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_722),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_722),
.B(n_596),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_730),
.B(n_624),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_808),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_730),
.B(n_734),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_734),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_773),
.B(n_364),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_738),
.B(n_739),
.Y(n_955)
);

OR2x6_ASAP7_75t_L g956 ( 
.A(n_793),
.B(n_295),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_777),
.B(n_364),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_738),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_671),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_739),
.B(n_624),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_681),
.B(n_663),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_742),
.B(n_318),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_742),
.B(n_624),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_744),
.B(n_624),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_744),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_777),
.B(n_376),
.Y(n_966)
);

INVxp67_ASAP7_75t_SL g967 ( 
.A(n_755),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_777),
.B(n_376),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_777),
.B(n_384),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_759),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_749),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_759),
.B(n_626),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_762),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_749),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_671),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_762),
.B(n_626),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_767),
.B(n_626),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_753),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_707),
.Y(n_979)
);

OR2x6_ASAP7_75t_L g980 ( 
.A(n_712),
.B(n_301),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_767),
.B(n_626),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_751),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_681),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_751),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_768),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_777),
.B(n_384),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_755),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_768),
.B(n_320),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_764),
.A2(n_385),
.B1(n_395),
.B2(n_392),
.Y(n_989)
);

BUFx6f_ASAP7_75t_SL g990 ( 
.A(n_681),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_775),
.B(n_322),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_775),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_779),
.B(n_385),
.Y(n_993)
);

BUFx8_ASAP7_75t_L g994 ( 
.A(n_799),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_757),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_780),
.B(n_603),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_780),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_757),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_682),
.B(n_663),
.Y(n_999)
);

BUFx4f_ASAP7_75t_L g1000 ( 
.A(n_712),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_784),
.B(n_789),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_710),
.B(n_665),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_784),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_829),
.A2(n_397),
.B1(n_392),
.B2(n_395),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_789),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_885),
.A2(n_720),
.B(n_779),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_864),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_857),
.B(n_829),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_831),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_831),
.Y(n_1010)
);

OAI21xp33_ASAP7_75t_L g1011 ( 
.A1(n_947),
.A2(n_799),
.B(n_712),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_890),
.B(n_710),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_857),
.B(n_791),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_906),
.B(n_779),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_890),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_919),
.B(n_791),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_874),
.A2(n_720),
.B(n_779),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_893),
.A2(n_932),
.B(n_879),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_932),
.A2(n_779),
.B(n_766),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_906),
.B(n_779),
.Y(n_1020)
);

NOR2x2_ASAP7_75t_L g1021 ( 
.A(n_980),
.B(n_712),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_867),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_899),
.A2(n_792),
.B(n_756),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_884),
.A2(n_809),
.B(n_794),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_943),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_832),
.A2(n_825),
.B(n_776),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_886),
.B(n_868),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_919),
.B(n_801),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_832),
.A2(n_740),
.B(n_804),
.C(n_801),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_884),
.A2(n_765),
.B(n_700),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_870),
.A2(n_765),
.B(n_700),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_1002),
.B(n_671),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_903),
.A2(n_754),
.B1(n_763),
.B2(n_752),
.Y(n_1033)
);

BUFx3_ASAP7_75t_L g1034 ( 
.A(n_925),
.Y(n_1034)
);

AOI21x1_ASAP7_75t_L g1035 ( 
.A1(n_866),
.A2(n_813),
.B(n_811),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_927),
.B(n_804),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_870),
.A2(n_765),
.B(n_700),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_856),
.A2(n_778),
.B(n_774),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_889),
.A2(n_891),
.B1(n_898),
.B2(n_839),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_961),
.B(n_927),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_897),
.A2(n_771),
.B(n_758),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_834),
.A2(n_807),
.B(n_810),
.C(n_806),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_889),
.A2(n_807),
.B1(n_810),
.B2(n_806),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_881),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_878),
.B(n_828),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_897),
.A2(n_771),
.B(n_758),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_979),
.B(n_811),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_942),
.A2(n_758),
.B(n_755),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_942),
.A2(n_758),
.B(n_755),
.Y(n_1049)
);

INVxp67_ASAP7_75t_L g1050 ( 
.A(n_928),
.Y(n_1050)
);

OAI321xp33_ASAP7_75t_L g1051 ( 
.A1(n_847),
.A2(n_449),
.A3(n_393),
.B1(n_389),
.B2(n_381),
.C(n_448),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_908),
.B(n_732),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_912),
.B(n_813),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_902),
.A2(n_758),
.B(n_755),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_923),
.B(n_732),
.Y(n_1055)
);

OAI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_830),
.A2(n_403),
.B1(n_413),
.B2(n_397),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_905),
.A2(n_782),
.B(n_814),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_915),
.A2(n_782),
.B(n_814),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_979),
.B(n_840),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_935),
.B(n_748),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_917),
.A2(n_967),
.B(n_873),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_834),
.A2(n_413),
.B(n_435),
.C(n_403),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_936),
.B(n_945),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_859),
.A2(n_782),
.B(n_689),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_891),
.A2(n_440),
.B1(n_450),
.B2(n_435),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_948),
.B(n_953),
.Y(n_1066)
);

NAND2x1p5_ASAP7_75t_L g1067 ( 
.A(n_979),
.B(n_748),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_894),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_869),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_864),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_842),
.A2(n_782),
.B(n_689),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_843),
.A2(n_782),
.B(n_691),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_864),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_846),
.B(n_341),
.Y(n_1074)
);

BUFx4f_ASAP7_75t_L g1075 ( 
.A(n_911),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_836),
.A2(n_691),
.B(n_688),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_907),
.B(n_341),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_979),
.B(n_748),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_900),
.A2(n_695),
.B(n_688),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_933),
.B(n_665),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_958),
.B(n_770),
.Y(n_1081)
);

AOI21x1_ASAP7_75t_L g1082 ( 
.A1(n_866),
.A2(n_704),
.B(n_695),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_838),
.A2(n_706),
.B(n_704),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_862),
.Y(n_1084)
);

NOR3xp33_ASAP7_75t_L g1085 ( 
.A(n_939),
.B(n_450),
.C(n_440),
.Y(n_1085)
);

AO21x1_ASAP7_75t_L g1086 ( 
.A1(n_930),
.A2(n_1004),
.B(n_836),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_848),
.A2(n_783),
.B(n_802),
.C(n_761),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_970),
.B(n_770),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_851),
.A2(n_854),
.B(n_952),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_876),
.B(n_510),
.Y(n_1090)
);

INVx1_ASAP7_75t_SL g1091 ( 
.A(n_863),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_849),
.A2(n_706),
.B1(n_785),
.B2(n_770),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_949),
.A2(n_721),
.B(n_709),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_910),
.A2(n_785),
.B(n_721),
.C(n_727),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_922),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_950),
.A2(n_727),
.B(n_709),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_955),
.A2(n_743),
.B(n_729),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_960),
.A2(n_743),
.B(n_729),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_1000),
.B(n_746),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_833),
.A2(n_761),
.B(n_823),
.C(n_822),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_910),
.A2(n_785),
.B(n_746),
.C(n_822),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_951),
.B(n_328),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_860),
.B(n_883),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_943),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_864),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_973),
.B(n_707),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_999),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_887),
.A2(n_783),
.B(n_823),
.C(n_816),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_985),
.B(n_707),
.Y(n_1109)
);

INVx3_ASAP7_75t_SL g1110 ( 
.A(n_978),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_860),
.B(n_511),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1001),
.A2(n_816),
.B(n_802),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_992),
.B(n_707),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_883),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_883),
.B(n_511),
.Y(n_1115)
);

BUFx8_ASAP7_75t_L g1116 ( 
.A(n_850),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_922),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_924),
.A2(n_707),
.B1(n_790),
.B2(n_342),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_855),
.A2(n_358),
.B1(n_353),
.B2(n_349),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_887),
.A2(n_337),
.B(n_350),
.C(n_343),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_997),
.B(n_707),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_1000),
.B(n_363),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_865),
.A2(n_579),
.B(n_606),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_845),
.B(n_329),
.Y(n_1124)
);

AND2x2_ASAP7_75t_SL g1125 ( 
.A(n_989),
.B(n_301),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_865),
.A2(n_579),
.B(n_612),
.Y(n_1126)
);

AOI21x1_ASAP7_75t_L g1127 ( 
.A1(n_914),
.A2(n_613),
.B(n_612),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_1003),
.A2(n_312),
.B(n_407),
.C(n_421),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_965),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_965),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1005),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_853),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_865),
.A2(n_613),
.B(n_612),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_904),
.A2(n_312),
.B(n_307),
.C(n_367),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_956),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_SL g1136 ( 
.A(n_983),
.B(n_333),
.C(n_331),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_841),
.B(n_363),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_875),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_956),
.Y(n_1139)
);

INVx4_ASAP7_75t_L g1140 ( 
.A(n_865),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_SL g1141 ( 
.A(n_850),
.B(n_852),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_872),
.A2(n_618),
.B(n_613),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_872),
.A2(n_636),
.B(n_618),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_872),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_872),
.A2(n_636),
.B(n_618),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_844),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_918),
.A2(n_987),
.B(n_996),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_934),
.B(n_707),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_963),
.A2(n_790),
.B(n_827),
.Y(n_1149)
);

NOR3xp33_ASAP7_75t_L g1150 ( 
.A(n_892),
.B(n_340),
.C(n_334),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_959),
.B(n_307),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_877),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_934),
.B(n_514),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_999),
.B(n_918),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_937),
.B(n_790),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_918),
.A2(n_638),
.B(n_636),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_929),
.A2(n_425),
.B1(n_359),
.B2(n_361),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_918),
.A2(n_640),
.B(n_638),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_987),
.B(n_363),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_880),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_835),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_956),
.A2(n_790),
.B1(n_402),
.B2(n_367),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_895),
.A2(n_429),
.B1(n_365),
.B2(n_366),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_964),
.A2(n_790),
.B(n_827),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_987),
.A2(n_640),
.B(n_638),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_916),
.B(n_345),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_896),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_987),
.A2(n_640),
.B(n_605),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_909),
.A2(n_790),
.B1(n_827),
.B2(n_651),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_972),
.A2(n_605),
.B(n_603),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_976),
.A2(n_605),
.B(n_603),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_937),
.B(n_514),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_977),
.A2(n_652),
.B(n_647),
.Y(n_1173)
);

OAI21xp33_ASAP7_75t_L g1174 ( 
.A1(n_946),
.A2(n_371),
.B(n_369),
.Y(n_1174)
);

NOR2xp67_ASAP7_75t_L g1175 ( 
.A(n_946),
.B(n_98),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_895),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_981),
.A2(n_790),
.B(n_827),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_920),
.A2(n_406),
.B1(n_373),
.B2(n_381),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_901),
.A2(n_605),
.B(n_603),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_901),
.A2(n_605),
.B(n_603),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_962),
.B(n_529),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_962),
.A2(n_398),
.B(n_393),
.C(n_389),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_988),
.B(n_652),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_988),
.B(n_653),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_944),
.A2(n_407),
.B1(n_373),
.B2(n_398),
.Y(n_1185)
);

AND2x2_ASAP7_75t_SL g1186 ( 
.A(n_837),
.B(n_399),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_861),
.B(n_858),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_861),
.B(n_575),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_991),
.B(n_372),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_991),
.B(n_653),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_913),
.A2(n_605),
.B(n_603),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_971),
.B(n_653),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_913),
.A2(n_629),
.B(n_643),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_871),
.A2(n_827),
.B1(n_623),
.B2(n_661),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_974),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_975),
.A2(n_827),
.B1(n_623),
.B2(n_661),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_980),
.B(n_379),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1025),
.B(n_926),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_SL g1199 ( 
.A1(n_1059),
.A2(n_966),
.B(n_921),
.C(n_993),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1015),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1153),
.B(n_982),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1009),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1022),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_1015),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1189),
.A2(n_911),
.B(n_995),
.C(n_998),
.Y(n_1205)
);

BUFx12f_ASAP7_75t_L g1206 ( 
.A(n_1116),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1027),
.B(n_980),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1172),
.B(n_984),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1016),
.A2(n_926),
.B1(n_990),
.B2(n_911),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1065),
.A2(n_442),
.B1(n_399),
.B2(n_402),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1018),
.A2(n_931),
.B(n_921),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1181),
.B(n_882),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1040),
.B(n_888),
.Y(n_1213)
);

OAI21xp33_ASAP7_75t_L g1214 ( 
.A1(n_1189),
.A2(n_938),
.B(n_383),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1124),
.A2(n_954),
.B(n_993),
.C(n_931),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1068),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1025),
.B(n_835),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1028),
.B(n_940),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1036),
.B(n_940),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1008),
.A2(n_990),
.B1(n_968),
.B2(n_986),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1027),
.B(n_852),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_1069),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1007),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1069),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1039),
.A2(n_954),
.B(n_941),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_1104),
.B(n_941),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1012),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1124),
.A2(n_957),
.B(n_986),
.C(n_969),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1074),
.B(n_529),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1007),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1056),
.A2(n_449),
.B(n_406),
.C(n_418),
.Y(n_1231)
);

INVx1_ASAP7_75t_SL g1232 ( 
.A(n_1110),
.Y(n_1232)
);

BUFx4f_ASAP7_75t_SL g1233 ( 
.A(n_1110),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1010),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1034),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1007),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1090),
.B(n_957),
.Y(n_1237)
);

OAI21xp33_ASAP7_75t_L g1238 ( 
.A1(n_1174),
.A2(n_387),
.B(n_382),
.Y(n_1238)
);

AO32x1_ASAP7_75t_L g1239 ( 
.A1(n_1043),
.A2(n_448),
.A3(n_421),
.B1(n_442),
.B2(n_444),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1044),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1104),
.A2(n_966),
.B1(n_969),
.B2(n_968),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1103),
.Y(n_1242)
);

OA22x2_ASAP7_75t_L g1243 ( 
.A1(n_1011),
.A2(n_418),
.B1(n_444),
.B2(n_388),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1130),
.Y(n_1244)
);

NAND3xp33_ASAP7_75t_SL g1245 ( 
.A(n_1182),
.B(n_443),
.C(n_391),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1135),
.Y(n_1246)
);

INVxp67_ASAP7_75t_L g1247 ( 
.A(n_1053),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1107),
.B(n_994),
.Y(n_1248)
);

OR2x6_ASAP7_75t_L g1249 ( 
.A(n_1161),
.B(n_994),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1023),
.A2(n_629),
.B(n_649),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1050),
.B(n_390),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1032),
.A2(n_642),
.B1(n_827),
.B2(n_661),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1183),
.B(n_642),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1024),
.A2(n_629),
.B(n_649),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1186),
.A2(n_446),
.B1(n_396),
.B2(n_401),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1095),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1116),
.Y(n_1257)
);

BUFx4f_ASAP7_75t_L g1258 ( 
.A(n_1114),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1107),
.B(n_1013),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1032),
.B(n_394),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1117),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1063),
.B(n_655),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1111),
.B(n_530),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1066),
.B(n_408),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1131),
.B(n_655),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1080),
.B(n_409),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1080),
.B(n_1146),
.Y(n_1267)
);

NOR2x1_ASAP7_75t_L g1268 ( 
.A(n_1136),
.B(n_655),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1075),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1175),
.B(n_1084),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1129),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1053),
.B(n_1045),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1139),
.B(n_416),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1007),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1186),
.A2(n_419),
.B1(n_420),
.B2(n_423),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1089),
.A2(n_629),
.B(n_649),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1184),
.B(n_668),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1038),
.A2(n_629),
.B(n_647),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1190),
.B(n_668),
.Y(n_1279)
);

OAI21xp33_ASAP7_75t_L g1280 ( 
.A1(n_1102),
.A2(n_424),
.B(n_426),
.Y(n_1280)
);

AOI22x1_ASAP7_75t_L g1281 ( 
.A1(n_1097),
.A2(n_668),
.B1(n_647),
.B2(n_643),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1155),
.A2(n_430),
.B1(n_432),
.B2(n_436),
.Y(n_1282)
);

NAND2x1p5_ASAP7_75t_L g1283 ( 
.A(n_1140),
.B(n_575),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1132),
.Y(n_1284)
);

OR2x6_ASAP7_75t_L g1285 ( 
.A(n_1154),
.B(n_530),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1077),
.B(n_531),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1056),
.A2(n_542),
.B(n_537),
.C(n_536),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_R g1288 ( 
.A(n_1075),
.B(n_447),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_SL g1289 ( 
.A1(n_1059),
.A2(n_542),
.B(n_537),
.C(n_536),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1167),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1166),
.B(n_531),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_1115),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1166),
.A2(n_533),
.B(n_643),
.C(n_575),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1102),
.B(n_575),
.Y(n_1294)
);

BUFx12f_ASAP7_75t_L g1295 ( 
.A(n_1151),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_1151),
.B(n_533),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_1091),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1061),
.A2(n_629),
.B(n_575),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1070),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1138),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1152),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1187),
.B(n_13),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1197),
.B(n_13),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1187),
.B(n_18),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1014),
.A2(n_575),
.B(n_623),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1160),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1125),
.B(n_623),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1021),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1125),
.B(n_623),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1052),
.Y(n_1310)
);

NAND3xp33_ASAP7_75t_L g1311 ( 
.A(n_1150),
.B(n_1197),
.C(n_1085),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1055),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1148),
.A2(n_111),
.B1(n_223),
.B2(n_222),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1150),
.A2(n_623),
.B1(n_103),
.B2(n_106),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1070),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_1141),
.Y(n_1316)
);

O2A1O1Ixp5_ASAP7_75t_L g1317 ( 
.A1(n_1086),
.A2(n_623),
.B(n_218),
.C(n_216),
.Y(n_1317)
);

NOR2xp67_ASAP7_75t_L g1318 ( 
.A(n_1122),
.B(n_113),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1176),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1060),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1154),
.A2(n_215),
.B1(n_214),
.B2(n_212),
.Y(n_1321)
);

NOR3xp33_ASAP7_75t_SL g1322 ( 
.A(n_1051),
.B(n_18),
.C(n_21),
.Y(n_1322)
);

BUFx4f_ASAP7_75t_L g1323 ( 
.A(n_1070),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1029),
.A2(n_1026),
.B(n_1042),
.C(n_1062),
.Y(n_1324)
);

OAI22x1_ASAP7_75t_L g1325 ( 
.A1(n_1122),
.A2(n_22),
.B1(n_29),
.B2(n_30),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1014),
.A2(n_1020),
.B1(n_1176),
.B2(n_1162),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1162),
.B(n_116),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1020),
.A2(n_623),
.B(n_210),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1137),
.B(n_22),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1006),
.A2(n_209),
.B(n_205),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1017),
.A2(n_201),
.B(n_197),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1030),
.A2(n_1037),
.B(n_1031),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1081),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1195),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1054),
.A2(n_192),
.B(n_188),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1163),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1070),
.Y(n_1337)
);

AO32x1_ASAP7_75t_L g1338 ( 
.A1(n_1092),
.A2(n_29),
.A3(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1147),
.A2(n_183),
.B(n_182),
.Y(n_1339)
);

NOR3xp33_ASAP7_75t_SL g1340 ( 
.A(n_1137),
.B(n_36),
.C(n_37),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1195),
.Y(n_1341)
);

OAI22x1_ASAP7_75t_L g1342 ( 
.A1(n_1159),
.A2(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1188),
.B(n_43),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1073),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1085),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1188),
.B(n_47),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1088),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1195),
.Y(n_1348)
);

NOR2xp67_ASAP7_75t_L g1349 ( 
.A(n_1159),
.B(n_181),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1072),
.A2(n_176),
.B(n_167),
.Y(n_1350)
);

O2A1O1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1120),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_SL g1352 ( 
.A(n_1073),
.B(n_165),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1033),
.B(n_50),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1157),
.A2(n_52),
.B1(n_53),
.B2(n_56),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_R g1355 ( 
.A(n_1035),
.B(n_162),
.Y(n_1355)
);

O2A1O1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1134),
.A2(n_56),
.B(n_57),
.C(n_59),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_SL g1357 ( 
.A(n_1073),
.B(n_158),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_L g1358 ( 
.A(n_1119),
.B(n_156),
.Y(n_1358)
);

NOR3xp33_ASAP7_75t_L g1359 ( 
.A(n_1128),
.B(n_1099),
.C(n_1121),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1118),
.A2(n_148),
.B1(n_147),
.B2(n_146),
.Y(n_1360)
);

OAI22x1_ASAP7_75t_L g1361 ( 
.A1(n_1099),
.A2(n_59),
.B1(n_62),
.B2(n_64),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1195),
.B(n_1106),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1071),
.A2(n_144),
.B(n_143),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1178),
.A2(n_66),
.B1(n_67),
.B2(n_71),
.Y(n_1364)
);

AOI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1311),
.A2(n_1260),
.B1(n_1207),
.B2(n_1336),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1272),
.A2(n_1108),
.B(n_1064),
.Y(n_1366)
);

AOI221xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1302),
.A2(n_1178),
.B1(n_1185),
.B2(n_1100),
.C(n_1101),
.Y(n_1367)
);

CKINVDCx9p33_ASAP7_75t_R g1368 ( 
.A(n_1221),
.Y(n_1368)
);

O2A1O1Ixp33_ASAP7_75t_L g1369 ( 
.A1(n_1353),
.A2(n_1094),
.B(n_1087),
.C(n_1113),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_SL g1370 ( 
.A1(n_1205),
.A2(n_1109),
.B(n_1047),
.C(n_1177),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1332),
.A2(n_1276),
.B(n_1254),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1202),
.Y(n_1372)
);

O2A1O1Ixp5_ASAP7_75t_L g1373 ( 
.A1(n_1317),
.A2(n_1173),
.B(n_1093),
.C(n_1096),
.Y(n_1373)
);

AO21x2_ASAP7_75t_L g1374 ( 
.A1(n_1324),
.A2(n_1098),
.B(n_1076),
.Y(n_1374)
);

BUFx3_ASAP7_75t_L g1375 ( 
.A(n_1233),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1269),
.B(n_1140),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_SL g1377 ( 
.A(n_1222),
.B(n_1105),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1211),
.A2(n_1079),
.B(n_1112),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1247),
.B(n_1185),
.Y(n_1379)
);

AND3x1_ASAP7_75t_SL g1380 ( 
.A(n_1354),
.B(n_74),
.C(n_76),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1277),
.A2(n_1057),
.B(n_1058),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1223),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1302),
.A2(n_1118),
.B1(n_1047),
.B2(n_1164),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1279),
.A2(n_1208),
.B(n_1201),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1278),
.A2(n_1298),
.B(n_1082),
.Y(n_1385)
);

BUFx10_ASAP7_75t_L g1386 ( 
.A(n_1221),
.Y(n_1386)
);

AOI221x1_ASAP7_75t_L g1387 ( 
.A1(n_1361),
.A2(n_1083),
.B1(n_1170),
.B2(n_1171),
.C(n_1145),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1304),
.A2(n_1149),
.B1(n_1192),
.B2(n_1073),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1212),
.A2(n_1049),
.B(n_1048),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1304),
.A2(n_1169),
.B(n_1194),
.C(n_1196),
.Y(n_1390)
);

O2A1O1Ixp5_ASAP7_75t_SL g1391 ( 
.A1(n_1291),
.A2(n_1247),
.B(n_1270),
.C(n_1220),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1227),
.B(n_1105),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1294),
.A2(n_1019),
.B(n_1144),
.Y(n_1393)
);

AO31x2_ASAP7_75t_L g1394 ( 
.A1(n_1293),
.A2(n_1143),
.A3(n_1156),
.B(n_1158),
.Y(n_1394)
);

O2A1O1Ixp5_ASAP7_75t_L g1395 ( 
.A1(n_1317),
.A2(n_1225),
.B(n_1326),
.C(n_1350),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1207),
.B(n_1105),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1323),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1233),
.Y(n_1398)
);

A2O1A1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1260),
.A2(n_1193),
.B(n_1126),
.C(n_1123),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1214),
.A2(n_1041),
.B(n_1046),
.C(n_1133),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1218),
.A2(n_1165),
.B(n_1142),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1292),
.A2(n_1144),
.B1(n_1105),
.B2(n_1179),
.Y(n_1402)
);

AOI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1292),
.A2(n_1144),
.B1(n_1180),
.B2(n_1191),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1258),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1234),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1245),
.A2(n_1144),
.B1(n_1078),
.B2(n_1067),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1323),
.Y(n_1407)
);

BUFx2_ASAP7_75t_R g1408 ( 
.A(n_1257),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1223),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1250),
.A2(n_1127),
.B(n_1168),
.Y(n_1410)
);

AOI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1259),
.A2(n_1219),
.B(n_1253),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1329),
.A2(n_1078),
.B(n_1067),
.C(n_82),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1256),
.Y(n_1413)
);

AOI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1262),
.A2(n_117),
.B(n_139),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1229),
.B(n_78),
.Y(n_1415)
);

AO31x2_ASAP7_75t_L g1416 ( 
.A1(n_1342),
.A2(n_78),
.A3(n_81),
.B(n_82),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1224),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1286),
.B(n_83),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1215),
.A2(n_1228),
.B(n_1199),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1237),
.A2(n_125),
.B(n_135),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1263),
.B(n_86),
.Y(n_1421)
);

NOR2x1_ASAP7_75t_L g1422 ( 
.A(n_1315),
.B(n_118),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1362),
.A2(n_127),
.B(n_132),
.Y(n_1423)
);

NAND3x1_ASAP7_75t_L g1424 ( 
.A(n_1303),
.B(n_87),
.C(n_91),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1258),
.Y(n_1425)
);

OAI22x1_ASAP7_75t_L g1426 ( 
.A1(n_1329),
.A2(n_91),
.B1(n_93),
.B2(n_140),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1359),
.A2(n_1213),
.B(n_1312),
.Y(n_1427)
);

OAI22x1_ASAP7_75t_L g1428 ( 
.A1(n_1217),
.A2(n_1308),
.B1(n_1200),
.B2(n_1242),
.Y(n_1428)
);

OR2x6_ASAP7_75t_L g1429 ( 
.A(n_1249),
.B(n_1248),
.Y(n_1429)
);

O2A1O1Ixp33_ASAP7_75t_SL g1430 ( 
.A1(n_1327),
.A2(n_1357),
.B(n_1352),
.C(n_1343),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_SL g1431 ( 
.A1(n_1360),
.A2(n_1313),
.B(n_1321),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1310),
.A2(n_1320),
.B(n_1347),
.Y(n_1432)
);

INVx4_ASAP7_75t_L g1433 ( 
.A(n_1223),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1267),
.A2(n_1333),
.B1(n_1271),
.B2(n_1261),
.Y(n_1434)
);

INVxp67_ASAP7_75t_L g1435 ( 
.A(n_1200),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1281),
.A2(n_1305),
.B(n_1363),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1267),
.A2(n_1290),
.B1(n_1364),
.B2(n_1306),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_SL g1438 ( 
.A(n_1232),
.B(n_1206),
.Y(n_1438)
);

AOI221x1_ASAP7_75t_L g1439 ( 
.A1(n_1325),
.A2(n_1359),
.B1(n_1245),
.B2(n_1345),
.C(n_1335),
.Y(n_1439)
);

O2A1O1Ixp33_ASAP7_75t_SL g1440 ( 
.A1(n_1346),
.A2(n_1309),
.B(n_1307),
.C(n_1264),
.Y(n_1440)
);

O2A1O1Ixp5_ASAP7_75t_L g1441 ( 
.A1(n_1339),
.A2(n_1330),
.B(n_1331),
.C(n_1328),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1224),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1358),
.A2(n_1280),
.B(n_1318),
.C(n_1238),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1241),
.A2(n_1265),
.B(n_1349),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_SL g1445 ( 
.A1(n_1198),
.A2(n_1351),
.B(n_1356),
.C(n_1231),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1203),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_SL g1447 ( 
.A1(n_1266),
.A2(n_1314),
.B(n_1341),
.C(n_1348),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1216),
.A2(n_1244),
.B(n_1252),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1284),
.Y(n_1449)
);

NOR4xp25_ASAP7_75t_L g1450 ( 
.A(n_1364),
.B(n_1255),
.C(n_1275),
.D(n_1210),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1300),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1283),
.A2(n_1226),
.B(n_1334),
.Y(n_1452)
);

NOR4xp25_ASAP7_75t_L g1453 ( 
.A(n_1255),
.B(n_1275),
.C(n_1210),
.D(n_1282),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1285),
.A2(n_1226),
.B(n_1239),
.Y(n_1454)
);

INVxp67_ASAP7_75t_SL g1455 ( 
.A(n_1223),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1285),
.A2(n_1239),
.B(n_1268),
.Y(n_1456)
);

AO31x2_ASAP7_75t_L g1457 ( 
.A1(n_1239),
.A2(n_1319),
.A3(n_1209),
.B(n_1273),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1301),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1285),
.A2(n_1289),
.B(n_1338),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1296),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1338),
.A2(n_1283),
.B(n_1230),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1296),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1242),
.B(n_1251),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1204),
.B(n_1246),
.Y(n_1464)
);

CKINVDCx11_ASAP7_75t_R g1465 ( 
.A(n_1249),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1230),
.A2(n_1274),
.B(n_1236),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1251),
.B(n_1243),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1344),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1299),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1204),
.B(n_1240),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1243),
.B(n_1322),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1338),
.A2(n_1230),
.B(n_1274),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1299),
.A2(n_1337),
.B(n_1287),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1240),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1337),
.A2(n_1355),
.B(n_1273),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1230),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1236),
.A2(n_1274),
.B(n_1322),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1354),
.B(n_1340),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1235),
.B(n_1340),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1297),
.Y(n_1480)
);

O2A1O1Ixp33_ASAP7_75t_SL g1481 ( 
.A1(n_1316),
.A2(n_1236),
.B(n_1274),
.C(n_1288),
.Y(n_1481)
);

NAND2xp33_ASAP7_75t_L g1482 ( 
.A(n_1236),
.B(n_1295),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1249),
.A2(n_1332),
.B(n_1013),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1269),
.B(n_1267),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1256),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1272),
.A2(n_1247),
.B1(n_1189),
.B2(n_1016),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1332),
.A2(n_1276),
.B(n_1254),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1272),
.B(n_1247),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1247),
.B(n_886),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1311),
.A2(n_1189),
.B1(n_886),
.B2(n_464),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1332),
.A2(n_1013),
.B(n_874),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1332),
.A2(n_1013),
.B(n_874),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1272),
.B(n_1247),
.Y(n_1493)
);

AO31x2_ASAP7_75t_L g1494 ( 
.A1(n_1324),
.A2(n_1086),
.A3(n_1039),
.B(n_1205),
.Y(n_1494)
);

O2A1O1Ixp33_ASAP7_75t_SL g1495 ( 
.A1(n_1353),
.A2(n_834),
.B(n_832),
.C(n_1205),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1332),
.A2(n_1013),
.B(n_874),
.Y(n_1496)
);

AO22x2_ASAP7_75t_L g1497 ( 
.A1(n_1311),
.A2(n_1353),
.B1(n_1245),
.B2(n_1122),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1332),
.A2(n_1013),
.B(n_874),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1323),
.Y(n_1499)
);

A2O1A1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1311),
.A2(n_1189),
.B(n_906),
.C(n_672),
.Y(n_1500)
);

AO31x2_ASAP7_75t_L g1501 ( 
.A1(n_1324),
.A2(n_1086),
.A3(n_1039),
.B(n_1205),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1224),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1332),
.A2(n_1276),
.B(n_1254),
.Y(n_1503)
);

AOI221x1_ASAP7_75t_L g1504 ( 
.A1(n_1353),
.A2(n_1189),
.B1(n_1311),
.B2(n_1361),
.C(n_1325),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1332),
.A2(n_1276),
.B(n_1254),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1332),
.A2(n_1013),
.B(n_874),
.Y(n_1506)
);

AOI221xp5_ASAP7_75t_SL g1507 ( 
.A1(n_1302),
.A2(n_1189),
.B1(n_1304),
.B2(n_1247),
.C(n_1011),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1233),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1224),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_SL g1510 ( 
.A(n_1222),
.B(n_886),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1233),
.Y(n_1511)
);

O2A1O1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1353),
.A2(n_1189),
.B(n_1304),
.C(n_1302),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1332),
.A2(n_1013),
.B(n_874),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1256),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1311),
.A2(n_1189),
.B1(n_886),
.B2(n_464),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1272),
.B(n_1247),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1332),
.A2(n_1013),
.B(n_874),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1332),
.A2(n_1276),
.B(n_1254),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1332),
.A2(n_1013),
.B(n_874),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1332),
.A2(n_1276),
.B(n_1254),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1332),
.A2(n_1276),
.B(n_1254),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1272),
.A2(n_1189),
.B(n_1040),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1332),
.A2(n_1013),
.B(n_874),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1272),
.B(n_1247),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1272),
.B(n_1247),
.Y(n_1525)
);

O2A1O1Ixp33_ASAP7_75t_SL g1526 ( 
.A1(n_1353),
.A2(n_834),
.B(n_832),
.C(n_1205),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1272),
.B(n_1247),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1202),
.Y(n_1528)
);

A2O1A1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1311),
.A2(n_1189),
.B(n_906),
.C(n_672),
.Y(n_1529)
);

AOI221xp5_ASAP7_75t_SL g1530 ( 
.A1(n_1302),
.A2(n_1189),
.B1(n_1304),
.B2(n_1247),
.C(n_1011),
.Y(n_1530)
);

OR2x6_ASAP7_75t_SL g1531 ( 
.A(n_1336),
.B(n_983),
.Y(n_1531)
);

A2O1A1Ixp33_ASAP7_75t_L g1532 ( 
.A1(n_1311),
.A2(n_1189),
.B(n_906),
.C(n_672),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1224),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1272),
.A2(n_1247),
.B1(n_1189),
.B2(n_1016),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1272),
.B(n_1247),
.Y(n_1535)
);

A2O1A1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1311),
.A2(n_1189),
.B(n_906),
.C(n_672),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1256),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1272),
.B(n_1247),
.Y(n_1538)
);

INVx3_ASAP7_75t_L g1539 ( 
.A(n_1223),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1223),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1478),
.A2(n_1486),
.B1(n_1534),
.B2(n_1365),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1372),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1405),
.Y(n_1543)
);

OAI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1490),
.A2(n_1515),
.B1(n_1471),
.B2(n_1493),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1413),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_SL g1546 ( 
.A1(n_1467),
.A2(n_1497),
.B1(n_1450),
.B2(n_1522),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1375),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1497),
.A2(n_1479),
.B1(n_1463),
.B2(n_1489),
.Y(n_1548)
);

BUFx12f_ASAP7_75t_L g1549 ( 
.A(n_1465),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1500),
.A2(n_1529),
.B1(n_1532),
.B2(n_1536),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1512),
.A2(n_1527),
.B1(n_1538),
.B2(n_1516),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1512),
.A2(n_1488),
.B1(n_1524),
.B2(n_1525),
.Y(n_1552)
);

INVx6_ASAP7_75t_L g1553 ( 
.A(n_1397),
.Y(n_1553)
);

CKINVDCx6p67_ASAP7_75t_R g1554 ( 
.A(n_1398),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1426),
.A2(n_1497),
.B1(n_1535),
.B2(n_1379),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_1480),
.Y(n_1556)
);

INVx6_ASAP7_75t_L g1557 ( 
.A(n_1397),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1417),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1418),
.A2(n_1415),
.B1(n_1419),
.B2(n_1427),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1380),
.A2(n_1419),
.B1(n_1424),
.B2(n_1453),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1392),
.B(n_1468),
.Y(n_1561)
);

INVx4_ASAP7_75t_L g1562 ( 
.A(n_1407),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1407),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_SL g1564 ( 
.A1(n_1421),
.A2(n_1437),
.B1(n_1429),
.B2(n_1386),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_SL g1565 ( 
.A1(n_1429),
.A2(n_1386),
.B1(n_1438),
.B2(n_1530),
.Y(n_1565)
);

CKINVDCx11_ASAP7_75t_R g1566 ( 
.A(n_1531),
.Y(n_1566)
);

BUFx12f_ASAP7_75t_L g1567 ( 
.A(n_1484),
.Y(n_1567)
);

CKINVDCx11_ASAP7_75t_R g1568 ( 
.A(n_1511),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1396),
.A2(n_1383),
.B1(n_1510),
.B2(n_1509),
.Y(n_1569)
);

BUFx12f_ASAP7_75t_L g1570 ( 
.A(n_1484),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1408),
.Y(n_1571)
);

INVx6_ASAP7_75t_L g1572 ( 
.A(n_1499),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1528),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1388),
.A2(n_1431),
.B1(n_1464),
.B2(n_1462),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1442),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1485),
.Y(n_1576)
);

AOI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1507),
.A2(n_1429),
.B1(n_1428),
.B2(n_1460),
.Y(n_1577)
);

INVx8_ASAP7_75t_L g1578 ( 
.A(n_1499),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1499),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1368),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1434),
.A2(n_1482),
.B1(n_1404),
.B2(n_1425),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1502),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1483),
.A2(n_1432),
.B1(n_1474),
.B2(n_1533),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1432),
.A2(n_1411),
.B1(n_1537),
.B2(n_1514),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1376),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1451),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1435),
.A2(n_1443),
.B1(n_1470),
.B2(n_1390),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1430),
.A2(n_1412),
.B1(n_1367),
.B2(n_1422),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1446),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1435),
.A2(n_1445),
.B1(n_1458),
.B2(n_1449),
.Y(n_1590)
);

CKINVDCx11_ASAP7_75t_R g1591 ( 
.A(n_1433),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1469),
.Y(n_1592)
);

INVxp67_ASAP7_75t_SL g1593 ( 
.A(n_1411),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1374),
.A2(n_1423),
.B1(n_1420),
.B2(n_1477),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1406),
.A2(n_1402),
.B1(n_1377),
.B2(n_1483),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1384),
.A2(n_1420),
.B1(n_1374),
.B2(n_1423),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1476),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1382),
.Y(n_1598)
);

INVxp67_ASAP7_75t_SL g1599 ( 
.A(n_1455),
.Y(n_1599)
);

INVx6_ASAP7_75t_L g1600 ( 
.A(n_1481),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1448),
.Y(n_1601)
);

BUFx2_ASAP7_75t_SL g1602 ( 
.A(n_1409),
.Y(n_1602)
);

OAI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1504),
.A2(n_1439),
.B1(n_1384),
.B2(n_1403),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1448),
.Y(n_1604)
);

BUFx2_ASAP7_75t_SL g1605 ( 
.A(n_1409),
.Y(n_1605)
);

CKINVDCx16_ASAP7_75t_R g1606 ( 
.A(n_1366),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1444),
.A2(n_1456),
.B1(n_1454),
.B2(n_1459),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1444),
.A2(n_1455),
.B1(n_1454),
.B2(n_1456),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1400),
.A2(n_1399),
.B1(n_1540),
.B2(n_1539),
.Y(n_1609)
);

CKINVDCx11_ASAP7_75t_R g1610 ( 
.A(n_1391),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1540),
.Y(n_1611)
);

CKINVDCx11_ASAP7_75t_R g1612 ( 
.A(n_1466),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1459),
.A2(n_1475),
.B1(n_1401),
.B2(n_1496),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1416),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1491),
.A2(n_1498),
.B1(n_1523),
.B2(n_1496),
.Y(n_1615)
);

OAI21xp33_ASAP7_75t_L g1616 ( 
.A1(n_1389),
.A2(n_1369),
.B(n_1523),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1416),
.Y(n_1617)
);

INVx6_ASAP7_75t_L g1618 ( 
.A(n_1447),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1452),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_SL g1620 ( 
.A1(n_1472),
.A2(n_1461),
.B1(n_1416),
.B2(n_1494),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1461),
.A2(n_1389),
.B1(n_1472),
.B2(n_1381),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1393),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1416),
.A2(n_1494),
.B1(n_1501),
.B2(n_1395),
.Y(n_1623)
);

CKINVDCx20_ASAP7_75t_R g1624 ( 
.A(n_1393),
.Y(n_1624)
);

OAI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1387),
.A2(n_1491),
.B1(n_1519),
.B2(n_1517),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1494),
.A2(n_1501),
.B1(n_1395),
.B2(n_1498),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1457),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1369),
.A2(n_1506),
.B1(n_1519),
.B2(n_1517),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1492),
.A2(n_1513),
.B1(n_1506),
.B2(n_1381),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1473),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1492),
.A2(n_1513),
.B1(n_1378),
.B2(n_1521),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1378),
.A2(n_1505),
.B1(n_1371),
.B2(n_1520),
.Y(n_1632)
);

CKINVDCx20_ASAP7_75t_R g1633 ( 
.A(n_1440),
.Y(n_1633)
);

BUFx4_ASAP7_75t_R g1634 ( 
.A(n_1457),
.Y(n_1634)
);

OAI22xp33_ASAP7_75t_SL g1635 ( 
.A1(n_1414),
.A2(n_1526),
.B1(n_1495),
.B2(n_1501),
.Y(n_1635)
);

INVx4_ASAP7_75t_L g1636 ( 
.A(n_1457),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1494),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1487),
.A2(n_1518),
.B1(n_1503),
.B2(n_1410),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1501),
.A2(n_1370),
.B1(n_1441),
.B2(n_1373),
.Y(n_1639)
);

BUFx12f_ASAP7_75t_L g1640 ( 
.A(n_1441),
.Y(n_1640)
);

BUFx2_ASAP7_75t_SL g1641 ( 
.A(n_1394),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_SL g1642 ( 
.A1(n_1373),
.A2(n_1436),
.B1(n_1394),
.B2(n_1385),
.Y(n_1642)
);

OAI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1478),
.A2(n_1365),
.B1(n_947),
.B2(n_1490),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1365),
.A2(n_1189),
.B1(n_1311),
.B2(n_947),
.Y(n_1644)
);

CKINVDCx6p67_ASAP7_75t_R g1645 ( 
.A(n_1375),
.Y(n_1645)
);

OAI22x1_ASAP7_75t_L g1646 ( 
.A1(n_1365),
.A2(n_1515),
.B1(n_1490),
.B2(n_1302),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1480),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1478),
.A2(n_1354),
.B1(n_1189),
.B2(n_1304),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1375),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1478),
.A2(n_1354),
.B1(n_1189),
.B2(n_1304),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1480),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1365),
.A2(n_1490),
.B1(n_1515),
.B2(n_710),
.Y(n_1652)
);

AOI21xp33_ASAP7_75t_L g1653 ( 
.A1(n_1512),
.A2(n_1189),
.B(n_1500),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1365),
.A2(n_1490),
.B1(n_1515),
.B2(n_710),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1486),
.B(n_1272),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1375),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1480),
.Y(n_1657)
);

BUFx2_ASAP7_75t_SL g1658 ( 
.A(n_1375),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1372),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1478),
.A2(n_1354),
.B1(n_1189),
.B2(n_1304),
.Y(n_1660)
);

INVx1_ASAP7_75t_SL g1661 ( 
.A(n_1480),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1478),
.A2(n_1354),
.B1(n_1189),
.B2(n_1304),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1478),
.A2(n_1354),
.B1(n_1189),
.B2(n_1304),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1365),
.A2(n_1490),
.B1(n_1515),
.B2(n_710),
.Y(n_1664)
);

CKINVDCx11_ASAP7_75t_R g1665 ( 
.A(n_1465),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1490),
.A2(n_1189),
.B1(n_1515),
.B2(n_1365),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1442),
.Y(n_1667)
);

INVx2_ASAP7_75t_SL g1668 ( 
.A(n_1375),
.Y(n_1668)
);

OAI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1500),
.A2(n_1532),
.B(n_1529),
.Y(n_1669)
);

CKINVDCx11_ASAP7_75t_R g1670 ( 
.A(n_1465),
.Y(n_1670)
);

CKINVDCx6p67_ASAP7_75t_R g1671 ( 
.A(n_1375),
.Y(n_1671)
);

INVx4_ASAP7_75t_L g1672 ( 
.A(n_1397),
.Y(n_1672)
);

CKINVDCx11_ASAP7_75t_R g1673 ( 
.A(n_1465),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1480),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1372),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1365),
.A2(n_1189),
.B1(n_1311),
.B2(n_947),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1480),
.Y(n_1677)
);

INVx6_ASAP7_75t_L g1678 ( 
.A(n_1397),
.Y(n_1678)
);

INVx6_ASAP7_75t_L g1679 ( 
.A(n_1397),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1413),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_SL g1681 ( 
.A1(n_1478),
.A2(n_710),
.B1(n_621),
.B2(n_947),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1413),
.Y(n_1682)
);

OAI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1478),
.A2(n_1365),
.B1(n_947),
.B2(n_1490),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1486),
.B(n_1272),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1365),
.A2(n_1490),
.B1(n_1515),
.B2(n_710),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1480),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_SL g1687 ( 
.A1(n_1478),
.A2(n_710),
.B1(n_621),
.B2(n_947),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1372),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1372),
.Y(n_1689)
);

CKINVDCx6p67_ASAP7_75t_R g1690 ( 
.A(n_1375),
.Y(n_1690)
);

CKINVDCx16_ASAP7_75t_R g1691 ( 
.A(n_1375),
.Y(n_1691)
);

CKINVDCx14_ASAP7_75t_R g1692 ( 
.A(n_1508),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1372),
.Y(n_1693)
);

INVx6_ASAP7_75t_L g1694 ( 
.A(n_1397),
.Y(n_1694)
);

BUFx2_ASAP7_75t_L g1695 ( 
.A(n_1442),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1372),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1397),
.Y(n_1697)
);

BUFx12f_ASAP7_75t_L g1698 ( 
.A(n_1465),
.Y(n_1698)
);

BUFx3_ASAP7_75t_L g1699 ( 
.A(n_1375),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1413),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1372),
.Y(n_1701)
);

BUFx3_ASAP7_75t_L g1702 ( 
.A(n_1375),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1365),
.A2(n_1189),
.B1(n_1311),
.B2(n_947),
.Y(n_1703)
);

INVx3_ASAP7_75t_SL g1704 ( 
.A(n_1508),
.Y(n_1704)
);

CKINVDCx11_ASAP7_75t_R g1705 ( 
.A(n_1465),
.Y(n_1705)
);

BUFx2_ASAP7_75t_SL g1706 ( 
.A(n_1375),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1372),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_1480),
.Y(n_1708)
);

OAI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1478),
.A2(n_1365),
.B1(n_947),
.B2(n_1490),
.Y(n_1709)
);

CKINVDCx20_ASAP7_75t_R g1710 ( 
.A(n_1480),
.Y(n_1710)
);

OAI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1478),
.A2(n_1365),
.B1(n_947),
.B2(n_1490),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1397),
.Y(n_1712)
);

BUFx3_ASAP7_75t_L g1713 ( 
.A(n_1375),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1480),
.Y(n_1714)
);

OAI21x1_ASAP7_75t_L g1715 ( 
.A1(n_1629),
.A2(n_1638),
.B(n_1631),
.Y(n_1715)
);

AO21x2_ASAP7_75t_L g1716 ( 
.A1(n_1653),
.A2(n_1625),
.B(n_1603),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1601),
.Y(n_1717)
);

OR2x6_ASAP7_75t_L g1718 ( 
.A(n_1641),
.B(n_1640),
.Y(n_1718)
);

BUFx2_ASAP7_75t_L g1719 ( 
.A(n_1622),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1666),
.A2(n_1650),
.B1(n_1660),
.B2(n_1648),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1604),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1637),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1614),
.Y(n_1723)
);

BUFx4f_ASAP7_75t_SL g1724 ( 
.A(n_1556),
.Y(n_1724)
);

INVx4_ASAP7_75t_L g1725 ( 
.A(n_1612),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1619),
.B(n_1624),
.Y(n_1726)
);

INVx1_ASAP7_75t_SL g1727 ( 
.A(n_1558),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1617),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1652),
.A2(n_1664),
.B1(n_1654),
.B2(n_1685),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_1619),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1593),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1606),
.B(n_1627),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1542),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1667),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1543),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1593),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1630),
.B(n_1669),
.Y(n_1737)
);

NOR2x1_ASAP7_75t_SL g1738 ( 
.A(n_1595),
.B(n_1550),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1630),
.Y(n_1739)
);

INVx3_ASAP7_75t_L g1740 ( 
.A(n_1630),
.Y(n_1740)
);

BUFx3_ASAP7_75t_L g1741 ( 
.A(n_1600),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1577),
.B(n_1599),
.Y(n_1742)
);

OA21x2_ASAP7_75t_L g1743 ( 
.A1(n_1607),
.A2(n_1621),
.B(n_1616),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1548),
.B(n_1607),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1600),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1546),
.B(n_1623),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1608),
.Y(n_1747)
);

AO21x2_ASAP7_75t_L g1748 ( 
.A1(n_1625),
.A2(n_1603),
.B(n_1628),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1646),
.A2(n_1676),
.B1(n_1703),
.B2(n_1644),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1551),
.B(n_1552),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1544),
.B(n_1655),
.Y(n_1751)
);

OAI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1648),
.A2(n_1660),
.B(n_1650),
.Y(n_1752)
);

BUFx2_ASAP7_75t_L g1753 ( 
.A(n_1599),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1573),
.Y(n_1754)
);

OAI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1662),
.A2(n_1663),
.B(n_1559),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1695),
.Y(n_1756)
);

OA21x2_ASAP7_75t_L g1757 ( 
.A1(n_1615),
.A2(n_1613),
.B(n_1596),
.Y(n_1757)
);

NAND2x1p5_ASAP7_75t_L g1758 ( 
.A(n_1588),
.B(n_1590),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1659),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1675),
.B(n_1688),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1684),
.B(n_1636),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1689),
.Y(n_1762)
);

CKINVDCx20_ASAP7_75t_R g1763 ( 
.A(n_1710),
.Y(n_1763)
);

OAI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1662),
.A2(n_1663),
.B(n_1559),
.Y(n_1764)
);

BUFx2_ASAP7_75t_L g1765 ( 
.A(n_1633),
.Y(n_1765)
);

OAI21x1_ASAP7_75t_L g1766 ( 
.A1(n_1632),
.A2(n_1615),
.B(n_1613),
.Y(n_1766)
);

AOI211x1_ASAP7_75t_L g1767 ( 
.A1(n_1643),
.A2(n_1683),
.B(n_1711),
.C(n_1709),
.Y(n_1767)
);

INVx3_ASAP7_75t_L g1768 ( 
.A(n_1636),
.Y(n_1768)
);

OAI21x1_ASAP7_75t_L g1769 ( 
.A1(n_1639),
.A2(n_1609),
.B(n_1596),
.Y(n_1769)
);

NAND2x1p5_ASAP7_75t_L g1770 ( 
.A(n_1693),
.B(n_1696),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1701),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1707),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1575),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1555),
.B(n_1541),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1642),
.Y(n_1775)
);

INVxp67_ASAP7_75t_SL g1776 ( 
.A(n_1584),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1620),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1544),
.B(n_1541),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1620),
.Y(n_1779)
);

AO31x2_ASAP7_75t_L g1780 ( 
.A1(n_1587),
.A2(n_1634),
.A3(n_1574),
.B(n_1623),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1589),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1584),
.B(n_1583),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1597),
.B(n_1585),
.Y(n_1783)
);

BUFx3_ASAP7_75t_L g1784 ( 
.A(n_1582),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1546),
.B(n_1555),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1626),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1626),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1618),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1709),
.B(n_1561),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1576),
.Y(n_1790)
);

OR2x6_ASAP7_75t_L g1791 ( 
.A(n_1618),
.B(n_1569),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1618),
.Y(n_1792)
);

OAI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1681),
.A2(n_1687),
.B1(n_1560),
.B2(n_1581),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1635),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1647),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1586),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1545),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1560),
.B(n_1565),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1681),
.A2(n_1687),
.B1(n_1564),
.B2(n_1565),
.Y(n_1799)
);

OAI21x1_ASAP7_75t_L g1800 ( 
.A1(n_1611),
.A2(n_1592),
.B(n_1700),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1680),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1682),
.B(n_1564),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1594),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1594),
.Y(n_1804)
);

OAI21x1_ASAP7_75t_L g1805 ( 
.A1(n_1579),
.A2(n_1697),
.B(n_1610),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1602),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1598),
.Y(n_1807)
);

OAI21x1_ASAP7_75t_L g1808 ( 
.A1(n_1579),
.A2(n_1697),
.B(n_1605),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1585),
.Y(n_1809)
);

AO21x1_ASAP7_75t_L g1810 ( 
.A1(n_1562),
.A2(n_1672),
.B(n_1591),
.Y(n_1810)
);

BUFx3_ASAP7_75t_L g1811 ( 
.A(n_1567),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1562),
.B(n_1672),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1566),
.A2(n_1549),
.B1(n_1698),
.B2(n_1570),
.Y(n_1813)
);

AO31x2_ASAP7_75t_L g1814 ( 
.A1(n_1580),
.A2(n_1563),
.A3(n_1712),
.B(n_1678),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1712),
.Y(n_1815)
);

OAI21x1_ASAP7_75t_L g1816 ( 
.A1(n_1578),
.A2(n_1572),
.B(n_1553),
.Y(n_1816)
);

OAI21x1_ASAP7_75t_L g1817 ( 
.A1(n_1578),
.A2(n_1572),
.B(n_1553),
.Y(n_1817)
);

BUFx3_ASAP7_75t_L g1818 ( 
.A(n_1557),
.Y(n_1818)
);

CKINVDCx11_ASAP7_75t_R g1819 ( 
.A(n_1665),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1691),
.B(n_1677),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1657),
.B(n_1661),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1679),
.Y(n_1822)
);

OAI21x1_ASAP7_75t_L g1823 ( 
.A1(n_1679),
.A2(n_1694),
.B(n_1658),
.Y(n_1823)
);

CKINVDCx6p67_ASAP7_75t_R g1824 ( 
.A(n_1670),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1651),
.B(n_1714),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1706),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1656),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1668),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1554),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1645),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1671),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1547),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1674),
.B(n_1708),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1649),
.A2(n_1713),
.B(n_1702),
.Y(n_1834)
);

OA21x2_ASAP7_75t_L g1835 ( 
.A1(n_1571),
.A2(n_1686),
.B(n_1690),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1699),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1704),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1568),
.Y(n_1838)
);

OA21x2_ASAP7_75t_L g1839 ( 
.A1(n_1704),
.A2(n_1692),
.B(n_1673),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1705),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_R g1841 ( 
.A(n_1571),
.B(n_925),
.Y(n_1841)
);

OAI21x1_ASAP7_75t_L g1842 ( 
.A1(n_1629),
.A2(n_1378),
.B(n_1371),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1546),
.B(n_1606),
.Y(n_1843)
);

NAND3xp33_ASAP7_75t_L g1844 ( 
.A(n_1749),
.B(n_1751),
.C(n_1778),
.Y(n_1844)
);

O2A1O1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1720),
.A2(n_1752),
.B(n_1793),
.C(n_1764),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1729),
.A2(n_1799),
.B1(n_1719),
.B2(n_1765),
.Y(n_1846)
);

OAI211xp5_ASAP7_75t_L g1847 ( 
.A1(n_1755),
.A2(n_1729),
.B(n_1767),
.C(n_1750),
.Y(n_1847)
);

NOR2x1_ASAP7_75t_L g1848 ( 
.A(n_1725),
.B(n_1719),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1726),
.B(n_1843),
.Y(n_1849)
);

A2O1A1Ixp33_ASAP7_75t_L g1850 ( 
.A1(n_1750),
.A2(n_1769),
.B(n_1798),
.C(n_1774),
.Y(n_1850)
);

AND2x4_ASAP7_75t_SL g1851 ( 
.A(n_1763),
.B(n_1725),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1732),
.B(n_1761),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1789),
.B(n_1791),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1732),
.B(n_1761),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1791),
.B(n_1738),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1758),
.A2(n_1774),
.B(n_1769),
.Y(n_1856)
);

OAI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1791),
.A2(n_1785),
.B(n_1776),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1753),
.B(n_1744),
.Y(n_1858)
);

OAI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1791),
.A2(n_1744),
.B(n_1766),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1734),
.B(n_1756),
.Y(n_1860)
);

NAND2xp33_ASAP7_75t_R g1861 ( 
.A(n_1791),
.B(n_1743),
.Y(n_1861)
);

INVx4_ASAP7_75t_SL g1862 ( 
.A(n_1814),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1753),
.Y(n_1863)
);

OR2x6_ASAP7_75t_L g1864 ( 
.A(n_1718),
.B(n_1742),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1760),
.B(n_1737),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_1795),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_SL g1867 ( 
.A1(n_1738),
.A2(n_1746),
.B1(n_1748),
.B2(n_1782),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1760),
.B(n_1790),
.Y(n_1868)
);

A2O1A1Ixp33_ASAP7_75t_L g1869 ( 
.A1(n_1782),
.A2(n_1804),
.B(n_1803),
.C(n_1747),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1814),
.B(n_1783),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1737),
.B(n_1773),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1733),
.B(n_1735),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1794),
.Y(n_1873)
);

OAI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1715),
.A2(n_1782),
.B(n_1802),
.Y(n_1874)
);

CKINVDCx20_ASAP7_75t_R g1875 ( 
.A(n_1819),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1757),
.A2(n_1743),
.B(n_1716),
.Y(n_1876)
);

A2O1A1Ixp33_ASAP7_75t_L g1877 ( 
.A1(n_1803),
.A2(n_1804),
.B(n_1747),
.C(n_1787),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1733),
.B(n_1735),
.Y(n_1878)
);

A2O1A1Ixp33_ASAP7_75t_L g1879 ( 
.A1(n_1786),
.A2(n_1787),
.B(n_1741),
.C(n_1779),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1757),
.A2(n_1743),
.B(n_1842),
.Y(n_1880)
);

OAI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1834),
.A2(n_1792),
.B(n_1743),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1781),
.Y(n_1882)
);

AO22x2_ASAP7_75t_L g1883 ( 
.A1(n_1767),
.A2(n_1775),
.B1(n_1779),
.B2(n_1777),
.Y(n_1883)
);

OA21x2_ASAP7_75t_L g1884 ( 
.A1(n_1775),
.A2(n_1786),
.B(n_1777),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1757),
.A2(n_1736),
.B(n_1731),
.Y(n_1885)
);

O2A1O1Ixp33_ASAP7_75t_SL g1886 ( 
.A1(n_1792),
.A2(n_1788),
.B(n_1826),
.C(n_1806),
.Y(n_1886)
);

AND2x6_ASAP7_75t_L g1887 ( 
.A(n_1788),
.B(n_1745),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1754),
.B(n_1759),
.Y(n_1888)
);

AO21x2_ASAP7_75t_L g1889 ( 
.A1(n_1731),
.A2(n_1736),
.B(n_1805),
.Y(n_1889)
);

A2O1A1Ixp33_ASAP7_75t_L g1890 ( 
.A1(n_1741),
.A2(n_1788),
.B(n_1745),
.C(n_1765),
.Y(n_1890)
);

OAI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1806),
.A2(n_1805),
.B(n_1823),
.Y(n_1891)
);

NAND3xp33_ASAP7_75t_L g1892 ( 
.A(n_1826),
.B(n_1745),
.C(n_1725),
.Y(n_1892)
);

OA21x2_ASAP7_75t_L g1893 ( 
.A1(n_1723),
.A2(n_1728),
.B(n_1722),
.Y(n_1893)
);

OAI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1823),
.A2(n_1808),
.B(n_1836),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1788),
.B(n_1725),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1814),
.B(n_1762),
.Y(n_1896)
);

NOR2x1p5_ASAP7_75t_L g1897 ( 
.A(n_1824),
.B(n_1840),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1771),
.B(n_1772),
.Y(n_1898)
);

A2O1A1Ixp33_ASAP7_75t_L g1899 ( 
.A1(n_1745),
.A2(n_1780),
.B(n_1757),
.C(n_1817),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1839),
.A2(n_1824),
.B1(n_1840),
.B2(n_1838),
.Y(n_1900)
);

AND2x4_ASAP7_75t_L g1901 ( 
.A(n_1814),
.B(n_1772),
.Y(n_1901)
);

O2A1O1Ixp33_ASAP7_75t_SL g1902 ( 
.A1(n_1829),
.A2(n_1831),
.B(n_1837),
.C(n_1827),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1814),
.B(n_1784),
.Y(n_1903)
);

AOI221xp5_ASAP7_75t_L g1904 ( 
.A1(n_1727),
.A2(n_1827),
.B1(n_1828),
.B2(n_1832),
.C(n_1801),
.Y(n_1904)
);

OAI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1800),
.A2(n_1821),
.B(n_1820),
.Y(n_1905)
);

NOR2x1_ASAP7_75t_SL g1906 ( 
.A(n_1718),
.B(n_1730),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1770),
.B(n_1780),
.Y(n_1907)
);

OAI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1820),
.A2(n_1832),
.B(n_1828),
.Y(n_1908)
);

A2O1A1Ixp33_ASAP7_75t_L g1909 ( 
.A1(n_1780),
.A2(n_1816),
.B(n_1817),
.C(n_1830),
.Y(n_1909)
);

BUFx2_ASAP7_75t_L g1910 ( 
.A(n_1815),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1780),
.B(n_1809),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1852),
.B(n_1728),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1893),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1870),
.B(n_1739),
.Y(n_1914)
);

INVxp67_ASAP7_75t_SL g1915 ( 
.A(n_1863),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1873),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1893),
.Y(n_1917)
);

INVx1_ASAP7_75t_SL g1918 ( 
.A(n_1910),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1884),
.B(n_1717),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1911),
.B(n_1768),
.Y(n_1920)
);

BUFx3_ASAP7_75t_L g1921 ( 
.A(n_1887),
.Y(n_1921)
);

INVx4_ASAP7_75t_L g1922 ( 
.A(n_1887),
.Y(n_1922)
);

HB1xp67_ASAP7_75t_L g1923 ( 
.A(n_1863),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1865),
.B(n_1907),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1882),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1854),
.B(n_1717),
.Y(n_1926)
);

HB1xp67_ASAP7_75t_L g1927 ( 
.A(n_1884),
.Y(n_1927)
);

INVxp67_ASAP7_75t_SL g1928 ( 
.A(n_1885),
.Y(n_1928)
);

INVxp67_ASAP7_75t_SL g1929 ( 
.A(n_1885),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1858),
.B(n_1721),
.Y(n_1930)
);

INVxp67_ASAP7_75t_L g1931 ( 
.A(n_1884),
.Y(n_1931)
);

NOR2x1p5_ASAP7_75t_L g1932 ( 
.A(n_1892),
.B(n_1830),
.Y(n_1932)
);

OAI222xp33_ASAP7_75t_L g1933 ( 
.A1(n_1845),
.A2(n_1718),
.B1(n_1801),
.B2(n_1797),
.C1(n_1796),
.C2(n_1838),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1844),
.A2(n_1839),
.B1(n_1810),
.B2(n_1811),
.Y(n_1934)
);

INVxp67_ASAP7_75t_L g1935 ( 
.A(n_1868),
.Y(n_1935)
);

BUFx3_ASAP7_75t_L g1936 ( 
.A(n_1887),
.Y(n_1936)
);

INVx1_ASAP7_75t_SL g1937 ( 
.A(n_1871),
.Y(n_1937)
);

AND2x4_ASAP7_75t_L g1938 ( 
.A(n_1862),
.B(n_1740),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1860),
.B(n_1835),
.Y(n_1939)
);

OAI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1846),
.A2(n_1839),
.B1(n_1835),
.B2(n_1718),
.Y(n_1940)
);

NOR2x1_ASAP7_75t_L g1941 ( 
.A(n_1881),
.B(n_1718),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1896),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1872),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1878),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1853),
.A2(n_1839),
.B1(n_1810),
.B2(n_1811),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1901),
.Y(n_1946)
);

OAI221xp5_ASAP7_75t_L g1947 ( 
.A1(n_1845),
.A2(n_1813),
.B1(n_1835),
.B2(n_1811),
.C(n_1829),
.Y(n_1947)
);

BUFx2_ASAP7_75t_L g1948 ( 
.A(n_1891),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1898),
.Y(n_1949)
);

BUFx3_ASAP7_75t_L g1950 ( 
.A(n_1887),
.Y(n_1950)
);

BUFx3_ASAP7_75t_L g1951 ( 
.A(n_1921),
.Y(n_1951)
);

AOI22xp33_ASAP7_75t_L g1952 ( 
.A1(n_1947),
.A2(n_1867),
.B1(n_1855),
.B2(n_1856),
.Y(n_1952)
);

OAI211xp5_ASAP7_75t_SL g1953 ( 
.A1(n_1947),
.A2(n_1934),
.B(n_1847),
.C(n_1905),
.Y(n_1953)
);

NOR2x1p5_ASAP7_75t_L g1954 ( 
.A(n_1922),
.B(n_1830),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1939),
.B(n_1900),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1927),
.Y(n_1956)
);

BUFx2_ASAP7_75t_L g1957 ( 
.A(n_1931),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1923),
.B(n_1876),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1923),
.B(n_1888),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1916),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1913),
.Y(n_1961)
);

INVxp67_ASAP7_75t_SL g1962 ( 
.A(n_1931),
.Y(n_1962)
);

INVx2_ASAP7_75t_SL g1963 ( 
.A(n_1914),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1942),
.B(n_1899),
.Y(n_1964)
);

BUFx3_ASAP7_75t_L g1965 ( 
.A(n_1921),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1916),
.Y(n_1966)
);

BUFx3_ASAP7_75t_L g1967 ( 
.A(n_1921),
.Y(n_1967)
);

INVx1_ASAP7_75t_SL g1968 ( 
.A(n_1918),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1942),
.B(n_1899),
.Y(n_1969)
);

AOI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1928),
.A2(n_1929),
.B(n_1880),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1935),
.B(n_1877),
.Y(n_1971)
);

NAND3xp33_ASAP7_75t_SL g1972 ( 
.A(n_1945),
.B(n_1900),
.C(n_1847),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1946),
.B(n_1859),
.Y(n_1973)
);

NOR2xp33_ASAP7_75t_L g1974 ( 
.A(n_1935),
.B(n_1835),
.Y(n_1974)
);

OAI31xp33_ASAP7_75t_L g1975 ( 
.A1(n_1940),
.A2(n_1850),
.A3(n_1879),
.B(n_1869),
.Y(n_1975)
);

AND2x4_ASAP7_75t_L g1976 ( 
.A(n_1938),
.B(n_1903),
.Y(n_1976)
);

INVx5_ASAP7_75t_SL g1977 ( 
.A(n_1938),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1925),
.Y(n_1978)
);

INVx4_ASAP7_75t_L g1979 ( 
.A(n_1922),
.Y(n_1979)
);

NOR2x1_ASAP7_75t_L g1980 ( 
.A(n_1932),
.B(n_1890),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1925),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1919),
.Y(n_1982)
);

NAND2x1_ASAP7_75t_L g1983 ( 
.A(n_1922),
.B(n_1864),
.Y(n_1983)
);

NAND3xp33_ASAP7_75t_L g1984 ( 
.A(n_1948),
.B(n_1867),
.C(n_1904),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1913),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1943),
.B(n_1877),
.Y(n_1986)
);

OAI21x1_ASAP7_75t_SL g1987 ( 
.A1(n_1941),
.A2(n_1906),
.B(n_1857),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1943),
.B(n_1874),
.Y(n_1988)
);

INVx1_ASAP7_75t_SL g1989 ( 
.A(n_1918),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1924),
.B(n_1889),
.Y(n_1990)
);

BUFx2_ASAP7_75t_L g1991 ( 
.A(n_1950),
.Y(n_1991)
);

OAI211xp5_ASAP7_75t_L g1992 ( 
.A1(n_1929),
.A2(n_1850),
.B(n_1879),
.C(n_1869),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1924),
.B(n_1889),
.Y(n_1993)
);

HB1xp67_ASAP7_75t_L g1994 ( 
.A(n_1919),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1938),
.B(n_1894),
.Y(n_1995)
);

OAI21xp33_ASAP7_75t_L g1996 ( 
.A1(n_1941),
.A2(n_1853),
.B(n_1883),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1949),
.B(n_1849),
.Y(n_1997)
);

HB1xp67_ASAP7_75t_L g1998 ( 
.A(n_1915),
.Y(n_1998)
);

AOI221xp5_ASAP7_75t_L g1999 ( 
.A1(n_1948),
.A2(n_1883),
.B1(n_1855),
.B2(n_1908),
.C(n_1902),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1961),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1990),
.B(n_1993),
.Y(n_2001)
);

INVxp67_ASAP7_75t_SL g2002 ( 
.A(n_1962),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1958),
.B(n_1912),
.Y(n_2003)
);

NAND2x1p5_ASAP7_75t_L g2004 ( 
.A(n_1983),
.B(n_1932),
.Y(n_2004)
);

BUFx2_ASAP7_75t_L g2005 ( 
.A(n_1980),
.Y(n_2005)
);

CKINVDCx16_ASAP7_75t_R g2006 ( 
.A(n_1980),
.Y(n_2006)
);

OR2x2_ASAP7_75t_L g2007 ( 
.A(n_1958),
.B(n_1912),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1964),
.B(n_1920),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1964),
.B(n_1937),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1964),
.B(n_1937),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1960),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1960),
.Y(n_2012)
);

NAND2x1p5_ASAP7_75t_L g2013 ( 
.A(n_1983),
.B(n_1936),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1966),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1969),
.B(n_1917),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1966),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1971),
.B(n_1944),
.Y(n_2017)
);

INVx1_ASAP7_75t_SL g2018 ( 
.A(n_1968),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1978),
.Y(n_2019)
);

INVxp33_ASAP7_75t_L g2020 ( 
.A(n_1974),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1978),
.Y(n_2021)
);

NAND2x1p5_ASAP7_75t_L g2022 ( 
.A(n_1979),
.B(n_1936),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1981),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1988),
.B(n_1926),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_1957),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1969),
.B(n_1914),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1961),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1998),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1969),
.B(n_1914),
.Y(n_2029)
);

AND2x4_ASAP7_75t_L g2030 ( 
.A(n_1976),
.B(n_1936),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1971),
.B(n_1986),
.Y(n_2031)
);

HB1xp67_ASAP7_75t_L g2032 ( 
.A(n_1957),
.Y(n_2032)
);

INVx1_ASAP7_75t_SL g2033 ( 
.A(n_1968),
.Y(n_2033)
);

O2A1O1Ixp33_ASAP7_75t_L g2034 ( 
.A1(n_1953),
.A2(n_1933),
.B(n_1902),
.C(n_1890),
.Y(n_2034)
);

INVx2_ASAP7_75t_SL g2035 ( 
.A(n_1954),
.Y(n_2035)
);

AND2x4_ASAP7_75t_L g2036 ( 
.A(n_1976),
.B(n_1950),
.Y(n_2036)
);

OAI21xp5_ASAP7_75t_L g2037 ( 
.A1(n_1984),
.A2(n_1933),
.B(n_1848),
.Y(n_2037)
);

NOR2xp33_ASAP7_75t_L g2038 ( 
.A(n_1955),
.B(n_1875),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_1986),
.B(n_1930),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1985),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1985),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1982),
.B(n_1915),
.Y(n_2042)
);

INVxp67_ASAP7_75t_L g2043 ( 
.A(n_2005),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2011),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2031),
.B(n_1989),
.Y(n_2045)
);

OR2x2_ASAP7_75t_L g2046 ( 
.A(n_2003),
.B(n_1959),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2030),
.B(n_1963),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_2030),
.B(n_2036),
.Y(n_2048)
);

INVx1_ASAP7_75t_SL g2049 ( 
.A(n_2005),
.Y(n_2049)
);

INVxp67_ASAP7_75t_SL g2050 ( 
.A(n_2025),
.Y(n_2050)
);

INVx3_ASAP7_75t_SL g2051 ( 
.A(n_2006),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2011),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_L g2053 ( 
.A(n_2038),
.B(n_1953),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2030),
.B(n_1963),
.Y(n_2054)
);

AOI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_2006),
.A2(n_1972),
.B1(n_1984),
.B2(n_1992),
.Y(n_2055)
);

NAND3xp33_ASAP7_75t_L g2056 ( 
.A(n_2037),
.B(n_1975),
.C(n_1999),
.Y(n_2056)
);

OAI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_2037),
.A2(n_1972),
.B(n_1992),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2012),
.Y(n_2058)
);

NOR2x1_ASAP7_75t_L g2059 ( 
.A(n_2018),
.B(n_1875),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_2000),
.Y(n_2060)
);

NOR2xp67_ASAP7_75t_L g2061 ( 
.A(n_2035),
.B(n_1963),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2012),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2014),
.Y(n_2063)
);

NOR2xp33_ASAP7_75t_R g2064 ( 
.A(n_2035),
.B(n_1724),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2014),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2031),
.B(n_1989),
.Y(n_2066)
);

NAND5xp2_ASAP7_75t_L g2067 ( 
.A(n_2034),
.B(n_1975),
.C(n_1999),
.D(n_1952),
.E(n_1996),
.Y(n_2067)
);

INVx1_ASAP7_75t_SL g2068 ( 
.A(n_2018),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2016),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_2000),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2033),
.B(n_1996),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2003),
.B(n_1959),
.Y(n_2072)
);

AOI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_2030),
.A2(n_1995),
.B1(n_1973),
.B2(n_1883),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2030),
.B(n_1977),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_L g2075 ( 
.A(n_2020),
.B(n_1831),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2016),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2033),
.B(n_1973),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2036),
.B(n_1977),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_2025),
.Y(n_2079)
);

XNOR2x2_ASAP7_75t_L g2080 ( 
.A(n_2034),
.B(n_2009),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_2007),
.B(n_1982),
.Y(n_2081)
);

INVxp67_ASAP7_75t_L g2082 ( 
.A(n_2017),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2032),
.Y(n_2083)
);

AOI21xp5_ASAP7_75t_L g2084 ( 
.A1(n_2017),
.A2(n_1987),
.B(n_1970),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2036),
.B(n_1977),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2039),
.B(n_1973),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2007),
.B(n_1994),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2032),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2019),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2019),
.Y(n_2090)
);

INVxp67_ASAP7_75t_SL g2091 ( 
.A(n_2004),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2039),
.B(n_1997),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2036),
.B(n_1977),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2021),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2021),
.Y(n_2095)
);

HB1xp67_ASAP7_75t_L g2096 ( 
.A(n_2028),
.Y(n_2096)
);

INVx2_ASAP7_75t_SL g2097 ( 
.A(n_2013),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2036),
.B(n_1977),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2023),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2062),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2060),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2062),
.Y(n_2102)
);

OR2x2_ASAP7_75t_L g2103 ( 
.A(n_2083),
.B(n_2002),
.Y(n_2103)
);

OR2x2_ASAP7_75t_L g2104 ( 
.A(n_2088),
.B(n_2002),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2055),
.B(n_2009),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2057),
.B(n_2009),
.Y(n_2106)
);

INVx2_ASAP7_75t_SL g2107 ( 
.A(n_2074),
.Y(n_2107)
);

HB1xp67_ASAP7_75t_L g2108 ( 
.A(n_2079),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2044),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2052),
.Y(n_2110)
);

OAI31xp33_ASAP7_75t_L g2111 ( 
.A1(n_2056),
.A2(n_2067),
.A3(n_2053),
.B(n_2071),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2053),
.B(n_2010),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2051),
.B(n_2048),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2068),
.B(n_2051),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2048),
.B(n_2035),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2058),
.Y(n_2116)
);

INVx1_ASAP7_75t_SL g2117 ( 
.A(n_2059),
.Y(n_2117)
);

OR2x2_ASAP7_75t_L g2118 ( 
.A(n_2092),
.B(n_2024),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_SL g2119 ( 
.A(n_2064),
.B(n_2004),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2074),
.B(n_2004),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2078),
.B(n_2004),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2075),
.B(n_2045),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2063),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2065),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2078),
.B(n_2026),
.Y(n_2125)
);

INVx1_ASAP7_75t_SL g2126 ( 
.A(n_2064),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2069),
.Y(n_2127)
);

INVxp67_ASAP7_75t_SL g2128 ( 
.A(n_2080),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2085),
.B(n_2026),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2076),
.Y(n_2130)
);

NOR2x1_ASAP7_75t_L g2131 ( 
.A(n_2049),
.B(n_1897),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2075),
.B(n_2010),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2066),
.B(n_2010),
.Y(n_2133)
);

OR2x6_ASAP7_75t_L g2134 ( 
.A(n_2043),
.B(n_2022),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2089),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2082),
.B(n_2008),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2060),
.Y(n_2137)
);

INVx2_ASAP7_75t_SL g2138 ( 
.A(n_2085),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2096),
.B(n_2008),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2090),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2113),
.B(n_2061),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_2131),
.B(n_2050),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2113),
.B(n_2117),
.Y(n_2143)
);

AOI221xp5_ASAP7_75t_L g2144 ( 
.A1(n_2128),
.A2(n_2111),
.B1(n_2105),
.B2(n_2106),
.C(n_2112),
.Y(n_2144)
);

INVx2_ASAP7_75t_SL g2145 ( 
.A(n_2115),
.Y(n_2145)
);

AOI21xp33_ASAP7_75t_SL g2146 ( 
.A1(n_2114),
.A2(n_2080),
.B(n_2013),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2131),
.B(n_2093),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2100),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2100),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2102),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2102),
.Y(n_2151)
);

AOI22xp33_ASAP7_75t_SL g2152 ( 
.A1(n_2120),
.A2(n_2091),
.B1(n_2084),
.B2(n_1987),
.Y(n_2152)
);

NAND2xp33_ASAP7_75t_L g2153 ( 
.A(n_2126),
.B(n_1841),
.Y(n_2153)
);

OAI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_2119),
.A2(n_2073),
.B1(n_2022),
.B2(n_2013),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2108),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2122),
.B(n_2008),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2109),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2109),
.Y(n_2158)
);

AOI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_2107),
.A2(n_2098),
.B1(n_2093),
.B2(n_2077),
.Y(n_2159)
);

OAI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_2132),
.A2(n_2022),
.B1(n_2013),
.B2(n_2097),
.Y(n_2160)
);

HB1xp67_ASAP7_75t_L g2161 ( 
.A(n_2103),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2110),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2110),
.Y(n_2163)
);

OR2x2_ASAP7_75t_L g2164 ( 
.A(n_2139),
.B(n_2086),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_2107),
.B(n_2097),
.Y(n_2165)
);

INVxp67_ASAP7_75t_L g2166 ( 
.A(n_2138),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2138),
.B(n_2115),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2116),
.Y(n_2168)
);

AOI22xp5_ASAP7_75t_L g2169 ( 
.A1(n_2120),
.A2(n_2098),
.B1(n_1995),
.B2(n_2047),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2125),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2161),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2141),
.Y(n_2172)
);

NAND2x1p5_ASAP7_75t_L g2173 ( 
.A(n_2142),
.B(n_1830),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2143),
.B(n_2125),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2144),
.B(n_2129),
.Y(n_2175)
);

AOI221xp5_ASAP7_75t_L g2176 ( 
.A1(n_2146),
.A2(n_2140),
.B1(n_2124),
.B2(n_2127),
.C(n_2135),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_2170),
.B(n_2133),
.Y(n_2177)
);

INVxp33_ASAP7_75t_L g2178 ( 
.A(n_2141),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2166),
.B(n_2129),
.Y(n_2179)
);

AOI32xp33_ASAP7_75t_L g2180 ( 
.A1(n_2142),
.A2(n_2121),
.A3(n_2136),
.B1(n_2103),
.B2(n_2104),
.Y(n_2180)
);

OAI21xp5_ASAP7_75t_L g2181 ( 
.A1(n_2142),
.A2(n_2104),
.B(n_2134),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2161),
.Y(n_2182)
);

XNOR2x1_ASAP7_75t_L g2183 ( 
.A(n_2155),
.B(n_2154),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2148),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2170),
.B(n_2118),
.Y(n_2185)
);

AOI22xp33_ASAP7_75t_L g2186 ( 
.A1(n_2152),
.A2(n_2121),
.B1(n_2118),
.B2(n_2134),
.Y(n_2186)
);

INVxp33_ASAP7_75t_L g2187 ( 
.A(n_2147),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_2145),
.B(n_2116),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2149),
.Y(n_2189)
);

AOI221xp5_ASAP7_75t_L g2190 ( 
.A1(n_2167),
.A2(n_2140),
.B1(n_2124),
.B2(n_2135),
.C(n_2123),
.Y(n_2190)
);

O2A1O1Ixp33_ASAP7_75t_L g2191 ( 
.A1(n_2165),
.A2(n_2134),
.B(n_2130),
.C(n_2127),
.Y(n_2191)
);

OAI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_2153),
.A2(n_2134),
.B(n_1970),
.Y(n_2192)
);

OAI32xp33_ASAP7_75t_L g2193 ( 
.A1(n_2147),
.A2(n_2022),
.A3(n_2130),
.B1(n_2123),
.B2(n_2081),
.Y(n_2193)
);

OAI31xp33_ASAP7_75t_L g2194 ( 
.A1(n_2175),
.A2(n_2160),
.A3(n_2145),
.B(n_2165),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2171),
.Y(n_2195)
);

AOI21xp33_ASAP7_75t_L g2196 ( 
.A1(n_2187),
.A2(n_2153),
.B(n_2159),
.Y(n_2196)
);

AOI21xp5_ASAP7_75t_L g2197 ( 
.A1(n_2191),
.A2(n_2134),
.B(n_2156),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2182),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2185),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2188),
.Y(n_2200)
);

OR2x2_ASAP7_75t_L g2201 ( 
.A(n_2174),
.B(n_2164),
.Y(n_2201)
);

A2O1A1Ixp33_ASAP7_75t_L g2202 ( 
.A1(n_2180),
.A2(n_2168),
.B(n_2163),
.C(n_2162),
.Y(n_2202)
);

O2A1O1Ixp5_ASAP7_75t_L g2203 ( 
.A1(n_2181),
.A2(n_2158),
.B(n_2157),
.C(n_2151),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2184),
.Y(n_2204)
);

NAND3xp33_ASAP7_75t_SL g2205 ( 
.A(n_2186),
.B(n_2169),
.C(n_2150),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2189),
.Y(n_2206)
);

OAI211xp5_ASAP7_75t_L g2207 ( 
.A1(n_2176),
.A2(n_2137),
.B(n_2101),
.C(n_2081),
.Y(n_2207)
);

OA21x2_ASAP7_75t_SL g2208 ( 
.A1(n_2178),
.A2(n_2042),
.B(n_1995),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2172),
.B(n_2101),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2199),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2196),
.B(n_2179),
.Y(n_2211)
);

NOR2xp67_ASAP7_75t_SL g2212 ( 
.A(n_2200),
.B(n_2181),
.Y(n_2212)
);

BUFx2_ASAP7_75t_L g2213 ( 
.A(n_2195),
.Y(n_2213)
);

NOR2xp67_ASAP7_75t_L g2214 ( 
.A(n_2207),
.B(n_2192),
.Y(n_2214)
);

HB1xp67_ASAP7_75t_L g2215 ( 
.A(n_2198),
.Y(n_2215)
);

O2A1O1Ixp33_ASAP7_75t_SL g2216 ( 
.A1(n_2202),
.A2(n_2193),
.B(n_2192),
.C(n_2190),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_2201),
.B(n_2183),
.Y(n_2217)
);

NAND4xp25_ASAP7_75t_L g2218 ( 
.A(n_2194),
.B(n_2177),
.C(n_1833),
.D(n_2137),
.Y(n_2218)
);

NAND4xp25_ASAP7_75t_L g2219 ( 
.A(n_2197),
.B(n_1895),
.C(n_1825),
.D(n_2173),
.Y(n_2219)
);

NOR3xp33_ASAP7_75t_L g2220 ( 
.A(n_2205),
.B(n_1866),
.C(n_2173),
.Y(n_2220)
);

XOR2xp5_ASAP7_75t_L g2221 ( 
.A(n_2209),
.B(n_1807),
.Y(n_2221)
);

OAI21xp5_ASAP7_75t_L g2222 ( 
.A1(n_2203),
.A2(n_1962),
.B(n_2087),
.Y(n_2222)
);

AOI221xp5_ASAP7_75t_L g2223 ( 
.A1(n_2216),
.A2(n_2202),
.B1(n_2203),
.B2(n_2204),
.C(n_2206),
.Y(n_2223)
);

AOI221xp5_ASAP7_75t_L g2224 ( 
.A1(n_2212),
.A2(n_2208),
.B1(n_2070),
.B2(n_2095),
.C(n_2094),
.Y(n_2224)
);

OAI221xp5_ASAP7_75t_SL g2225 ( 
.A1(n_2220),
.A2(n_2087),
.B1(n_2054),
.B2(n_2047),
.C(n_2046),
.Y(n_2225)
);

AOI211xp5_ASAP7_75t_SL g2226 ( 
.A1(n_2217),
.A2(n_1895),
.B(n_1886),
.C(n_2054),
.Y(n_2226)
);

AOI211xp5_ASAP7_75t_L g2227 ( 
.A1(n_2214),
.A2(n_1965),
.B(n_1951),
.C(n_1967),
.Y(n_2227)
);

AOI221xp5_ASAP7_75t_L g2228 ( 
.A1(n_2218),
.A2(n_2070),
.B1(n_2099),
.B2(n_2042),
.C(n_2001),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_SL g2229 ( 
.A(n_2222),
.B(n_2046),
.Y(n_2229)
);

O2A1O1Ixp33_ASAP7_75t_L g2230 ( 
.A1(n_2223),
.A2(n_2215),
.B(n_2213),
.C(n_2210),
.Y(n_2230)
);

OAI21xp5_ASAP7_75t_L g2231 ( 
.A1(n_2229),
.A2(n_2211),
.B(n_2222),
.Y(n_2231)
);

OAI21x1_ASAP7_75t_SL g2232 ( 
.A1(n_2224),
.A2(n_2221),
.B(n_2219),
.Y(n_2232)
);

AOI211xp5_ASAP7_75t_L g2233 ( 
.A1(n_2225),
.A2(n_1951),
.B(n_1965),
.C(n_1967),
.Y(n_2233)
);

O2A1O1Ixp33_ASAP7_75t_L g2234 ( 
.A1(n_2227),
.A2(n_2072),
.B(n_1994),
.C(n_2001),
.Y(n_2234)
);

O2A1O1Ixp33_ASAP7_75t_L g2235 ( 
.A1(n_2226),
.A2(n_2072),
.B(n_2001),
.C(n_1886),
.Y(n_2235)
);

OAI221xp5_ASAP7_75t_SL g2236 ( 
.A1(n_2228),
.A2(n_1991),
.B1(n_1967),
.B2(n_1951),
.C(n_1965),
.Y(n_2236)
);

AOI22xp5_ASAP7_75t_L g2237 ( 
.A1(n_2233),
.A2(n_1851),
.B1(n_1991),
.B2(n_1954),
.Y(n_2237)
);

NOR2x1_ASAP7_75t_L g2238 ( 
.A(n_2230),
.B(n_2000),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2231),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2234),
.B(n_2015),
.Y(n_2240)
);

NOR2x1_ASAP7_75t_L g2241 ( 
.A(n_2235),
.B(n_2027),
.Y(n_2241)
);

INVxp67_ASAP7_75t_SL g2242 ( 
.A(n_2236),
.Y(n_2242)
);

NAND3x1_ASAP7_75t_L g2243 ( 
.A(n_2239),
.B(n_2232),
.C(n_2015),
.Y(n_2243)
);

AND4x1_ASAP7_75t_L g2244 ( 
.A(n_2238),
.B(n_1909),
.C(n_2015),
.D(n_2026),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_2242),
.B(n_2029),
.Y(n_2245)
);

XNOR2x1_ASAP7_75t_L g2246 ( 
.A(n_2245),
.B(n_2241),
.Y(n_2246)
);

BUFx2_ASAP7_75t_L g2247 ( 
.A(n_2246),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2247),
.Y(n_2248)
);

OAI21xp5_ASAP7_75t_L g2249 ( 
.A1(n_2247),
.A2(n_2243),
.B(n_2240),
.Y(n_2249)
);

OAI22xp5_ASAP7_75t_L g2250 ( 
.A1(n_2248),
.A2(n_2237),
.B1(n_2244),
.B2(n_2024),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_2249),
.B(n_2029),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2251),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2250),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2252),
.Y(n_2254)
);

AOI22xp33_ASAP7_75t_L g2255 ( 
.A1(n_2254),
.A2(n_2253),
.B1(n_1979),
.B2(n_1956),
.Y(n_2255)
);

AOI22xp5_ASAP7_75t_L g2256 ( 
.A1(n_2255),
.A2(n_2029),
.B1(n_2027),
.B2(n_2041),
.Y(n_2256)
);

OAI221xp5_ASAP7_75t_R g2257 ( 
.A1(n_2256),
.A2(n_1861),
.B1(n_2027),
.B2(n_2040),
.C(n_2041),
.Y(n_2257)
);

AOI211xp5_ASAP7_75t_L g2258 ( 
.A1(n_2257),
.A2(n_1812),
.B(n_1818),
.C(n_1822),
.Y(n_2258)
);


endmodule