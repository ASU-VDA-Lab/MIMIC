module fake_jpeg_20606_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_0),
.B(n_1),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_L g19 ( 
.A1(n_10),
.A2(n_0),
.B(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_2),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_20),
.Y(n_39)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_3),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_40),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_19),
.B1(n_27),
.B2(n_16),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_19),
.B(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_18),
.Y(n_47)
);

OR2x2_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_27),
.B1(n_16),
.B2(n_25),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_27),
.B1(n_32),
.B2(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_62),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_42),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_41),
.B(n_38),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_57),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_61),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_45),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_18),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_45),
.C(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_47),
.B(n_37),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_73),
.B(n_26),
.Y(n_91)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_71),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_77),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_78),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_42),
.B1(n_26),
.B2(n_24),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_42),
.B1(n_17),
.B2(n_14),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_55),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_51),
.C(n_56),
.Y(n_82)
);

NOR4xp25_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_67),
.C(n_74),
.D(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_17),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_86),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_90),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_56),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_41),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_67),
.C(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_92),
.B(n_14),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_89),
.B(n_72),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_104),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_70),
.C(n_69),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_78),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_93),
.Y(n_104)
);

FAx1_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_86),
.CI(n_84),
.CON(n_105),
.SN(n_105)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_107),
.B(n_78),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_88),
.B(n_90),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_103),
.C(n_95),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_111),
.C(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_112),
.B(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_116),
.B(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_105),
.Y(n_124)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_9),
.C(n_12),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_120),
.B(n_118),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_105),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_123),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_122),
.B(n_124),
.Y(n_129)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_13),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_121),
.A2(n_115),
.B1(n_108),
.B2(n_13),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_126),
.A2(n_48),
.A3(n_5),
.B1(n_4),
.B2(n_10),
.C1(n_11),
.C2(n_7),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_3),
.B(n_4),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_127),
.B(n_8),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_131),
.A2(n_132),
.B(n_129),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_126),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_134),
.Y(n_136)
);


endmodule