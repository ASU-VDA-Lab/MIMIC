module real_aes_148_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_798, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_798;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_755;
wire n_656;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_0), .B(n_139), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_1), .A2(n_148), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_2), .B(n_792), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_3), .B(n_139), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_4), .B(n_155), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_5), .B(n_155), .Y(n_218) );
INVx1_ASAP7_75t_L g146 ( .A(n_6), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_7), .B(n_155), .Y(n_193) );
CKINVDCx16_ASAP7_75t_R g792 ( .A(n_8), .Y(n_792) );
NAND2xp33_ASAP7_75t_L g156 ( .A(n_9), .B(n_157), .Y(n_156) );
AND2x2_ASAP7_75t_L g474 ( .A(n_10), .B(n_165), .Y(n_474) );
AND2x2_ASAP7_75t_L g534 ( .A(n_11), .B(n_134), .Y(n_534) );
INVx2_ASAP7_75t_L g136 ( .A(n_12), .Y(n_136) );
AOI221x1_ASAP7_75t_L g234 ( .A1(n_13), .A2(n_24), .B1(n_139), .B2(n_148), .C(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_14), .B(n_155), .Y(n_508) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_15), .Y(n_116) );
NOR3xp33_ASAP7_75t_L g790 ( .A(n_15), .B(n_791), .C(n_793), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_16), .B(n_139), .Y(n_138) );
AO21x2_ASAP7_75t_L g133 ( .A1(n_17), .A2(n_134), .B(n_137), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_18), .B(n_173), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_19), .B(n_155), .Y(n_182) );
AO21x1_ASAP7_75t_L g213 ( .A1(n_20), .A2(n_139), .B(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_21), .B(n_139), .Y(n_539) );
INVx1_ASAP7_75t_L g120 ( .A(n_22), .Y(n_120) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_23), .A2(n_90), .B1(n_139), .B2(n_479), .Y(n_478) );
NAND2x1_ASAP7_75t_L g204 ( .A(n_25), .B(n_155), .Y(n_204) );
NAND2x1_ASAP7_75t_L g192 ( .A(n_26), .B(n_157), .Y(n_192) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_27), .A2(n_87), .B(n_136), .Y(n_135) );
OR2x2_ASAP7_75t_L g160 ( .A(n_27), .B(n_87), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_28), .B(n_157), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_29), .B(n_155), .Y(n_154) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_30), .A2(n_165), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_31), .B(n_157), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_32), .A2(n_148), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_33), .B(n_155), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_34), .A2(n_148), .B(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g145 ( .A(n_35), .B(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g149 ( .A(n_35), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g487 ( .A(n_35), .Y(n_487) );
OR2x6_ASAP7_75t_L g118 ( .A(n_36), .B(n_119), .Y(n_118) );
INVxp67_ASAP7_75t_L g793 ( .A(n_36), .Y(n_793) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_37), .B(n_139), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_38), .B(n_139), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_39), .B(n_155), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_40), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_41), .B(n_157), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_42), .B(n_139), .Y(n_460) );
XNOR2xp5_ASAP7_75t_L g760 ( .A(n_43), .B(n_761), .Y(n_760) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_44), .A2(n_148), .B(n_470), .Y(n_469) );
OAI22xp5_ASAP7_75t_SL g781 ( .A1(n_45), .A2(n_782), .B1(n_783), .B2(n_784), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_45), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_46), .A2(n_148), .B(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_47), .B(n_157), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_48), .B(n_157), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_49), .B(n_139), .Y(n_505) );
INVx1_ASAP7_75t_L g142 ( .A(n_50), .Y(n_142) );
INVx1_ASAP7_75t_L g152 ( .A(n_50), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_51), .B(n_155), .Y(n_472) );
AND2x2_ASAP7_75t_L g494 ( .A(n_52), .B(n_173), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_53), .B(n_157), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_54), .B(n_155), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_55), .B(n_157), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_56), .A2(n_148), .B(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_57), .B(n_139), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_58), .B(n_139), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_59), .A2(n_148), .B(n_513), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_60), .A2(n_100), .B1(n_762), .B2(n_763), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_60), .Y(n_763) );
AO21x1_ASAP7_75t_L g215 ( .A1(n_61), .A2(n_148), .B(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g545 ( .A(n_62), .B(n_174), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_63), .B(n_139), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_64), .B(n_157), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_65), .B(n_139), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_66), .A2(n_79), .B1(n_785), .B2(n_786), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_66), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_67), .B(n_157), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_68), .A2(n_94), .B1(n_148), .B2(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_69), .Y(n_769) );
AND2x2_ASAP7_75t_L g228 ( .A(n_70), .B(n_174), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_71), .B(n_155), .Y(n_542) );
INVx1_ASAP7_75t_L g144 ( .A(n_72), .Y(n_144) );
INVx1_ASAP7_75t_L g150 ( .A(n_72), .Y(n_150) );
AND2x2_ASAP7_75t_L g196 ( .A(n_73), .B(n_165), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_74), .B(n_157), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_75), .A2(n_148), .B(n_498), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_76), .A2(n_148), .B(n_462), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_77), .A2(n_148), .B(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g517 ( .A(n_78), .B(n_174), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_79), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_80), .B(n_173), .Y(n_476) );
INVx1_ASAP7_75t_L g121 ( .A(n_81), .Y(n_121) );
AND2x2_ASAP7_75t_L g164 ( .A(n_82), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_83), .B(n_139), .Y(n_184) );
AND2x2_ASAP7_75t_L g465 ( .A(n_84), .B(n_134), .Y(n_465) );
AND2x2_ASAP7_75t_L g214 ( .A(n_85), .B(n_159), .Y(n_214) );
INVxp33_ASAP7_75t_L g796 ( .A(n_86), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_88), .B(n_157), .Y(n_183) );
AND2x2_ASAP7_75t_L g208 ( .A(n_89), .B(n_165), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_91), .B(n_155), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_92), .A2(n_148), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_93), .B(n_157), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_95), .A2(n_148), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_96), .B(n_155), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_97), .B(n_155), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_98), .Y(n_122) );
BUFx2_ASAP7_75t_L g544 ( .A(n_99), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_100), .Y(n_762) );
BUFx2_ASAP7_75t_L g108 ( .A(n_101), .Y(n_108) );
BUFx2_ASAP7_75t_SL g775 ( .A(n_101), .Y(n_775) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_102), .A2(n_148), .B(n_153), .Y(n_147) );
AOI21xp33_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_787), .B(n_795), .Y(n_103) );
OA21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_123), .B(n_772), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AOI21xp33_ASAP7_75t_SL g776 ( .A1(n_110), .A2(n_777), .B(n_780), .Y(n_776) );
NOR2xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_122), .Y(n_110) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g779 ( .A(n_115), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
OR2x6_ASAP7_75t_SL g451 ( .A(n_116), .B(n_117), .Y(n_451) );
AND2x6_ASAP7_75t_SL g759 ( .A(n_116), .B(n_118), .Y(n_759) );
OR2x2_ASAP7_75t_L g771 ( .A(n_116), .B(n_118), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_120), .B(n_121), .Y(n_794) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_760), .B(n_764), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22x1_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_449), .B1(n_452), .B2(n_756), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_127), .A2(n_453), .B1(n_766), .B2(n_767), .Y(n_765) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_370), .Y(n_127) );
NOR3xp33_ASAP7_75t_SL g128 ( .A(n_129), .B(n_282), .C(n_322), .Y(n_128) );
OAI221xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_197), .B1(n_246), .B2(n_261), .C(n_264), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_161), .Y(n_131) );
INVx2_ASAP7_75t_L g279 ( .A(n_132), .Y(n_279) );
AND2x2_ASAP7_75t_L g309 ( .A(n_132), .B(n_310), .Y(n_309) );
BUFx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g247 ( .A(n_133), .B(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g254 ( .A(n_133), .B(n_187), .Y(n_254) );
INVx2_ASAP7_75t_L g260 ( .A(n_133), .Y(n_260) );
AND2x2_ASAP7_75t_L g269 ( .A(n_133), .B(n_163), .Y(n_269) );
INVx1_ASAP7_75t_L g285 ( .A(n_133), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_133), .B(n_331), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_134), .A2(n_539), .B(n_540), .Y(n_538) );
BUFx4f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx3_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
AND2x4_ASAP7_75t_L g159 ( .A(n_136), .B(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_136), .B(n_160), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_147), .B(n_159), .Y(n_137) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_145), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
AND2x6_ASAP7_75t_L g157 ( .A(n_141), .B(n_150), .Y(n_157) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x4_ASAP7_75t_L g155 ( .A(n_143), .B(n_152), .Y(n_155) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx5_ASAP7_75t_L g158 ( .A(n_145), .Y(n_158) );
AND2x2_ASAP7_75t_L g151 ( .A(n_146), .B(n_152), .Y(n_151) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_146), .Y(n_482) );
AND2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
BUFx3_ASAP7_75t_L g483 ( .A(n_149), .Y(n_483) );
INVx2_ASAP7_75t_L g489 ( .A(n_150), .Y(n_489) );
AND2x4_ASAP7_75t_L g485 ( .A(n_151), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g481 ( .A(n_152), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_156), .B(n_158), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_157), .B(n_544), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_158), .A2(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_158), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_158), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_158), .A2(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_158), .A2(n_217), .B(n_218), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_158), .A2(n_225), .B(n_226), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_158), .A2(n_236), .B(n_237), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_158), .A2(n_463), .B(n_464), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_158), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_158), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_158), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_158), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_158), .A2(n_531), .B(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_158), .A2(n_542), .B(n_543), .Y(n_541) );
INVx1_ASAP7_75t_SL g178 ( .A(n_159), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_159), .B(n_220), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_159), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_159), .A2(n_505), .B(n_506), .Y(n_504) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_162), .B(n_175), .Y(n_161) );
INVx4_ASAP7_75t_L g250 ( .A(n_162), .Y(n_250) );
AND2x2_ASAP7_75t_L g281 ( .A(n_162), .B(n_188), .Y(n_281) );
AND2x2_ASAP7_75t_L g357 ( .A(n_162), .B(n_331), .Y(n_357) );
NAND2x1p5_ASAP7_75t_L g399 ( .A(n_162), .B(n_187), .Y(n_399) );
INVx5_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_163), .B(n_187), .Y(n_286) );
AND2x2_ASAP7_75t_L g310 ( .A(n_163), .B(n_188), .Y(n_310) );
BUFx2_ASAP7_75t_L g326 ( .A(n_163), .Y(n_326) );
NOR2x1_ASAP7_75t_SL g429 ( .A(n_163), .B(n_331), .Y(n_429) );
OR2x6_ASAP7_75t_L g163 ( .A(n_164), .B(n_167), .Y(n_163) );
INVx3_ASAP7_75t_L g207 ( .A(n_165), .Y(n_207) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_166), .A2(n_468), .B(n_474), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_173), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_173), .Y(n_195) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_173), .A2(n_234), .B(n_238), .Y(n_233) );
OA21x2_ASAP7_75t_L g296 ( .A1(n_173), .A2(n_234), .B(n_238), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_173), .A2(n_460), .B(n_461), .Y(n_459) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_173), .A2(n_478), .B(n_484), .Y(n_477) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g306 ( .A(n_175), .Y(n_306) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_175), .A2(n_373), .B1(n_375), .B2(n_377), .C(n_382), .Y(n_372) );
AND2x2_ASAP7_75t_L g392 ( .A(n_175), .B(n_285), .Y(n_392) );
AND2x4_ASAP7_75t_L g175 ( .A(n_176), .B(n_187), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g248 ( .A(n_177), .Y(n_248) );
INVx1_ASAP7_75t_L g301 ( .A(n_177), .Y(n_301) );
AO21x2_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_185), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_178), .B(n_186), .Y(n_185) );
AO21x2_ASAP7_75t_L g331 ( .A1(n_178), .A2(n_179), .B(n_185), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_184), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_187), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g270 ( .A(n_187), .B(n_258), .Y(n_270) );
INVx2_ASAP7_75t_L g312 ( .A(n_187), .Y(n_312) );
AND2x2_ASAP7_75t_L g445 ( .A(n_187), .B(n_260), .Y(n_445) );
INVx4_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_188), .Y(n_302) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_195), .B(n_196), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_194), .Y(n_189) );
AOI21x1_ASAP7_75t_L g527 ( .A1(n_195), .A2(n_528), .B(n_534), .Y(n_527) );
NOR3xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_229), .C(n_244), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_209), .Y(n_198) );
INVx2_ASAP7_75t_L g359 ( .A(n_199), .Y(n_359) );
AND2x2_ASAP7_75t_L g404 ( .A(n_199), .B(n_281), .Y(n_404) );
BUFx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g349 ( .A(n_200), .Y(n_349) );
AND2x4_ASAP7_75t_SL g364 ( .A(n_200), .B(n_276), .Y(n_364) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_207), .B(n_208), .Y(n_200) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_201), .A2(n_207), .B(n_208), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_206), .Y(n_201) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_207), .A2(n_222), .B(n_228), .Y(n_221) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_207), .A2(n_222), .B(n_228), .Y(n_241) );
AO21x1_ASAP7_75t_SL g510 ( .A1(n_207), .A2(n_511), .B(n_517), .Y(n_510) );
AO21x2_ASAP7_75t_L g568 ( .A1(n_207), .A2(n_511), .B(n_517), .Y(n_568) );
INVx2_ASAP7_75t_L g318 ( .A(n_209), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_209), .B(n_348), .Y(n_374) );
AND2x4_ASAP7_75t_L g407 ( .A(n_209), .B(n_354), .Y(n_407) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_221), .Y(n_209) );
AND2x2_ASAP7_75t_L g245 ( .A(n_210), .B(n_240), .Y(n_245) );
OR2x2_ASAP7_75t_L g275 ( .A(n_210), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_SL g344 ( .A(n_210), .B(n_296), .Y(n_344) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
BUFx2_ASAP7_75t_L g289 ( .A(n_211), .Y(n_289) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g263 ( .A(n_212), .Y(n_263) );
OAI21x1_ASAP7_75t_SL g212 ( .A1(n_213), .A2(n_215), .B(n_219), .Y(n_212) );
INVx1_ASAP7_75t_L g220 ( .A(n_214), .Y(n_220) );
INVx2_ASAP7_75t_L g276 ( .A(n_221), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_223), .B(n_227), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_229), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_239), .Y(n_230) );
AND2x2_ASAP7_75t_L g244 ( .A(n_231), .B(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g317 ( .A(n_231), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g402 ( .A(n_231), .Y(n_402) );
BUFx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x4_ASAP7_75t_L g262 ( .A(n_232), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g381 ( .A(n_232), .B(n_241), .Y(n_381) );
AND2x2_ASAP7_75t_L g385 ( .A(n_232), .B(n_251), .Y(n_385) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g354 ( .A(n_233), .Y(n_354) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_233), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_239), .B(n_262), .Y(n_338) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_240), .B(n_263), .Y(n_448) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g252 ( .A(n_241), .B(n_243), .Y(n_252) );
AND2x2_ASAP7_75t_L g334 ( .A(n_241), .B(n_296), .Y(n_334) );
AND2x2_ASAP7_75t_L g353 ( .A(n_241), .B(n_242), .Y(n_353) );
BUFx2_ASAP7_75t_L g274 ( .A(n_242), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_242), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
BUFx3_ASAP7_75t_L g251 ( .A(n_243), .Y(n_251) );
INVxp67_ASAP7_75t_L g294 ( .A(n_243), .Y(n_294) );
INVx1_ASAP7_75t_L g267 ( .A(n_245), .Y(n_267) );
AND2x2_ASAP7_75t_L g303 ( .A(n_245), .B(n_274), .Y(n_303) );
NAND2xp33_ASAP7_75t_L g384 ( .A(n_245), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g421 ( .A(n_245), .B(n_422), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_249), .B1(n_252), .B2(n_253), .C(n_255), .Y(n_246) );
AND2x2_ASAP7_75t_L g350 ( .A(n_247), .B(n_250), .Y(n_350) );
AND2x2_ASAP7_75t_SL g369 ( .A(n_247), .B(n_310), .Y(n_369) );
AND2x2_ASAP7_75t_L g387 ( .A(n_247), .B(n_312), .Y(n_387) );
AND2x2_ASAP7_75t_L g442 ( .A(n_247), .B(n_281), .Y(n_442) );
INVx1_ASAP7_75t_L g258 ( .A(n_248), .Y(n_258) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_248), .Y(n_314) );
CKINVDCx16_ASAP7_75t_R g394 ( .A(n_249), .Y(n_394) );
AND2x4_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_250), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_250), .B(n_301), .Y(n_376) );
AND2x2_ASAP7_75t_L g343 ( .A(n_251), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g379 ( .A(n_251), .Y(n_379) );
AND2x2_ASAP7_75t_L g288 ( .A(n_252), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_252), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g430 ( .A(n_252), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_252), .B(n_354), .Y(n_440) );
AND2x4_ASAP7_75t_L g356 ( .A(n_253), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g427 ( .A(n_254), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
OR2x2_ASAP7_75t_L g298 ( .A(n_259), .B(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g305 ( .A(n_260), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g336 ( .A(n_260), .B(n_310), .Y(n_336) );
AND2x2_ASAP7_75t_L g410 ( .A(n_260), .B(n_331), .Y(n_410) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g358 ( .A(n_262), .B(n_359), .Y(n_358) );
OAI32xp33_ASAP7_75t_L g423 ( .A1(n_262), .A2(n_424), .A3(n_426), .B1(n_427), .B2(n_430), .Y(n_423) );
AND2x4_ASAP7_75t_L g295 ( .A(n_263), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g393 ( .A(n_263), .B(n_296), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_268), .B1(n_271), .B2(n_277), .Y(n_264) );
INVxp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_SL g382 ( .A1(n_266), .A2(n_280), .B(n_383), .C(n_384), .Y(n_382) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g366 ( .A(n_267), .B(n_294), .Y(n_366) );
INVx1_ASAP7_75t_SL g437 ( .A(n_268), .Y(n_437) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
AND2x4_ASAP7_75t_L g340 ( .A(n_270), .B(n_279), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_270), .A2(n_419), .B1(n_420), .B2(n_421), .C(n_423), .Y(n_418) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_275), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OAI22xp33_ASAP7_75t_L g360 ( .A1(n_278), .A2(n_308), .B1(n_361), .B2(n_362), .Y(n_360) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
OAI211xp5_ASAP7_75t_SL g396 ( .A1(n_279), .A2(n_397), .B(n_405), .C(n_418), .Y(n_396) );
INVx2_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g316 ( .A(n_281), .B(n_285), .Y(n_316) );
OAI211xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_287), .B(n_290), .C(n_319), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g313 ( .A(n_285), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g433 ( .A(n_285), .B(n_429), .Y(n_433) );
OAI32xp33_ASAP7_75t_L g390 ( .A1(n_286), .A2(n_391), .A3(n_393), .B1(n_394), .B2(n_395), .Y(n_390) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_SL g380 ( .A(n_289), .B(n_381), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_297), .B1(n_303), .B2(n_304), .C(n_307), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g447 ( .A(n_294), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_295), .B(n_359), .Y(n_361) );
A2O1A1O1Ixp25_ASAP7_75t_L g432 ( .A1(n_295), .A2(n_364), .B(n_380), .C(n_426), .D(n_433), .Y(n_432) );
AOI31xp33_ASAP7_75t_L g434 ( .A1(n_295), .A2(n_316), .A3(n_426), .B(n_433), .Y(n_434) );
AND2x2_ASAP7_75t_L g348 ( .A(n_296), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_298), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx2_ASAP7_75t_L g425 ( .A(n_300), .Y(n_425) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g420 ( .A(n_301), .B(n_312), .Y(n_420) );
INVx1_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
AND2x2_ASAP7_75t_L g320 ( .A(n_304), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
AOI31xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_311), .A3(n_315), .B(n_317), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_310), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g443 ( .A(n_310), .B(n_389), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AND2x2_ASAP7_75t_L g388 ( .A(n_312), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g414 ( .A(n_312), .Y(n_414) );
INVxp67_ASAP7_75t_L g383 ( .A(n_313), .Y(n_383) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g321 ( .A(n_317), .Y(n_321) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND3xp33_ASAP7_75t_SL g322 ( .A(n_323), .B(n_339), .C(n_355), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_332), .B1(n_336), .B2(n_337), .Y(n_323) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx2_ASAP7_75t_L g409 ( .A(n_326), .Y(n_409) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVxp67_ASAP7_75t_SL g389 ( .A(n_330), .Y(n_389) );
INVxp67_ASAP7_75t_SL g415 ( .A(n_330), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_330), .B(n_399), .Y(n_416) );
NAND2xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
INVx1_ASAP7_75t_L g367 ( .A(n_334), .Y(n_367) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_350), .B2(n_351), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g341 ( .A(n_342), .B(n_345), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_348), .A2(n_353), .B1(n_387), .B2(n_388), .C(n_390), .Y(n_386) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2x1_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g426 ( .A(n_353), .Y(n_426) );
AND2x2_ASAP7_75t_L g363 ( .A(n_354), .B(n_364), .Y(n_363) );
O2A1O1Ixp33_ASAP7_75t_SL g411 ( .A1(n_354), .A2(n_412), .B(n_416), .C(n_417), .Y(n_411) );
AOI211xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_358), .B(n_360), .C(n_365), .Y(n_355) );
AND2x2_ASAP7_75t_L g406 ( .A(n_359), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g417 ( .A(n_364), .Y(n_417) );
AOI21xp33_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_367), .B(n_368), .Y(n_365) );
INVx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NOR3xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_396), .C(n_431), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_372), .B(n_386), .Y(n_371) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g395 ( .A(n_380), .Y(n_395) );
INVxp67_ASAP7_75t_L g419 ( .A(n_384), .Y(n_419) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g403 ( .A(n_393), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B1(n_403), .B2(n_404), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B(n_411), .Y(n_405) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g444 ( .A(n_429), .B(n_445), .Y(n_444) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .B1(n_435), .B2(n_438), .C(n_441), .Y(n_431) );
INVxp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI31xp33_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_443), .A3(n_444), .B(n_446), .Y(n_441) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx4f_ASAP7_75t_SL g766 ( .A(n_449), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
CKINVDCx11_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
INVx3_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
XNOR2xp5_ASAP7_75t_L g780 ( .A(n_453), .B(n_781), .Y(n_780) );
AND2x4_ASAP7_75t_SL g453 ( .A(n_454), .B(n_652), .Y(n_453) );
NOR3xp33_ASAP7_75t_SL g454 ( .A(n_455), .B(n_561), .C(n_593), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_490), .B1(n_518), .B2(n_535), .C(n_546), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_466), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g524 ( .A(n_458), .B(n_467), .Y(n_524) );
INVx4_ASAP7_75t_L g552 ( .A(n_458), .Y(n_552) );
AND2x4_ASAP7_75t_SL g592 ( .A(n_458), .B(n_526), .Y(n_592) );
BUFx2_ASAP7_75t_L g602 ( .A(n_458), .Y(n_602) );
NOR2x1_ASAP7_75t_L g668 ( .A(n_458), .B(n_607), .Y(n_668) );
AND2x2_ASAP7_75t_L g677 ( .A(n_458), .B(n_605), .Y(n_677) );
OR2x2_ASAP7_75t_L g685 ( .A(n_458), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g711 ( .A(n_458), .B(n_550), .Y(n_711) );
AND2x4_ASAP7_75t_L g730 ( .A(n_458), .B(n_731), .Y(n_730) );
OR2x6_ASAP7_75t_L g458 ( .A(n_459), .B(n_465), .Y(n_458) );
INVx2_ASAP7_75t_SL g643 ( .A(n_466), .Y(n_643) );
OR2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_475), .Y(n_466) );
AND2x2_ASAP7_75t_L g550 ( .A(n_467), .B(n_527), .Y(n_550) );
INVx2_ASAP7_75t_L g577 ( .A(n_467), .Y(n_577) );
INVx2_ASAP7_75t_L g607 ( .A(n_467), .Y(n_607) );
AND2x2_ASAP7_75t_L g621 ( .A(n_467), .B(n_526), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_473), .Y(n_468) );
AND2x2_ASAP7_75t_L g551 ( .A(n_475), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g574 ( .A(n_475), .Y(n_574) );
BUFx3_ASAP7_75t_L g588 ( .A(n_475), .Y(n_588) );
AND2x2_ASAP7_75t_L g617 ( .A(n_475), .B(n_618), .Y(n_617) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
AND2x4_ASAP7_75t_L g522 ( .A(n_476), .B(n_477), .Y(n_522) );
AND2x4_ASAP7_75t_L g479 ( .A(n_480), .B(n_483), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
NOR2x1p5_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g623 ( .A(n_490), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_501), .Y(n_490) );
OR2x2_ASAP7_75t_L g734 ( .A(n_491), .B(n_535), .Y(n_734) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g590 ( .A(n_492), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_492), .B(n_501), .Y(n_651) );
OR2x2_ASAP7_75t_L g749 ( .A(n_492), .B(n_671), .Y(n_749) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g560 ( .A(n_493), .B(n_536), .Y(n_560) );
OR2x2_ASAP7_75t_SL g570 ( .A(n_493), .B(n_571), .Y(n_570) );
INVx4_ASAP7_75t_L g581 ( .A(n_493), .Y(n_581) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_493), .Y(n_632) );
NAND2x1_ASAP7_75t_L g638 ( .A(n_493), .B(n_537), .Y(n_638) );
AND2x2_ASAP7_75t_L g663 ( .A(n_493), .B(n_503), .Y(n_663) );
OR2x2_ASAP7_75t_L g684 ( .A(n_493), .B(n_567), .Y(n_684) );
OR2x6_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g579 ( .A(n_501), .Y(n_579) );
O2A1O1Ixp33_ASAP7_75t_L g672 ( .A1(n_501), .A2(n_673), .B(n_676), .C(n_678), .Y(n_672) );
AND2x2_ASAP7_75t_L g745 ( .A(n_501), .B(n_521), .Y(n_745) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_510), .Y(n_501) );
INVx1_ASAP7_75t_L g612 ( .A(n_502), .Y(n_612) );
AND2x2_ASAP7_75t_L g682 ( .A(n_502), .B(n_537), .Y(n_682) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g556 ( .A(n_503), .Y(n_556) );
OR2x2_ASAP7_75t_L g571 ( .A(n_503), .B(n_537), .Y(n_571) );
INVx1_ASAP7_75t_L g587 ( .A(n_503), .Y(n_587) );
AND2x2_ASAP7_75t_L g599 ( .A(n_503), .B(n_510), .Y(n_599) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_503), .Y(n_705) );
NOR2x1_ASAP7_75t_SL g536 ( .A(n_510), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_516), .Y(n_511) );
INVxp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_523), .Y(n_519) );
OR2x2_ASAP7_75t_L g669 ( .A(n_520), .B(n_604), .Y(n_669) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_521), .B(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g751 ( .A(n_521), .B(n_648), .Y(n_751) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g596 ( .A(n_522), .B(n_577), .Y(n_596) );
AND2x2_ASAP7_75t_L g692 ( .A(n_522), .B(n_605), .Y(n_692) );
INVx1_ASAP7_75t_L g609 ( .A(n_523), .Y(n_609) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
INVx1_ASAP7_75t_L g659 ( .A(n_524), .Y(n_659) );
INVx2_ASAP7_75t_L g626 ( .A(n_525), .Y(n_626) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g576 ( .A(n_526), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g606 ( .A(n_526), .Y(n_606) );
INVx1_ASAP7_75t_L g731 ( .A(n_526), .Y(n_731) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_527), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_533), .Y(n_528) );
OR2x2_ASAP7_75t_L g702 ( .A(n_535), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_SL g557 ( .A(n_537), .Y(n_557) );
OR2x2_ASAP7_75t_L g580 ( .A(n_537), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g591 ( .A(n_537), .B(n_567), .Y(n_591) );
AND2x2_ASAP7_75t_L g665 ( .A(n_537), .B(n_581), .Y(n_665) );
BUFx2_ASAP7_75t_L g748 ( .A(n_537), .Y(n_748) );
OR2x6_ASAP7_75t_L g537 ( .A(n_538), .B(n_545), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_553), .B(n_558), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_551), .Y(n_548) );
AND2x2_ASAP7_75t_L g700 ( .A(n_549), .B(n_622), .Y(n_700) );
BUFx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g559 ( .A(n_550), .B(n_552), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_551), .B(n_621), .Y(n_722) );
INVx1_ASAP7_75t_L g752 ( .A(n_551), .Y(n_752) );
NAND2x1p5_ASAP7_75t_L g648 ( .A(n_552), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_552), .B(n_688), .Y(n_725) );
INVxp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
AND2x4_ASAP7_75t_SL g589 ( .A(n_555), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_555), .B(n_583), .Y(n_736) );
INVx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_556), .B(n_638), .Y(n_694) );
AND2x2_ASAP7_75t_L g712 ( .A(n_556), .B(n_665), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_557), .B(n_599), .Y(n_615) );
A2O1A1Ixp33_ASAP7_75t_L g644 ( .A1(n_557), .A2(n_603), .B(n_645), .C(n_650), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_557), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_559), .A2(n_632), .B1(n_740), .B2(n_746), .C(n_750), .Y(n_739) );
INVx1_ASAP7_75t_SL g727 ( .A(n_560), .Y(n_727) );
OAI221xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_572), .B1(n_578), .B2(n_582), .C(n_798), .Y(n_561) );
INVx2_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_569), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g637 ( .A(n_566), .Y(n_637) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g611 ( .A(n_567), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g642 ( .A(n_567), .B(n_587), .Y(n_642) );
INVx2_ASAP7_75t_L g675 ( .A(n_567), .Y(n_675) );
INVx3_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI32xp33_ASAP7_75t_L g726 ( .A1(n_570), .A2(n_617), .A3(n_648), .B1(n_727), .B2(n_728), .Y(n_726) );
OR2x2_ASAP7_75t_L g697 ( .A(n_571), .B(n_684), .Y(n_697) );
INVx1_ASAP7_75t_L g707 ( .A(n_572), .Y(n_707) );
OR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
INVx2_ASAP7_75t_L g622 ( .A(n_573), .Y(n_622) );
AND2x2_ASAP7_75t_L g693 ( .A(n_573), .B(n_668), .Y(n_693) );
OR2x2_ASAP7_75t_L g724 ( .A(n_573), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_574), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g618 ( .A(n_577), .Y(n_618) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx2_ASAP7_75t_SL g583 ( .A(n_580), .Y(n_583) );
OR2x2_ASAP7_75t_L g670 ( .A(n_580), .B(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_581), .B(n_599), .Y(n_598) );
NOR2xp67_ASAP7_75t_L g704 ( .A(n_581), .B(n_705), .Y(n_704) );
BUFx2_ASAP7_75t_L g717 ( .A(n_581), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B(n_589), .C(n_592), .Y(n_582) );
AND2x2_ASAP7_75t_L g732 ( .A(n_584), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g658 ( .A(n_588), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_588), .B(n_592), .Y(n_679) );
AND2x2_ASAP7_75t_L g710 ( .A(n_588), .B(n_711), .Y(n_710) );
O2A1O1Ixp33_ASAP7_75t_L g720 ( .A1(n_590), .A2(n_721), .B(n_723), .C(n_726), .Y(n_720) );
AOI222xp33_ASAP7_75t_L g594 ( .A1(n_591), .A2(n_595), .B1(n_597), .B2(n_600), .C1(n_608), .C2(n_610), .Y(n_594) );
AND2x2_ASAP7_75t_L g662 ( .A(n_591), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g595 ( .A(n_592), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_SL g616 ( .A(n_592), .Y(n_616) );
NAND4xp25_ASAP7_75t_L g593 ( .A(n_594), .B(n_613), .C(n_634), .D(n_644), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_596), .B(n_602), .Y(n_656) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g664 ( .A(n_599), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_SL g671 ( .A(n_599), .Y(n_671) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_601), .A2(n_635), .B(n_639), .C(n_643), .Y(n_634) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_602), .B(n_617), .Y(n_738) );
OR2x2_ASAP7_75t_L g742 ( .A(n_602), .B(n_628), .Y(n_742) );
INVx1_ASAP7_75t_L g715 ( .A(n_603), .Y(n_715) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_SL g649 ( .A(n_606), .Y(n_649) );
INVx1_ASAP7_75t_L g629 ( .A(n_607), .Y(n_629) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_609), .B(n_646), .Y(n_645) );
BUFx2_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g633 ( .A(n_611), .Y(n_633) );
AOI322xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .A3(n_617), .B1(n_619), .B2(n_623), .C1(n_624), .C2(n_630), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_SL g695 ( .A1(n_616), .A2(n_696), .B(n_697), .C(n_698), .Y(n_695) );
INVx1_ASAP7_75t_L g718 ( .A(n_617), .Y(n_718) );
NOR2xp67_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g676 ( .A(n_622), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_628), .Y(n_698) );
INVx2_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx3_ASAP7_75t_L g641 ( .A(n_638), .Y(n_641) );
OR2x2_ASAP7_75t_L g709 ( .A(n_638), .B(n_671), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_638), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_SL g741 ( .A(n_642), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_643), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND3xp33_ASAP7_75t_SL g746 ( .A(n_651), .B(n_747), .C(n_749), .Y(n_746) );
NOR3xp33_ASAP7_75t_SL g652 ( .A(n_653), .B(n_690), .C(n_719), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_654), .B(n_672), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .B(n_660), .C(n_666), .Y(n_654) );
OAI31xp33_ASAP7_75t_L g699 ( .A1(n_655), .A2(n_677), .A3(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
INVx2_ASAP7_75t_L g714 ( .A(n_662), .Y(n_714) );
INVx1_ASAP7_75t_L g689 ( .A(n_664), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B(n_670), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g716 ( .A(n_674), .B(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g755 ( .A(n_675), .Y(n_755) );
OAI22xp33_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_680), .B1(n_685), .B2(n_689), .Y(n_678) );
INVx3_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x4_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_684), .Y(n_696) );
OR2x2_ASAP7_75t_L g747 ( .A(n_684), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND3xp33_ASAP7_75t_SL g690 ( .A(n_691), .B(n_699), .C(n_706), .Y(n_690) );
O2A1O1Ixp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B(n_694), .C(n_695), .Y(n_691) );
INVx2_ASAP7_75t_L g728 ( .A(n_692), .Y(n_728) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B1(n_710), .B2(n_712), .C(n_713), .Y(n_706) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI22xp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B1(n_716), .B2(n_718), .Y(n_713) );
NAND3xp33_ASAP7_75t_SL g719 ( .A(n_720), .B(n_729), .C(n_739), .Y(n_719) );
INVxp33_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_732), .B1(n_735), .B2(n_737), .Y(n_729) );
INVx2_ASAP7_75t_L g743 ( .A(n_730), .Y(n_743) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_742), .B1(n_743), .B2(n_744), .Y(n_740) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI22xp33_ASAP7_75t_SL g750 ( .A1(n_749), .A2(n_751), .B1(n_752), .B2(n_753), .Y(n_750) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
CKINVDCx6p67_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
INVx4_ASAP7_75t_SL g767 ( .A(n_757), .Y(n_767) );
INVx3_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_759), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_760), .A2(n_765), .B(n_768), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
BUFx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_776), .Y(n_772) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
CKINVDCx16_ASAP7_75t_R g783 ( .A(n_784), .Y(n_783) );
BUFx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_788), .B(n_796), .Y(n_795) );
INVx3_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g789 ( .A(n_790), .B(n_794), .Y(n_789) );
endmodule