module fake_jpeg_28260_n_240 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_240);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_240;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_32),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_5),
.C(n_9),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_22),
.B(n_20),
.C(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_18),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_16),
.B1(n_14),
.B2(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_20),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_16),
.B1(n_19),
.B2(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_50),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_49),
.Y(n_64)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_58),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_16),
.B1(n_18),
.B2(n_17),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_25),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_24),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_32),
.B1(n_28),
.B2(n_24),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_44),
.B1(n_36),
.B2(n_12),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_61),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_12),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_33),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_71),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_48),
.B1(n_57),
.B2(n_60),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_33),
.B1(n_38),
.B2(n_36),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_55),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_0),
.B(n_1),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_44),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_78),
.B1(n_48),
.B2(n_51),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_28),
.B1(n_24),
.B2(n_31),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_28),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_54),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_31),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_82),
.B(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_15),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_54),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_71),
.A2(n_55),
.B1(n_58),
.B2(n_52),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_85),
.A2(n_81),
.B1(n_53),
.B2(n_72),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_109),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_96),
.B(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_89),
.B(n_90),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_47),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_69),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_91),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_97),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_73),
.B1(n_81),
.B2(n_80),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_45),
.B(n_53),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_7),
.B(n_10),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_15),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_15),
.Y(n_98)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_69),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_30),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_101),
.B(n_105),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_30),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_0),
.Y(n_104)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

OA21x2_ASAP7_75t_L g106 ( 
.A1(n_83),
.A2(n_63),
.B(n_60),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_106),
.A2(n_66),
.B(n_73),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_70),
.B1(n_74),
.B2(n_65),
.Y(n_107)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_66),
.A2(n_63),
.B1(n_53),
.B2(n_6),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_84),
.B1(n_72),
.B2(n_75),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_0),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_112),
.B(n_119),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_64),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_64),
.C(n_80),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_117),
.C(n_90),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_116),
.B(n_124),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_88),
.C(n_109),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_128),
.B1(n_129),
.B2(n_132),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_103),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_120),
.A2(n_131),
.B1(n_108),
.B2(n_96),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_125),
.B(n_100),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_81),
.B1(n_75),
.B2(n_84),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_85),
.A2(n_84),
.B1(n_75),
.B2(n_6),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_102),
.A2(n_5),
.B1(n_9),
.B2(n_8),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_98),
.A2(n_5),
.B1(n_9),
.B2(n_8),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_89),
.B1(n_106),
.B2(n_108),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_10),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_126),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_115),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_88),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_141),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_101),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_104),
.C(n_85),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_148),
.C(n_163),
.Y(n_166)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_146),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_92),
.C(n_97),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_SL g181 ( 
.A(n_145),
.B(n_159),
.C(n_132),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_91),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_95),
.C(n_107),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_95),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_114),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_150),
.A2(n_153),
.B1(n_161),
.B2(n_162),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_94),
.Y(n_151)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_99),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_152),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_96),
.B1(n_107),
.B2(n_106),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_157),
.A2(n_161),
.B1(n_156),
.B2(n_120),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_110),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_160),
.B(n_144),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_106),
.C(n_4),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_169),
.B1(n_173),
.B2(n_150),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_176),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_163),
.A2(n_135),
.B1(n_119),
.B2(n_112),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_135),
.B1(n_112),
.B2(n_119),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_178),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_115),
.C(n_133),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_175),
.B(n_123),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_133),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_123),
.Y(n_178)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_140),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_184),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_147),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_155),
.B(n_158),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_185),
.A2(n_195),
.B(n_157),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_162),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_193),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_172),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_187),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_164),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_155),
.B(n_148),
.C(n_144),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_190),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_151),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_193),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_202),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_166),
.C(n_175),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_167),
.C(n_189),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_178),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_205),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_166),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_206),
.A2(n_169),
.B1(n_188),
.B2(n_185),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_183),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_170),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_174),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_176),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_214),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_203),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_213),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_211),
.B(n_216),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_198),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_171),
.C(n_179),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_204),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_200),
.B(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_200),
.B(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_206),
.B1(n_121),
.B2(n_196),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_156),
.B1(n_125),
.B2(n_134),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_181),
.B(n_196),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_225),
.B(n_215),
.Y(n_226)
);

NOR3xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_228),
.C(n_218),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_205),
.C(n_208),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_231),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_4),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_L g236 ( 
.A1(n_232),
.A2(n_235),
.A3(n_228),
.B1(n_3),
.B2(n_7),
.C1(n_1),
.C2(n_2),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_221),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_3),
.B(n_1),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g235 ( 
.A1(n_229),
.A2(n_160),
.A3(n_6),
.B1(n_3),
.B2(n_7),
.C1(n_9),
.C2(n_2),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_236),
.A2(n_237),
.B(n_233),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_0),
.C(n_1),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_2),
.Y(n_240)
);


endmodule