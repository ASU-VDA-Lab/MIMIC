module fake_ibex_951_n_751 (n_85, n_84, n_64, n_3, n_73, n_65, n_103, n_95, n_55, n_63, n_98, n_29, n_106, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_93, n_13, n_61, n_14, n_0, n_94, n_12, n_42, n_77, n_112, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_100, n_72, n_26, n_34, n_97, n_102, n_15, n_24, n_52, n_99, n_105, n_1, n_111, n_25, n_36, n_104, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_107, n_50, n_11, n_92, n_101, n_113, n_96, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_751);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_103;
input n_95;
input n_55;
input n_63;
input n_98;
input n_29;
input n_106;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_93;
input n_13;
input n_61;
input n_14;
input n_0;
input n_94;
input n_12;
input n_42;
input n_77;
input n_112;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_34;
input n_97;
input n_102;
input n_15;
input n_24;
input n_52;
input n_99;
input n_105;
input n_1;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_50;
input n_11;
input n_92;
input n_101;
input n_113;
input n_96;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_751;

wire n_151;
wire n_599;
wire n_507;
wire n_743;
wire n_540;
wire n_395;
wire n_171;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_688;
wire n_130;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_124;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_638;
wire n_398;
wire n_304;
wire n_125;
wire n_191;
wire n_593;
wire n_153;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_134;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_412;
wire n_357;
wire n_457;
wire n_494;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_421;
wire n_738;
wire n_475;
wire n_166;
wire n_163;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_114;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_375;
wire n_340;
wire n_698;
wire n_187;
wire n_667;
wire n_154;
wire n_682;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_723;
wire n_144;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_561;
wire n_117;
wire n_417;
wire n_471;
wire n_739;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_147;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_598;
wire n_143;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_127;
wire n_121;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_120;
wire n_168;
wire n_526;
wire n_155;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_122;
wire n_523;
wire n_116;
wire n_694;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_750;
wire n_746;
wire n_136;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_355;
wire n_474;
wire n_281;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_156;
wire n_570;
wire n_126;
wire n_623;
wire n_585;
wire n_715;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_141;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_454;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_146;
wire n_207;
wire n_438;
wire n_689;
wire n_167;
wire n_676;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_618;
wire n_514;
wire n_139;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_129;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_347;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_262;
wire n_433;
wire n_299;
wire n_439;
wire n_704;
wire n_643;
wire n_137;
wire n_679;
wire n_338;
wire n_173;
wire n_696;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_257;
wire n_718;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_140;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_546;
wire n_199;
wire n_592;
wire n_495;
wire n_410;
wire n_308;
wire n_675;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_135;
wire n_520;
wire n_684;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_115;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_138;
wire n_650;
wire n_409;
wire n_582;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_332;
wire n_517;
wire n_211;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_132;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_247;
wire n_379;
wire n_320;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_148;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_118;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_198;
wire n_264;
wire n_616;
wire n_217;
wire n_324;
wire n_391;
wire n_537;
wire n_728;
wire n_670;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_668;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_119;
wire n_361;
wire n_455;
wire n_419;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_131;
wire n_123;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_462;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_149;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_159;
wire n_231;
wire n_202;
wire n_298;
wire n_587;
wire n_160;
wire n_657;
wire n_184;
wire n_492;
wire n_649;
wire n_232;
wire n_380;
wire n_749;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g114 ( 
.A(n_24),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVxp33_ASAP7_75t_SL g116 ( 
.A(n_85),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_23),
.Y(n_117)
);

INVxp67_ASAP7_75t_SL g118 ( 
.A(n_93),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_42),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_18),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_19),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_41),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_29),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_11),
.Y(n_129)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_30),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_51),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_68),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_10),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_38),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_53),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_21),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_1),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

BUFx10_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_109),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

BUFx2_ASAP7_75t_SL g143 ( 
.A(n_58),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_28),
.Y(n_144)
);

BUFx2_ASAP7_75t_SL g145 ( 
.A(n_47),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_0),
.Y(n_148)
);

INVxp33_ASAP7_75t_SL g149 ( 
.A(n_84),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_10),
.Y(n_151)
);

NOR2xp67_ASAP7_75t_L g152 ( 
.A(n_81),
.B(n_86),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

BUFx2_ASAP7_75t_SL g155 ( 
.A(n_77),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_76),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_26),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_11),
.Y(n_159)
);

INVxp67_ASAP7_75t_SL g160 ( 
.A(n_69),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_2),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_56),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_50),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_110),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_79),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_60),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_22),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_80),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_96),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_17),
.Y(n_174)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_57),
.Y(n_175)
);

INVxp67_ASAP7_75t_SL g176 ( 
.A(n_20),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_3),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_48),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_101),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_14),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_78),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_31),
.Y(n_183)
);

NOR2xp67_ASAP7_75t_L g184 ( 
.A(n_3),
.B(n_2),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_32),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

INVxp33_ASAP7_75t_SL g188 ( 
.A(n_25),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_14),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_62),
.Y(n_191)
);

INVx4_ASAP7_75t_R g192 ( 
.A(n_43),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_19),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_17),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_67),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_4),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_83),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_54),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_194),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_126),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_124),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_147),
.B(n_0),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_129),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_140),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_1),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_124),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_186),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_138),
.Y(n_216)
);

NAND2xp33_ASAP7_75t_SL g217 ( 
.A(n_130),
.B(n_4),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_127),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

NOR2xp67_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_5),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_140),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_133),
.B(n_130),
.Y(n_222)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_140),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_127),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_123),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_134),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_141),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_134),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_142),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_5),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_148),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_141),
.B(n_45),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_151),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_156),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_162),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_133),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_142),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_114),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_114),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_156),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_191),
.Y(n_247)
);

AND2x4_ASAP7_75t_L g248 ( 
.A(n_161),
.B(n_6),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_161),
.B(n_6),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_128),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_191),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_128),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_120),
.B(n_7),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_135),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_159),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_135),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_197),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_136),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_136),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_143),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_197),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_165),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_115),
.B(n_7),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_165),
.B(n_117),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_116),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_116),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_121),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_149),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_122),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_149),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_125),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_139),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_131),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_144),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_248),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_230),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_222),
.B(n_146),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_230),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_230),
.Y(n_279)
);

AND2x4_ASAP7_75t_L g280 ( 
.A(n_214),
.B(n_150),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_208),
.B(n_132),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_199),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_231),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_231),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_206),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_224),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_237),
.Y(n_287)
);

AND2x6_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_210),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_206),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_224),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_211),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_221),
.B(n_260),
.Y(n_293)
);

AND2x4_ASAP7_75t_L g294 ( 
.A(n_221),
.B(n_209),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_211),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_246),
.B(n_188),
.Y(n_297)
);

AND2x6_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_198),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_199),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_199),
.Y(n_300)
);

NAND2x1p5_ASAP7_75t_L g301 ( 
.A(n_244),
.B(n_195),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_199),
.Y(n_302)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_207),
.Y(n_303)
);

BUFx4f_ASAP7_75t_L g304 ( 
.A(n_207),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_226),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_228),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_255),
.B(n_137),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_267),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_246),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_212),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_247),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_267),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_267),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g314 ( 
.A(n_233),
.B(n_249),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_256),
.B(n_273),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_267),
.Y(n_316)
);

AND2x6_ASAP7_75t_L g317 ( 
.A(n_204),
.B(n_169),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_212),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_212),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_207),
.B(n_173),
.Y(n_321)
);

AND2x4_ASAP7_75t_L g322 ( 
.A(n_203),
.B(n_153),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_250),
.B(n_168),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_247),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_252),
.B(n_170),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_271),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_218),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_223),
.B(n_205),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_215),
.A2(n_188),
.B1(n_160),
.B2(n_118),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_223),
.B(n_143),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_241),
.Y(n_331)
);

AND2x6_ASAP7_75t_L g332 ( 
.A(n_243),
.B(n_171),
.Y(n_332)
);

A2O1A1Ixp33_ASAP7_75t_L g333 ( 
.A1(n_243),
.A2(n_178),
.B(n_189),
.C(n_187),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_271),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_229),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_254),
.B(n_164),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_271),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_227),
.Y(n_338)
);

NOR2x1p5_ASAP7_75t_L g339 ( 
.A(n_201),
.B(n_175),
.Y(n_339)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_241),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_241),
.Y(n_341)
);

NAND2x1p5_ASAP7_75t_L g342 ( 
.A(n_258),
.B(n_163),
.Y(n_342)
);

NAND3xp33_ASAP7_75t_L g343 ( 
.A(n_216),
.B(n_166),
.C(n_185),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_241),
.Y(n_344)
);

NAND3x1_ASAP7_75t_L g345 ( 
.A(n_253),
.B(n_182),
.C(n_154),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_262),
.B(n_180),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_257),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_235),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_232),
.B(n_157),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_225),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_257),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_257),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_259),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_251),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_223),
.Y(n_355)
);

AND2x2_ASAP7_75t_SL g356 ( 
.A(n_253),
.B(n_179),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_259),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_234),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_264),
.B(n_176),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_236),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_225),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_219),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_272),
.B(n_158),
.Y(n_363)
);

NAND2x1p5_ASAP7_75t_L g364 ( 
.A(n_264),
.B(n_239),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_269),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_269),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_238),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_217),
.A2(n_155),
.B1(n_145),
.B2(n_152),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_240),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_263),
.Y(n_370)
);

AOI22x1_ASAP7_75t_L g371 ( 
.A1(n_274),
.A2(n_155),
.B1(n_145),
.B2(n_192),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_311),
.B(n_201),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_370),
.B(n_268),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_309),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_370),
.B(n_268),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_370),
.B(n_265),
.Y(n_376)
);

NOR3xp33_ASAP7_75t_SL g377 ( 
.A(n_286),
.B(n_265),
.C(n_266),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_291),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_275),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_270),
.Y(n_380)
);

NAND2x1p5_ASAP7_75t_L g381 ( 
.A(n_327),
.B(n_304),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_322),
.B(n_220),
.Y(n_382)
);

NAND2x1p5_ASAP7_75t_L g383 ( 
.A(n_304),
.B(n_242),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_277),
.B(n_215),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_291),
.Y(n_385)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_288),
.Y(n_386)
);

AO22x1_ASAP7_75t_L g387 ( 
.A1(n_309),
.A2(n_245),
.B1(n_200),
.B2(n_217),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_283),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_322),
.B(n_200),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_284),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_315),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_277),
.B(n_8),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_8),
.Y(n_393)
);

NOR2x1p5_ASAP7_75t_L g394 ( 
.A(n_290),
.B(n_213),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_285),
.Y(n_395)
);

NOR2x1_ASAP7_75t_L g396 ( 
.A(n_343),
.B(n_213),
.Y(n_396)
);

OR2x6_ASAP7_75t_L g397 ( 
.A(n_348),
.B(n_202),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_349),
.B(n_9),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_307),
.B(n_202),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_335),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_R g401 ( 
.A(n_324),
.B(n_9),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_294),
.B(n_12),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_354),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_R g404 ( 
.A(n_297),
.B(n_49),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_289),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_292),
.Y(n_407)
);

CKINVDCx8_ASAP7_75t_R g408 ( 
.A(n_280),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_359),
.B(n_52),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_294),
.B(n_12),
.Y(n_410)
);

NOR2x2_ASAP7_75t_L g411 ( 
.A(n_339),
.B(n_13),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_354),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_328),
.B(n_55),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_300),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_328),
.B(n_13),
.Y(n_415)
);

BUFx4f_ASAP7_75t_L g416 ( 
.A(n_288),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_359),
.B(n_15),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_295),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_295),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_338),
.Y(n_420)
);

NOR3xp33_ASAP7_75t_SL g421 ( 
.A(n_333),
.B(n_287),
.C(n_323),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_293),
.B(n_59),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_275),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_338),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_SL g425 ( 
.A(n_329),
.B(n_15),
.C(n_16),
.Y(n_425)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_298),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_301),
.B(n_64),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_321),
.B(n_16),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_363),
.B(n_18),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_305),
.B(n_27),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_301),
.B(n_33),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_350),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_280),
.B(n_34),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_363),
.Y(n_434)
);

CKINVDCx6p67_ASAP7_75t_R g435 ( 
.A(n_317),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_365),
.Y(n_436)
);

OR2x6_ASAP7_75t_L g437 ( 
.A(n_355),
.B(n_342),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_281),
.B(n_35),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_300),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_330),
.B(n_36),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_300),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_300),
.Y(n_442)
);

OR2x6_ASAP7_75t_SL g443 ( 
.A(n_287),
.B(n_37),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_355),
.B(n_39),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_350),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_296),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_303),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_365),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_356),
.A2(n_40),
.B1(n_46),
.B2(n_65),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_361),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_293),
.B(n_71),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_362),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_306),
.B(n_72),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_366),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_288),
.A2(n_74),
.B1(n_75),
.B2(n_82),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_303),
.B(n_356),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_426),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_426),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_426),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_437),
.B(n_360),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_385),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_385),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_373),
.A2(n_279),
.B(n_276),
.Y(n_463)
);

CKINVDCx8_ASAP7_75t_R g464 ( 
.A(n_397),
.Y(n_464)
);

NOR3xp33_ASAP7_75t_L g465 ( 
.A(n_384),
.B(n_333),
.C(n_323),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_385),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_434),
.B(n_288),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_412),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_386),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_430),
.A2(n_342),
.B(n_371),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_373),
.B(n_317),
.Y(n_471)
);

A2O1A1Ixp33_ASAP7_75t_L g472 ( 
.A1(n_421),
.A2(n_278),
.B(n_358),
.C(n_346),
.Y(n_472)
);

OAI221xp5_ASAP7_75t_L g473 ( 
.A1(n_408),
.A2(n_368),
.B1(n_364),
.B2(n_346),
.C(n_369),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_386),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_374),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_420),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_416),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_393),
.A2(n_314),
.B1(n_368),
.B2(n_353),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_437),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_388),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_390),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_393),
.A2(n_314),
.B1(n_298),
.B2(n_317),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_379),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_403),
.Y(n_484)
);

AO32x1_ASAP7_75t_L g485 ( 
.A1(n_438),
.A2(n_310),
.A3(n_331),
.B1(n_344),
.B2(n_320),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_391),
.B(n_367),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_375),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_379),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_395),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_424),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_375),
.A2(n_352),
.B(n_351),
.Y(n_491)
);

NOR2xp67_ASAP7_75t_L g492 ( 
.A(n_455),
.B(n_357),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_398),
.A2(n_298),
.B1(n_317),
.B2(n_332),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_437),
.B(n_298),
.Y(n_494)
);

A2O1A1Ixp33_ASAP7_75t_L g495 ( 
.A1(n_392),
.A2(n_325),
.B(n_336),
.C(n_347),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_389),
.B(n_364),
.Y(n_496)
);

BUFx5_ASAP7_75t_L g497 ( 
.A(n_454),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_380),
.B(n_317),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_405),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_398),
.A2(n_298),
.B1(n_336),
.B2(n_325),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_407),
.Y(n_501)
);

BUFx4f_ASAP7_75t_L g502 ( 
.A(n_389),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_399),
.B(n_303),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_423),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_397),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_402),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_402),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_416),
.A2(n_345),
.B1(n_347),
.B2(n_316),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_446),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_397),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_452),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_380),
.B(n_332),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_428),
.A2(n_456),
.B1(n_410),
.B2(n_425),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_410),
.B(n_332),
.Y(n_514)
);

AOI221xp5_ASAP7_75t_L g515 ( 
.A1(n_387),
.A2(n_316),
.B1(n_326),
.B2(n_334),
.C(n_337),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_440),
.B(n_340),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_377),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_372),
.B(n_326),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_435),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_423),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_448),
.Y(n_521)
);

NOR2xp67_ASAP7_75t_L g522 ( 
.A(n_455),
.B(n_340),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_417),
.A2(n_332),
.B1(n_313),
.B2(n_312),
.Y(n_523)
);

INVx3_ASAP7_75t_SL g524 ( 
.A(n_411),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_450),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_428),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_376),
.B(n_332),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_447),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_443),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_433),
.B(n_340),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_451),
.B(n_318),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_453),
.A2(n_308),
.B(n_310),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_449),
.A2(n_451),
.B1(n_440),
.B2(n_429),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_378),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_418),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_382),
.B(n_299),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_381),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_401),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_448),
.Y(n_539)
);

OR2x2_ASAP7_75t_SL g540 ( 
.A(n_394),
.B(n_282),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_400),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_479),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_475),
.B(n_396),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_480),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_481),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_502),
.A2(n_396),
.B1(n_415),
.B2(n_409),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_489),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_468),
.B(n_419),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_502),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_476),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_SL g551 ( 
.A(n_494),
.B(n_404),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_529),
.A2(n_444),
.B1(n_445),
.B2(n_432),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_533),
.A2(n_422),
.B(n_436),
.Y(n_553)
);

CKINVDCx11_ASAP7_75t_R g554 ( 
.A(n_464),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_482),
.A2(n_413),
.B1(n_431),
.B2(n_427),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_499),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_533),
.A2(n_522),
.B1(n_493),
.B2(n_478),
.Y(n_557)
);

AOI221xp5_ASAP7_75t_L g558 ( 
.A1(n_465),
.A2(n_383),
.B1(n_406),
.B2(n_341),
.C(n_319),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_L g559 ( 
.A1(n_484),
.A2(n_319),
.B1(n_341),
.B2(n_302),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_501),
.Y(n_560)
);

AOI32xp33_ASAP7_75t_L g561 ( 
.A1(n_513),
.A2(n_87),
.A3(n_88),
.B1(n_89),
.B2(n_95),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_490),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_509),
.B(n_414),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_486),
.B(n_460),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_460),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_525),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_496),
.A2(n_414),
.B1(n_439),
.B2(n_441),
.Y(n_567)
);

NAND2x1_ASAP7_75t_L g568 ( 
.A(n_458),
.B(n_414),
.Y(n_568)
);

AO21x1_ASAP7_75t_L g569 ( 
.A1(n_478),
.A2(n_302),
.B(n_319),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_522),
.A2(n_302),
.B1(n_319),
.B2(n_341),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_524),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_479),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_503),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_517),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_511),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_462),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_493),
.A2(n_302),
.B1(n_439),
.B2(n_442),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_506),
.B(n_442),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_494),
.B(n_507),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_492),
.A2(n_472),
.B1(n_487),
.B2(n_500),
.Y(n_580)
);

OAI22xp33_ASAP7_75t_L g581 ( 
.A1(n_505),
.A2(n_510),
.B1(n_487),
.B2(n_538),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_526),
.A2(n_473),
.B1(n_467),
.B2(n_514),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_527),
.A2(n_508),
.B1(n_492),
.B2(n_498),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_528),
.Y(n_584)
);

NAND3xp33_ASAP7_75t_SL g585 ( 
.A(n_515),
.B(n_508),
.C(n_518),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_516),
.A2(n_523),
.B1(n_495),
.B2(n_531),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_469),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_540),
.B(n_537),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_SL g589 ( 
.A(n_463),
.B(n_523),
.C(n_530),
.Y(n_589)
);

OAI22xp33_ASAP7_75t_L g590 ( 
.A1(n_519),
.A2(n_471),
.B1(n_512),
.B2(n_535),
.Y(n_590)
);

OA21x2_ASAP7_75t_L g591 ( 
.A1(n_470),
.A2(n_532),
.B(n_491),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_520),
.Y(n_592)
);

INVx4_ASAP7_75t_SL g593 ( 
.A(n_457),
.Y(n_593)
);

AO21x2_ASAP7_75t_L g594 ( 
.A1(n_485),
.A2(n_539),
.B(n_521),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_527),
.B(n_536),
.Y(n_595)
);

INVxp33_ASAP7_75t_L g596 ( 
.A(n_536),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_504),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_534),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_534),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_497),
.B(n_488),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_519),
.B(n_483),
.Y(n_601)
);

CKINVDCx14_ASAP7_75t_R g602 ( 
.A(n_477),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_462),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_497),
.B(n_488),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_541),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_541),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_497),
.B(n_483),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_L g608 ( 
.A(n_497),
.B(n_474),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_497),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_462),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_466),
.Y(n_611)
);

BUFx12f_ASAP7_75t_L g612 ( 
.A(n_477),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_469),
.B(n_474),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_477),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_461),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_458),
.B(n_469),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_466),
.B(n_474),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_466),
.Y(n_618)
);

AO22x1_ASAP7_75t_SL g619 ( 
.A1(n_457),
.A2(n_524),
.B1(n_464),
.B2(n_389),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_457),
.B(n_459),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_459),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_459),
.B(n_485),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_564),
.B(n_565),
.Y(n_623)
);

AOI221xp5_ASAP7_75t_L g624 ( 
.A1(n_557),
.A2(n_573),
.B1(n_556),
.B2(n_560),
.C(n_545),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_557),
.A2(n_585),
.B1(n_582),
.B2(n_543),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_544),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_591),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_583),
.A2(n_580),
.B1(n_553),
.B2(n_552),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g629 ( 
.A(n_550),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_612),
.Y(n_630)
);

AOI222xp33_ASAP7_75t_L g631 ( 
.A1(n_554),
.A2(n_566),
.B1(n_562),
.B2(n_547),
.C1(n_575),
.C2(n_581),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_591),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_576),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_596),
.B(n_549),
.Y(n_634)
);

AOI221xp5_ASAP7_75t_L g635 ( 
.A1(n_580),
.A2(n_586),
.B1(n_592),
.B2(n_546),
.C(n_551),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_548),
.B(n_588),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_589),
.A2(n_586),
.B1(n_595),
.B2(n_558),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_602),
.Y(n_638)
);

NOR2x1_ASAP7_75t_SL g639 ( 
.A(n_542),
.B(n_572),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_579),
.B(n_542),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_579),
.B(n_572),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_571),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_553),
.A2(n_590),
.B1(n_577),
.B2(n_607),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_555),
.A2(n_577),
.B(n_569),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_584),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_597),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_600),
.A2(n_604),
.B1(n_607),
.B2(n_563),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_576),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_614),
.B(n_601),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_598),
.A2(n_606),
.B1(n_605),
.B2(n_599),
.Y(n_650)
);

OAI221xp5_ASAP7_75t_SL g651 ( 
.A1(n_561),
.A2(n_558),
.B1(n_619),
.B2(n_563),
.C(n_600),
.Y(n_651)
);

OAI211xp5_ASAP7_75t_L g652 ( 
.A1(n_574),
.A2(n_615),
.B(n_621),
.C(n_604),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_555),
.B(n_609),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_578),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_570),
.A2(n_613),
.B1(n_567),
.B2(n_559),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_620),
.B(n_616),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_616),
.A2(n_622),
.B1(n_594),
.B2(n_570),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_594),
.A2(n_587),
.B1(n_608),
.B2(n_618),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_613),
.Y(n_659)
);

BUFx4f_ASAP7_75t_SL g660 ( 
.A(n_587),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_593),
.Y(n_661)
);

AOI211xp5_ASAP7_75t_L g662 ( 
.A1(n_617),
.A2(n_603),
.B(n_610),
.C(n_611),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_593),
.B(n_568),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_593),
.Y(n_664)
);

OAI221xp5_ASAP7_75t_L g665 ( 
.A1(n_582),
.A2(n_384),
.B1(n_408),
.B2(n_464),
.C(n_434),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_557),
.A2(n_529),
.B1(n_465),
.B2(n_478),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_557),
.A2(n_482),
.B1(n_493),
.B2(n_522),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_557),
.A2(n_529),
.B1(n_465),
.B2(n_478),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_564),
.B(n_513),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_659),
.B(n_625),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_629),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_SL g672 ( 
.A(n_631),
.B(n_652),
.C(n_665),
.Y(n_672)
);

OAI31xp33_ASAP7_75t_L g673 ( 
.A1(n_628),
.A2(n_667),
.A3(n_651),
.B(n_668),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_644),
.A2(n_643),
.B(n_647),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_627),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_625),
.B(n_668),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_632),
.Y(n_677)
);

AOI221xp5_ASAP7_75t_L g678 ( 
.A1(n_624),
.A2(n_666),
.B1(n_669),
.B2(n_636),
.C(n_635),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_623),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_626),
.Y(n_680)
);

OAI221xp5_ASAP7_75t_L g681 ( 
.A1(n_666),
.A2(n_636),
.B1(n_637),
.B2(n_634),
.C(n_649),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_656),
.B(n_654),
.Y(n_682)
);

AO21x2_ASAP7_75t_L g683 ( 
.A1(n_653),
.A2(n_655),
.B(n_650),
.Y(n_683)
);

INVxp67_ASAP7_75t_SL g684 ( 
.A(n_639),
.Y(n_684)
);

AOI211xp5_ASAP7_75t_L g685 ( 
.A1(n_638),
.A2(n_634),
.B(n_641),
.C(n_653),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_646),
.B(n_640),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_661),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_637),
.A2(n_657),
.B1(n_662),
.B2(n_658),
.Y(n_688)
);

OAI221xp5_ASAP7_75t_L g689 ( 
.A1(n_630),
.A2(n_657),
.B1(n_645),
.B2(n_658),
.C(n_664),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_660),
.A2(n_633),
.B1(n_648),
.B2(n_663),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_670),
.B(n_648),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_675),
.Y(n_692)
);

OAI211xp5_ASAP7_75t_L g693 ( 
.A1(n_672),
.A2(n_642),
.B(n_633),
.C(n_648),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_680),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_677),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_679),
.B(n_678),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_680),
.Y(n_697)
);

OAI33xp33_ASAP7_75t_L g698 ( 
.A1(n_688),
.A2(n_633),
.A3(n_648),
.B1(n_686),
.B2(n_682),
.B3(n_670),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_683),
.B(n_676),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_684),
.B(n_687),
.Y(n_700)
);

OAI21xp5_ASAP7_75t_SL g701 ( 
.A1(n_690),
.A2(n_673),
.B(n_676),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_685),
.A2(n_681),
.B1(n_689),
.B2(n_671),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_685),
.B(n_673),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_687),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_699),
.B(n_687),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_694),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_697),
.B(n_677),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_699),
.B(n_677),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_692),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_696),
.B(n_683),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_703),
.B(n_688),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_700),
.B(n_683),
.Y(n_712)
);

AOI211xp5_ASAP7_75t_SL g713 ( 
.A1(n_711),
.A2(n_693),
.B(n_702),
.C(n_701),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_708),
.B(n_695),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_711),
.B(n_683),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_710),
.B(n_700),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_708),
.B(n_691),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_705),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_706),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_707),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_712),
.B(n_700),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_709),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_718),
.B(n_691),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_715),
.B(n_704),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_718),
.A2(n_716),
.B1(n_717),
.B2(n_721),
.Y(n_725)
);

NOR2x1_ASAP7_75t_L g726 ( 
.A(n_719),
.B(n_690),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_SL g727 ( 
.A(n_714),
.B(n_695),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_720),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_714),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_722),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_717),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_730),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_724),
.Y(n_733)
);

NAND3xp33_ASAP7_75t_L g734 ( 
.A(n_727),
.B(n_713),
.C(n_674),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_723),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_725),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_725),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_731),
.Y(n_738)
);

INVxp67_ASAP7_75t_SL g739 ( 
.A(n_726),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_732),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_733),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_736),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_742),
.A2(n_736),
.B1(n_737),
.B2(n_734),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_741),
.B(n_733),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_744),
.Y(n_745)
);

A2O1A1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_745),
.A2(n_743),
.B(n_739),
.C(n_728),
.Y(n_746)
);

OR2x6_ASAP7_75t_L g747 ( 
.A(n_746),
.B(n_735),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_747),
.Y(n_748)
);

NOR2xp67_ASAP7_75t_L g749 ( 
.A(n_747),
.B(n_740),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_748),
.A2(n_738),
.B1(n_740),
.B2(n_735),
.Y(n_750)
);

AOI221xp5_ASAP7_75t_L g751 ( 
.A1(n_750),
.A2(n_749),
.B1(n_698),
.B2(n_732),
.C(n_729),
.Y(n_751)
);


endmodule