module fake_jpeg_17652_n_316 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_20),
.B1(n_21),
.B2(n_32),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_16),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_46),
.B(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_48),
.B(n_27),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_25),
.B1(n_18),
.B2(n_21),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_24),
.B1(n_29),
.B2(n_23),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_36),
.B1(n_32),
.B2(n_18),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_28),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_28),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_24),
.B1(n_29),
.B2(n_3),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_17),
.B1(n_27),
.B2(n_34),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_63),
.B(n_66),
.Y(n_108)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_59),
.B(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_67),
.B(n_97),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_36),
.B1(n_20),
.B2(n_31),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_68),
.A2(n_74),
.B1(n_77),
.B2(n_98),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_38),
.B1(n_46),
.B2(n_25),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_69),
.A2(n_82),
.B1(n_88),
.B2(n_91),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_70),
.A2(n_96),
.B1(n_15),
.B2(n_13),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_71),
.A2(n_33),
.B1(n_30),
.B2(n_12),
.Y(n_113)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_73),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_56),
.B1(n_47),
.B2(n_62),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_1),
.Y(n_128)
);

FAx1_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_45),
.CI(n_42),
.CON(n_76),
.SN(n_76)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_40),
.B(n_55),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_28),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_86),
.Y(n_121)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_60),
.A2(n_53),
.B1(n_50),
.B2(n_62),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_37),
.C(n_44),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_55),
.C(n_19),
.Y(n_110)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_27),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_28),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_45),
.B1(n_42),
.B2(n_41),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_62),
.A2(n_41),
.B1(n_17),
.B2(n_29),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_94),
.B1(n_99),
.B2(n_40),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

BUFx4f_ASAP7_75t_SL g125 ( 
.A(n_90),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_47),
.A2(n_29),
.B1(n_17),
.B2(n_33),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_100),
.B1(n_55),
.B2(n_37),
.Y(n_107)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_54),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_54),
.A2(n_33),
.B1(n_30),
.B2(n_19),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_102),
.A2(n_64),
.B(n_92),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_103),
.A2(n_63),
.B1(n_88),
.B2(n_79),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_106),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_96),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_70),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_114),
.B1(n_127),
.B2(n_88),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_76),
.A2(n_34),
.B1(n_30),
.B2(n_19),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_28),
.C(n_19),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_90),
.C(n_95),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_SL g119 ( 
.A(n_67),
.B(n_34),
.C(n_19),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_124),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_126),
.B1(n_71),
.B2(n_97),
.Y(n_133)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_76),
.A2(n_15),
.B1(n_2),
.B2(n_3),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_76),
.A2(n_82),
.B1(n_83),
.B2(n_65),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_1),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_131),
.A2(n_136),
.B(n_141),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_121),
.B(n_78),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_138),
.C(n_146),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_117),
.B1(n_115),
.B2(n_101),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_116),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_137),
.C(n_142),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_73),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_127),
.A2(n_88),
.B1(n_80),
.B2(n_81),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_144),
.B1(n_148),
.B2(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_122),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_154),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_109),
.B(n_87),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_147),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_121),
.B(n_15),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_109),
.B(n_84),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_64),
.B1(n_72),
.B2(n_94),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_151),
.C(n_156),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_127),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_2),
.C(n_4),
.Y(n_151)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_130),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_153),
.A2(n_113),
.B1(n_105),
.B2(n_104),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_4),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_122),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_SL g182 ( 
.A(n_155),
.B(n_157),
.C(n_6),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_5),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_106),
.B(n_5),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_129),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_161),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_116),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_170),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_102),
.B(n_126),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_165),
.A2(n_171),
.B(n_187),
.Y(n_203)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_157),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_168),
.B(n_185),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_112),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_105),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_120),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_186),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_128),
.B(n_119),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_7),
.B(n_8),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_144),
.B1(n_145),
.B2(n_151),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_101),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_179),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_177),
.A2(n_142),
.B1(n_146),
.B2(n_156),
.Y(n_195)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_178),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_111),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_117),
.B1(n_111),
.B2(n_123),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_125),
.B1(n_7),
.B2(n_8),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_182),
.A2(n_188),
.B1(n_166),
.B2(n_168),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_124),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_187),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_136),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_125),
.C(n_123),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_136),
.B(n_6),
.Y(n_187)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_153),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_193),
.A2(n_199),
.B1(n_205),
.B2(n_214),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_201),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_197),
.B(n_212),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_7),
.B1(n_8),
.B2(n_125),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_200),
.A2(n_166),
.B1(n_159),
.B2(n_182),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_125),
.B(n_178),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_202),
.A2(n_203),
.B(n_206),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_169),
.A2(n_188),
.B1(n_177),
.B2(n_185),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_164),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_210),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_158),
.Y(n_211)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_184),
.C(n_171),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_169),
.B1(n_189),
.B2(n_175),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_180),
.A2(n_174),
.B1(n_179),
.B2(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_181),
.B(n_170),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_216),
.B(n_181),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_162),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_222),
.C(n_226),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_192),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_231),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_171),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_192),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_224),
.B(n_230),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_186),
.C(n_163),
.Y(n_226)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_208),
.B(n_176),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_198),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_196),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_233),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_198),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_163),
.C(n_172),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_239),
.Y(n_249)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_194),
.Y(n_236)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_238),
.A2(n_191),
.B1(n_207),
.B2(n_209),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_195),
.B(n_173),
.C(n_176),
.Y(n_239)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_225),
.B(n_216),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_244),
.B(n_236),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_211),
.Y(n_245)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_210),
.Y(n_246)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g247 ( 
.A(n_239),
.B(n_217),
.CI(n_209),
.CON(n_247),
.SN(n_247)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_247),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_205),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_251),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_237),
.B(n_235),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_202),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_257),
.C(n_237),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_229),
.A2(n_204),
.B1(n_207),
.B2(n_214),
.Y(n_254)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_215),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_228),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_265),
.C(n_269),
.Y(n_286)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_251),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_220),
.Y(n_264)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_222),
.C(n_229),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_233),
.Y(n_268)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_217),
.C(n_221),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_242),
.A2(n_204),
.B(n_223),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_255),
.B1(n_238),
.B2(n_191),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_234),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_256),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_277),
.C(n_263),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_278),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_273),
.Y(n_278)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_272),
.A2(n_271),
.B(n_270),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_280),
.A2(n_283),
.B(n_267),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_200),
.B1(n_196),
.B2(n_247),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_247),
.Y(n_292)
);

O2A1O1Ixp33_ASAP7_75t_SL g287 ( 
.A1(n_266),
.A2(n_254),
.B(n_253),
.C(n_221),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_287),
.A2(n_267),
.B(n_213),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_277),
.B(n_252),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_290),
.Y(n_301)
);

NOR2x1_ASAP7_75t_SL g291 ( 
.A(n_278),
.B(n_268),
.Y(n_291)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_292),
.A3(n_294),
.B1(n_285),
.B2(n_289),
.C1(n_281),
.C2(n_196),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_276),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_269),
.C(n_260),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_286),
.C(n_265),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_298),
.C(n_249),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_260),
.C(n_249),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_282),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_299),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_304),
.B(n_213),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_303),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_287),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_288),
.B(n_261),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_297),
.A2(n_232),
.B(n_275),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_305),
.A2(n_301),
.B(n_298),
.Y(n_311)
);

AOI21xp33_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_308),
.B(n_309),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_311),
.B(n_312),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_193),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_199),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_197),
.C(n_167),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_167),
.Y(n_316)
);


endmodule