module fake_jpeg_10841_n_409 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_409);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_409;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_45),
.B(n_48),
.Y(n_97)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_46),
.Y(n_139)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_47),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g48 ( 
.A(n_23),
.B(n_13),
.C(n_12),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_13),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_50),
.B(n_73),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_51),
.B(n_62),
.Y(n_107)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_57),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_63),
.B(n_65),
.Y(n_131)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_11),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_77),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_25),
.B(n_1),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_88),
.Y(n_101)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

NAND2x1_ASAP7_75t_SL g137 ( 
.A(n_79),
.B(n_80),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_18),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_83),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_20),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_87),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_17),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_90),
.Y(n_98)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_44),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_20),
.B1(n_24),
.B2(n_37),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_93),
.A2(n_95),
.B1(n_109),
.B2(n_25),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_47),
.A2(n_88),
.B1(n_58),
.B2(n_77),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_94),
.A2(n_118),
.B1(n_135),
.B2(n_57),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_20),
.B1(n_24),
.B2(n_37),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_24),
.B1(n_39),
.B2(n_33),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_75),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_110),
.B(n_127),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_115),
.B(n_80),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_58),
.A2(n_44),
.B1(n_42),
.B2(n_36),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_48),
.B(n_39),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_124),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_53),
.B(n_33),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_56),
.B(n_29),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_76),
.B(n_29),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_90),
.A2(n_24),
.B1(n_44),
.B2(n_30),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_130),
.A2(n_134),
.B1(n_30),
.B2(n_21),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_87),
.A2(n_21),
.B1(n_42),
.B2(n_36),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_52),
.A2(n_21),
.B1(n_42),
.B2(n_36),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_72),
.B(n_28),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_79),
.B(n_28),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_137),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_135),
.A2(n_91),
.B1(n_89),
.B2(n_44),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_145),
.A2(n_168),
.B1(n_177),
.B2(n_183),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_146),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_149),
.B(n_173),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_137),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_153),
.B(n_174),
.Y(n_220)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_158),
.A2(n_94),
.B1(n_98),
.B2(n_138),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_SL g226 ( 
.A1(n_159),
.A2(n_138),
.B(n_140),
.Y(n_226)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_161),
.Y(n_219)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_92),
.B(n_22),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_164),
.B(n_176),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_35),
.C(n_60),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_130),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_118),
.A2(n_21),
.B1(n_42),
.B2(n_36),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_172),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_112),
.Y(n_170)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_114),
.Y(n_171)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_46),
.B1(n_30),
.B2(n_79),
.Y(n_175)
);

AO22x1_ASAP7_75t_L g201 ( 
.A1(n_175),
.A2(n_102),
.B1(n_119),
.B2(n_106),
.Y(n_201)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_97),
.A2(n_30),
.B1(n_35),
.B2(n_66),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_189),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_181),
.Y(n_195)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_131),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_184),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_101),
.A2(n_49),
.B1(n_2),
.B2(n_3),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_99),
.B(n_1),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_187),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_188),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_128),
.B(n_4),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_100),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_142),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_194),
.A2(n_197),
.B1(n_206),
.B2(n_208),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_158),
.A2(n_108),
.B1(n_100),
.B2(n_113),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_201),
.A2(n_175),
.B(n_187),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_217),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_159),
.A2(n_108),
.B1(n_125),
.B2(n_134),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_154),
.A2(n_164),
.B1(n_145),
.B2(n_168),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_148),
.A2(n_125),
.B1(n_142),
.B2(n_117),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_213),
.A2(n_226),
.B1(n_102),
.B2(n_175),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_139),
.Y(n_217)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_167),
.A2(n_139),
.B1(n_119),
.B2(n_106),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_152),
.B1(n_157),
.B2(n_147),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_209),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_232),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_180),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_230),
.B(n_254),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_185),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_239),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_221),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_191),
.B(n_179),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_234),
.B(n_241),
.Y(n_271)
);

NOR2x1_ASAP7_75t_L g235 ( 
.A(n_194),
.B(n_171),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_235),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_170),
.B(n_165),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_253),
.Y(n_284)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_240),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_193),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_207),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_247),
.Y(n_276)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_243),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_246),
.B1(n_249),
.B2(n_223),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_208),
.A2(n_184),
.B1(n_176),
.B2(n_173),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_210),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_215),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_259),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_198),
.A2(n_163),
.B1(n_188),
.B2(n_156),
.Y(n_249)
);

NAND2x1p5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_162),
.Y(n_250)
);

AND2x4_ASAP7_75t_L g288 ( 
.A(n_250),
.B(n_199),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_212),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_252),
.B(n_257),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_191),
.A2(n_146),
.B(n_96),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_214),
.B(n_161),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_255),
.A2(n_206),
.B1(n_197),
.B2(n_198),
.Y(n_264)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_256),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_198),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_205),
.Y(n_258)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_192),
.B(n_169),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_203),
.B(n_169),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_219),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_211),
.C(n_223),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_285),
.C(n_287),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_264),
.A2(n_267),
.B1(n_268),
.B2(n_279),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_211),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_266),
.B(n_236),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_201),
.B1(n_216),
.B2(n_212),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_237),
.A2(n_201),
.B1(n_202),
.B2(n_200),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_269),
.A2(n_274),
.B1(n_255),
.B2(n_243),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_236),
.A2(n_200),
.B1(n_225),
.B2(n_202),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_237),
.A2(n_225),
.B1(n_205),
.B2(n_219),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_281),
.B(n_288),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_229),
.A2(n_218),
.B1(n_199),
.B2(n_204),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_289),
.B(n_238),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_204),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_244),
.B(n_218),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_260),
.A2(n_49),
.B1(n_6),
.B2(n_7),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_272),
.A2(n_260),
.B1(n_235),
.B2(n_241),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_272),
.A2(n_235),
.B1(n_254),
.B2(n_250),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_276),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_294),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_234),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_296),
.B(n_297),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_263),
.B(n_242),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_286),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_298),
.B(n_301),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_279),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_299),
.B(n_306),
.Y(n_323)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_300),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_248),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_250),
.C(n_253),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_313),
.C(n_288),
.Y(n_320)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_284),
.A2(n_239),
.B(n_245),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_305),
.A2(n_289),
.B(n_282),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_307),
.Y(n_328)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_308),
.Y(n_333)
);

AND2x6_ASAP7_75t_L g309 ( 
.A(n_261),
.B(n_247),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_309),
.B(n_310),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_266),
.B(n_246),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_231),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_311),
.Y(n_315)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_251),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_240),
.C(n_233),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_302),
.A2(n_265),
.B1(n_284),
.B2(n_288),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_316),
.A2(n_329),
.B1(n_306),
.B2(n_312),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_265),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_311),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_327),
.C(n_330),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_307),
.A2(n_305),
.B1(n_293),
.B2(n_290),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_325),
.A2(n_332),
.B1(n_335),
.B2(n_291),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_326),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_295),
.B(n_303),
.C(n_313),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_302),
.A2(n_288),
.B1(n_264),
.B2(n_268),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_281),
.C(n_278),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_331),
.A2(n_5),
.B(n_6),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_298),
.A2(n_267),
.B1(n_249),
.B2(n_262),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_292),
.A2(n_262),
.B1(n_273),
.B2(n_251),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_337),
.B(n_345),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_325),
.A2(n_314),
.B1(n_294),
.B2(n_299),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_339),
.A2(n_342),
.B1(n_348),
.B2(n_331),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_314),
.C(n_309),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_340),
.B(n_341),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_308),
.C(n_300),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_320),
.B(n_330),
.C(n_316),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_344),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_317),
.B(n_304),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_310),
.C(n_258),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_324),
.Y(n_346)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_346),
.Y(n_357)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_334),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_349),
.Y(n_365)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_318),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_350),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_351),
.A2(n_345),
.B1(n_328),
.B2(n_315),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_336),
.B(n_273),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_323),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_353),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_355),
.A2(n_368),
.B1(n_354),
.B2(n_343),
.Y(n_372)
);

INVx13_ASAP7_75t_L g356 ( 
.A(n_354),
.Y(n_356)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_356),
.Y(n_370)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_341),
.Y(n_362)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_362),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_340),
.A2(n_328),
.B1(n_323),
.B2(n_335),
.Y(n_364)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_364),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_367),
.B(n_337),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_372),
.A2(n_375),
.B1(n_360),
.B2(n_364),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_374),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_362),
.B(n_338),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_368),
.A2(n_318),
.B1(n_333),
.B2(n_321),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_338),
.C(n_329),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_377),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_321),
.C(n_333),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_359),
.B(n_5),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_378),
.B(n_369),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_365),
.Y(n_381)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_381),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_382),
.A2(n_383),
.B1(n_380),
.B2(n_370),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_380),
.A2(n_357),
.B1(n_361),
.B2(n_363),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_366),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_5),
.Y(n_394)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_386),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_369),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_387),
.A2(n_389),
.B(n_363),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_376),
.B(n_367),
.C(n_356),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_391),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_379),
.C(n_372),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_392),
.A2(n_394),
.B(n_395),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_384),
.B(n_5),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_393),
.A2(n_381),
.B(n_389),
.Y(n_399)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_399),
.Y(n_403)
);

AOI21x1_ASAP7_75t_L g400 ( 
.A1(n_391),
.A2(n_388),
.B(n_8),
.Y(n_400)
);

AO221x1_ASAP7_75t_L g402 ( 
.A1(n_400),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.C(n_394),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_397),
.B(n_396),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_401),
.Y(n_404)
);

O2A1O1Ixp33_ASAP7_75t_SL g405 ( 
.A1(n_402),
.A2(n_398),
.B(n_8),
.C(n_9),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_405),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_403),
.C(n_404),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_407),
.B(n_7),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_9),
.Y(n_409)
);


endmodule