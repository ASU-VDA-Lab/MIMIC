module fake_jpeg_25746_n_166 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_166);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

CKINVDCx6p67_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_25),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_27),
.Y(n_53)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_53),
.Y(n_58)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_22),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_38),
.B1(n_37),
.B2(n_30),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_54),
.B1(n_37),
.B2(n_38),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_29),
.B1(n_20),
.B2(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_24),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_65),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_14),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_18),
.B1(n_28),
.B2(n_19),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_72),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_15),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_27),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_31),
.C(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_32),
.Y(n_85)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_14),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_78),
.B(n_82),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_74),
.A2(n_44),
.B1(n_34),
.B2(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_86),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_59),
.B(n_23),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_73),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_33),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_33),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_23),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_58),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_44),
.B1(n_48),
.B2(n_56),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_65),
.B1(n_67),
.B2(n_75),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_93),
.B1(n_48),
.B2(n_24),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_48),
.B1(n_28),
.B2(n_19),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_94),
.B(n_95),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_101),
.Y(n_110)
);

BUFx4f_ASAP7_75t_SL g99 ( 
.A(n_81),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_77),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_100),
.B(n_108),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_62),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_105),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_66),
.B1(n_18),
.B2(n_16),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_80),
.B1(n_84),
.B2(n_92),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_87),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_42),
.C(n_39),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_84),
.C(n_42),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_122),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_82),
.Y(n_117)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_102),
.B1(n_94),
.B2(n_114),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_107),
.C(n_92),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_78),
.B(n_76),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_9),
.B(n_12),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_60),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_127),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_101),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_130),
.C(n_39),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_135),
.B(n_0),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_91),
.B1(n_76),
.B2(n_109),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_133),
.B1(n_121),
.B2(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_99),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_119),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_134),
.B(n_112),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_99),
.B(n_60),
.C(n_39),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_1),
.Y(n_149)
);

NAND2x1_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_118),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_137),
.A2(n_138),
.B(n_142),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_112),
.B1(n_110),
.B2(n_118),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_141),
.B(n_144),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_130),
.C(n_135),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_137),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_135),
.C(n_128),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_148),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_124),
.C(n_10),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_2),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_154),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

OAI221xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.C(n_154),
.Y(n_159)
);

O2A1O1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_145),
.A2(n_137),
.B(n_144),
.C(n_136),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_156),
.B(n_2),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_158),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_155),
.A2(n_151),
.B(n_8),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_156),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_3),
.C(n_5),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_162),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_163),
.Y(n_166)
);


endmodule