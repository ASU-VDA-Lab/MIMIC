module fake_jpeg_12165_n_104 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_13),
.B(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_51),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_39),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_34),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_60),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_37),
.B1(n_39),
.B2(n_29),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_61),
.A2(n_42),
.B(n_36),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_29),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_37),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_1),
.B(n_2),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_74),
.Y(n_83)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_31),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_70),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_61),
.B(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_64),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_10),
.B1(n_12),
.B2(n_16),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_18),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_76),
.B(n_8),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_3),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_84),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_85),
.B1(n_26),
.B2(n_28),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_86),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_17),
.C(n_20),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_91),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_21),
.B(n_22),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_23),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_93),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_94),
.C(n_90),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_87),
.Y(n_100)
);

AOI21x1_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_90),
.B(n_95),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_89),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_77),
.Y(n_104)
);


endmodule