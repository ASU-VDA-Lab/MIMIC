module fake_jpeg_24122_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx16_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_24),
.Y(n_35)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_26),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_14),
.B(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_2),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_28),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_2),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_36),
.B(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_19),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_34),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_24),
.B1(n_21),
.B2(n_12),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_41),
.B1(n_43),
.B2(n_30),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_10),
.B1(n_20),
.B2(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_29),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_55),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_51),
.B(n_53),
.Y(n_61)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_56),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_43),
.B(n_13),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_59),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_50),
.B(n_39),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_44),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_60),
.Y(n_67)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_63),
.A2(n_66),
.B1(n_30),
.B2(n_54),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_43),
.B1(n_16),
.B2(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_70),
.B(n_20),
.C(n_6),
.Y(n_74)
);

BUFx24_ASAP7_75t_SL g73 ( 
.A(n_72),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_74),
.B(n_16),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_18),
.A3(n_52),
.B1(n_5),
.B2(n_6),
.C1(n_47),
.C2(n_46),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_5),
.Y(n_77)
);


endmodule