module fake_jpeg_30381_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_20),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_9),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_76),
.Y(n_83)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_0),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_66),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_56),
.Y(n_78)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_69),
.B(n_59),
.C(n_63),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_89),
.B(n_52),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_50),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_67),
.B1(n_66),
.B2(n_60),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_92),
.B1(n_53),
.B2(n_25),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_68),
.B1(n_64),
.B2(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_53),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_67),
.B1(n_60),
.B2(n_68),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_101),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_55),
.Y(n_96)
);

FAx1_ASAP7_75t_SL g121 ( 
.A(n_96),
.B(n_99),
.CI(n_4),
.CON(n_121),
.SN(n_121)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_77),
.B1(n_72),
.B2(n_78),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_85),
.B1(n_84),
.B2(n_80),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_89),
.B1(n_52),
.B2(n_93),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_28),
.B1(n_46),
.B2(n_45),
.Y(n_120)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_51),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_106),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_0),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_12),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_2),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_2),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_84),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_119),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_125),
.B1(n_35),
.B2(n_36),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_128),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_107),
.B1(n_95),
.B2(n_102),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_6),
.B(n_7),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_129),
.B(n_27),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_18),
.C(n_19),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_13),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_13),
.B(n_16),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_17),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_130),
.B(n_32),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_133),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_111),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_143),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_113),
.B(n_22),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_23),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_129),
.C(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_137),
.B(n_145),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_123),
.A2(n_30),
.B(n_31),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_138),
.B(n_140),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_34),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_126),
.B(n_37),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_144),
.Y(n_146)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_131),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_139),
.B(n_136),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_153),
.A2(n_148),
.B1(n_142),
.B2(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_155),
.Y(n_156)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_141),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_156),
.B(n_148),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_147),
.B(n_134),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_146),
.C(n_151),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_38),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_48),
.Y(n_164)
);


endmodule