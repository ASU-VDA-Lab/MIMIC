module real_aes_8216_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g465 ( .A1(n_0), .A2(n_166), .B(n_466), .C(n_469), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_1), .B(n_460), .Y(n_471) );
INVx1_ASAP7_75t_L g429 ( .A(n_2), .Y(n_429) );
INVx1_ASAP7_75t_L g215 ( .A(n_3), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_4), .B(n_154), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_5), .A2(n_444), .B(n_514), .Y(n_513) );
OAI22xp5_ASAP7_75t_SL g753 ( .A1(n_6), .A2(n_9), .B1(n_424), .B2(n_754), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_6), .Y(n_754) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_7), .A2(n_171), .B(n_523), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_8), .A2(n_39), .B1(n_127), .B2(n_139), .Y(n_165) );
AOI22xp5_ASAP7_75t_L g110 ( .A1(n_9), .A2(n_111), .B1(n_112), .B2(n_424), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_9), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_10), .B(n_171), .Y(n_204) );
AND2x6_ASAP7_75t_L g142 ( .A(n_11), .B(n_143), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_12), .A2(n_142), .B(n_447), .C(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_13), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_14), .B(n_40), .Y(n_430) );
INVx1_ASAP7_75t_L g123 ( .A(n_15), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_16), .B(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g209 ( .A(n_17), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_18), .B(n_154), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_19), .B(n_169), .Y(n_187) );
AO32x2_ASAP7_75t_L g163 ( .A1(n_20), .A2(n_164), .A3(n_168), .B1(n_170), .B2(n_171), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g104 ( .A1(n_21), .A2(n_99), .B1(n_105), .B2(n_106), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_21), .Y(n_106) );
AND2x2_ASAP7_75t_L g508 ( .A(n_22), .B(n_119), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_23), .B(n_127), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_24), .B(n_169), .Y(n_217) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_25), .A2(n_55), .B1(n_127), .B2(n_139), .Y(n_167) );
AOI22xp33_ASAP7_75t_SL g180 ( .A1(n_26), .A2(n_81), .B1(n_127), .B2(n_131), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_27), .B(n_127), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_28), .A2(n_170), .B(n_447), .C(n_449), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_29), .A2(n_170), .B(n_447), .C(n_526), .Y(n_525) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_30), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_31), .B(n_119), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_32), .A2(n_444), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_33), .B(n_119), .Y(n_161) );
INVx2_ASAP7_75t_L g129 ( .A(n_34), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_35), .A2(n_478), .B(n_479), .C(n_483), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_36), .B(n_127), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_37), .B(n_119), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_38), .B(n_134), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_41), .B(n_443), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_42), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_43), .B(n_154), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_44), .B(n_444), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_45), .A2(n_478), .B(n_483), .C(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_46), .B(n_127), .Y(n_197) );
INVx1_ASAP7_75t_L g467 ( .A(n_47), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_48), .B(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_49), .A2(n_89), .B1(n_139), .B2(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g506 ( .A(n_50), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_51), .B(n_127), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_52), .B(n_127), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_53), .B(n_444), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_54), .B(n_202), .Y(n_201) );
AOI22xp33_ASAP7_75t_SL g191 ( .A1(n_56), .A2(n_60), .B1(n_127), .B2(n_131), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_57), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_58), .B(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_59), .B(n_127), .Y(n_228) );
INVx1_ASAP7_75t_L g143 ( .A(n_61), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_62), .B(n_444), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_63), .B(n_460), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_64), .A2(n_202), .B(n_212), .C(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_65), .B(n_127), .Y(n_216) );
INVx1_ASAP7_75t_L g122 ( .A(n_66), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_67), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_68), .B(n_154), .Y(n_481) );
AO32x2_ASAP7_75t_L g176 ( .A1(n_69), .A2(n_170), .A3(n_171), .B1(n_177), .B2(n_181), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_70), .B(n_155), .Y(n_537) );
INVx1_ASAP7_75t_L g227 ( .A(n_71), .Y(n_227) );
INVx1_ASAP7_75t_L g152 ( .A(n_72), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g463 ( .A(n_73), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_74), .B(n_451), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_75), .A2(n_447), .B(n_483), .C(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_76), .B(n_751), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_76), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_76), .B(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_77), .B(n_131), .Y(n_153) );
CKINVDCx16_ASAP7_75t_R g515 ( .A(n_78), .Y(n_515) );
INVx1_ASAP7_75t_L g739 ( .A(n_79), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_80), .B(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_82), .B(n_139), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_83), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_84), .B(n_131), .Y(n_158) );
INVx2_ASAP7_75t_L g120 ( .A(n_85), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_86), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_87), .B(n_141), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_88), .B(n_131), .Y(n_198) );
OR2x2_ASAP7_75t_L g427 ( .A(n_90), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g725 ( .A(n_90), .Y(n_725) );
OR2x2_ASAP7_75t_L g743 ( .A(n_90), .B(n_734), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_91), .A2(n_100), .B1(n_131), .B2(n_132), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_92), .B(n_444), .Y(n_476) );
INVx1_ASAP7_75t_L g480 ( .A(n_93), .Y(n_480) );
INVxp67_ASAP7_75t_L g518 ( .A(n_94), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_95), .B(n_131), .Y(n_225) );
INVx1_ASAP7_75t_L g493 ( .A(n_96), .Y(n_493) );
INVx1_ASAP7_75t_L g533 ( .A(n_97), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_98), .B(n_739), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_99), .Y(n_105) );
O2A1O1Ixp33_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_730), .B(n_735), .C(n_744), .Y(n_101) );
HB1xp67_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_107), .B1(n_726), .B2(n_727), .Y(n_103) );
INVx1_ASAP7_75t_L g726 ( .A(n_104), .Y(n_726) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OAI22x1_ASAP7_75t_SL g108 ( .A1(n_109), .A2(n_425), .B1(n_431), .B2(n_722), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_110), .A2(n_432), .B1(n_722), .B2(n_729), .Y(n_728) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_111), .A2(n_112), .B1(n_752), .B2(n_753), .Y(n_751) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_346), .Y(n_112) );
NAND5xp2_ASAP7_75t_L g113 ( .A(n_114), .B(n_265), .C(n_280), .D(n_306), .E(n_328), .Y(n_113) );
NOR2xp33_ASAP7_75t_SL g114 ( .A(n_115), .B(n_245), .Y(n_114) );
OAI221xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_182), .B1(n_218), .B2(n_234), .C(n_235), .Y(n_115) );
NOR2xp33_ASAP7_75t_SL g116 ( .A(n_117), .B(n_172), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_117), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_SL g422 ( .A(n_117), .Y(n_422) );
AND2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_145), .Y(n_117) );
INVx1_ASAP7_75t_L g262 ( .A(n_118), .Y(n_262) );
AND2x2_ASAP7_75t_L g264 ( .A(n_118), .B(n_163), .Y(n_264) );
AND2x2_ASAP7_75t_L g274 ( .A(n_118), .B(n_162), .Y(n_274) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_118), .Y(n_292) );
INVx1_ASAP7_75t_L g302 ( .A(n_118), .Y(n_302) );
OR2x2_ASAP7_75t_L g340 ( .A(n_118), .B(n_239), .Y(n_340) );
INVx2_ASAP7_75t_L g390 ( .A(n_118), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_118), .B(n_238), .Y(n_407) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_144), .Y(n_118) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_119), .A2(n_149), .B(n_161), .Y(n_148) );
INVx2_ASAP7_75t_L g181 ( .A(n_119), .Y(n_181) );
INVx1_ASAP7_75t_L g457 ( .A(n_119), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_119), .A2(n_476), .B(n_477), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_119), .A2(n_503), .B(n_504), .Y(n_502) );
AND2x2_ASAP7_75t_SL g119 ( .A(n_120), .B(n_121), .Y(n_119) );
AND2x2_ASAP7_75t_L g169 ( .A(n_120), .B(n_121), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
OAI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_136), .B(n_142), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_130), .B(n_133), .Y(n_125) );
INVx3_ASAP7_75t_L g151 ( .A(n_127), .Y(n_151) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_127), .Y(n_495) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g139 ( .A(n_128), .Y(n_139) );
BUFx3_ASAP7_75t_L g179 ( .A(n_128), .Y(n_179) );
AND2x6_ASAP7_75t_L g447 ( .A(n_128), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g132 ( .A(n_129), .Y(n_132) );
INVx1_ASAP7_75t_L g203 ( .A(n_129), .Y(n_203) );
INVx2_ASAP7_75t_L g210 ( .A(n_131), .Y(n_210) );
INVx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
INVx3_ASAP7_75t_L g155 ( .A(n_135), .Y(n_155) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_135), .Y(n_160) );
AND2x2_ASAP7_75t_L g445 ( .A(n_135), .B(n_203), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_135), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B(n_140), .Y(n_136) );
O2A1O1Ixp5_ASAP7_75t_L g226 ( .A1(n_140), .A2(n_214), .B(n_227), .C(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g164 ( .A1(n_141), .A2(n_165), .B1(n_166), .B2(n_167), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g177 ( .A1(n_141), .A2(n_155), .B1(n_178), .B2(n_180), .Y(n_177) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_141), .A2(n_166), .B1(n_190), .B2(n_191), .Y(n_189) );
INVx4_ASAP7_75t_L g468 ( .A(n_141), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g149 ( .A1(n_142), .A2(n_150), .B(n_156), .Y(n_149) );
BUFx3_ASAP7_75t_L g170 ( .A(n_142), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g195 ( .A1(n_142), .A2(n_196), .B(n_199), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_142), .A2(n_208), .B(n_213), .Y(n_207) );
AND2x4_ASAP7_75t_L g444 ( .A(n_142), .B(n_445), .Y(n_444) );
INVx4_ASAP7_75t_SL g470 ( .A(n_142), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g534 ( .A(n_142), .B(n_445), .Y(n_534) );
NOR2xp67_ASAP7_75t_L g145 ( .A(n_146), .B(n_162), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_147), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_147), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_SL g322 ( .A(n_147), .B(n_262), .Y(n_322) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_148), .Y(n_174) );
INVx2_ASAP7_75t_L g239 ( .A(n_148), .Y(n_239) );
OR2x2_ASAP7_75t_L g301 ( .A(n_148), .B(n_302), .Y(n_301) );
O2A1O1Ixp5_ASAP7_75t_SL g150 ( .A1(n_151), .A2(n_152), .B(n_153), .C(n_154), .Y(n_150) );
INVx2_ASAP7_75t_L g166 ( .A(n_154), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_154), .A2(n_197), .B(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_154), .A2(n_224), .B(n_225), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_154), .B(n_518), .Y(n_517) );
INVx5_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_159), .Y(n_156) );
INVx1_ASAP7_75t_L g212 ( .A(n_159), .Y(n_212) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g451 ( .A(n_160), .Y(n_451) );
AND2x2_ASAP7_75t_L g240 ( .A(n_162), .B(n_176), .Y(n_240) );
AND2x2_ASAP7_75t_L g257 ( .A(n_162), .B(n_237), .Y(n_257) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g175 ( .A(n_163), .B(n_176), .Y(n_175) );
BUFx2_ASAP7_75t_L g260 ( .A(n_163), .Y(n_260) );
AND2x2_ASAP7_75t_L g389 ( .A(n_163), .B(n_390), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_166), .A2(n_200), .B(n_201), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_166), .A2(n_214), .B(n_215), .C(n_216), .Y(n_213) );
INVx2_ASAP7_75t_L g206 ( .A(n_168), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_168), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_169), .Y(n_171) );
NAND3xp33_ASAP7_75t_L g188 ( .A(n_170), .B(n_189), .C(n_192), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_170), .A2(n_223), .B(n_226), .Y(n_222) );
INVx4_ASAP7_75t_L g192 ( .A(n_171), .Y(n_192) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_171), .A2(n_195), .B(n_204), .Y(n_194) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_171), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_171), .A2(n_524), .B(n_525), .Y(n_523) );
INVx1_ASAP7_75t_L g234 ( .A(n_172), .Y(n_234) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_175), .Y(n_172) );
AND2x2_ASAP7_75t_L g352 ( .A(n_173), .B(n_240), .Y(n_352) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g353 ( .A(n_174), .B(n_264), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_L g320 ( .A1(n_175), .A2(n_321), .B(n_323), .C(n_325), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_175), .B(n_321), .Y(n_330) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_175), .A2(n_251), .B1(n_394), .B2(n_395), .C(n_397), .Y(n_393) );
INVx1_ASAP7_75t_L g237 ( .A(n_176), .Y(n_237) );
INVx1_ASAP7_75t_L g273 ( .A(n_176), .Y(n_273) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_176), .Y(n_282) );
INVx2_ASAP7_75t_L g469 ( .A(n_179), .Y(n_469) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_179), .Y(n_482) );
INVx1_ASAP7_75t_L g454 ( .A(n_181), .Y(n_454) );
INVx1_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_193), .Y(n_183) );
AND2x2_ASAP7_75t_L g299 ( .A(n_184), .B(n_244), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_184), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_185), .B(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g391 ( .A(n_185), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g423 ( .A(n_185), .Y(n_423) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx3_ASAP7_75t_L g253 ( .A(n_186), .Y(n_253) );
AND2x2_ASAP7_75t_L g279 ( .A(n_186), .B(n_233), .Y(n_279) );
NOR2x1_ASAP7_75t_L g288 ( .A(n_186), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g295 ( .A(n_186), .B(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
INVx1_ASAP7_75t_L g231 ( .A(n_187), .Y(n_231) );
AO21x1_ASAP7_75t_L g230 ( .A1(n_189), .A2(n_192), .B(n_231), .Y(n_230) );
INVx3_ASAP7_75t_L g460 ( .A(n_192), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_192), .B(n_485), .Y(n_484) );
AO21x2_ASAP7_75t_L g489 ( .A1(n_192), .A2(n_490), .B(n_497), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_192), .B(n_498), .Y(n_497) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_192), .A2(n_532), .B(n_539), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_193), .B(n_335), .Y(n_370) );
INVx1_ASAP7_75t_SL g374 ( .A(n_193), .Y(n_374) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_205), .Y(n_193) );
INVx3_ASAP7_75t_L g233 ( .A(n_194), .Y(n_233) );
AND2x2_ASAP7_75t_L g244 ( .A(n_194), .B(n_221), .Y(n_244) );
AND2x2_ASAP7_75t_L g266 ( .A(n_194), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g311 ( .A(n_194), .B(n_305), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_194), .B(n_243), .Y(n_392) );
INVx2_ASAP7_75t_L g214 ( .A(n_202), .Y(n_214) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g232 ( .A(n_205), .B(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g243 ( .A(n_205), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_205), .B(n_221), .Y(n_268) );
AND2x2_ASAP7_75t_L g304 ( .A(n_205), .B(n_305), .Y(n_304) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_217), .Y(n_205) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_206), .A2(n_222), .B(n_229), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_211), .C(n_212), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_210), .A2(n_527), .B(n_528), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_210), .A2(n_537), .B(n_538), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_212), .A2(n_493), .B(n_494), .C(n_495), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_214), .A2(n_450), .B(n_452), .Y(n_449) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_232), .Y(n_219) );
INVx1_ASAP7_75t_L g284 ( .A(n_220), .Y(n_284) );
AND2x2_ASAP7_75t_L g326 ( .A(n_220), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_220), .B(n_247), .Y(n_332) );
AOI21xp5_ASAP7_75t_SL g406 ( .A1(n_220), .A2(n_238), .B(n_261), .Y(n_406) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_230), .Y(n_220) );
OR2x2_ASAP7_75t_L g249 ( .A(n_221), .B(n_230), .Y(n_249) );
AND2x2_ASAP7_75t_L g296 ( .A(n_221), .B(n_233), .Y(n_296) );
INVx2_ASAP7_75t_L g305 ( .A(n_221), .Y(n_305) );
INVx1_ASAP7_75t_L g411 ( .A(n_221), .Y(n_411) );
AND2x2_ASAP7_75t_L g335 ( .A(n_230), .B(n_305), .Y(n_335) );
INVx1_ASAP7_75t_L g360 ( .A(n_230), .Y(n_360) );
AND2x2_ASAP7_75t_L g269 ( .A(n_232), .B(n_253), .Y(n_269) );
AND2x2_ASAP7_75t_L g281 ( .A(n_232), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_SL g399 ( .A(n_232), .Y(n_399) );
INVx2_ASAP7_75t_L g289 ( .A(n_233), .Y(n_289) );
AND2x2_ASAP7_75t_L g327 ( .A(n_233), .B(n_243), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_233), .B(n_411), .Y(n_410) );
OAI21xp33_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_240), .B(n_241), .Y(n_235) );
AND2x2_ASAP7_75t_L g342 ( .A(n_236), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g396 ( .A(n_236), .Y(n_396) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx1_ASAP7_75t_L g316 ( .A(n_237), .Y(n_316) );
BUFx2_ASAP7_75t_L g415 ( .A(n_237), .Y(n_415) );
BUFx2_ASAP7_75t_L g286 ( .A(n_238), .Y(n_286) );
AND2x2_ASAP7_75t_L g388 ( .A(n_238), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g371 ( .A(n_239), .Y(n_371) );
AND2x4_ASAP7_75t_L g298 ( .A(n_240), .B(n_261), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_240), .B(n_322), .Y(n_334) );
AOI32xp33_ASAP7_75t_L g258 ( .A1(n_241), .A2(n_259), .A3(n_261), .B1(n_263), .B2(n_264), .Y(n_258) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
INVx3_ASAP7_75t_L g247 ( .A(n_242), .Y(n_247) );
OR2x2_ASAP7_75t_L g383 ( .A(n_242), .B(n_339), .Y(n_383) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g252 ( .A(n_243), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g359 ( .A(n_243), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g251 ( .A(n_244), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g263 ( .A(n_244), .B(n_253), .Y(n_263) );
INVx1_ASAP7_75t_L g384 ( .A(n_244), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_244), .B(n_359), .Y(n_417) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_250), .B(n_254), .C(n_258), .Y(n_245) );
OAI322xp33_ASAP7_75t_L g354 ( .A1(n_246), .A2(n_291), .A3(n_355), .B1(n_357), .B2(n_361), .C1(n_362), .C2(n_366), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVxp67_ASAP7_75t_L g319 ( .A(n_247), .Y(n_319) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g373 ( .A(n_249), .B(n_374), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_249), .B(n_289), .Y(n_420) );
INVxp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g312 ( .A(n_252), .Y(n_312) );
OR2x2_ASAP7_75t_L g398 ( .A(n_253), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_256), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g307 ( .A(n_257), .B(n_286), .Y(n_307) );
AND2x2_ASAP7_75t_L g378 ( .A(n_257), .B(n_291), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_257), .B(n_365), .Y(n_400) );
AOI221xp5_ASAP7_75t_L g265 ( .A1(n_259), .A2(n_266), .B1(n_269), .B2(n_270), .C(n_275), .Y(n_265) );
OR2x2_ASAP7_75t_L g276 ( .A(n_259), .B(n_272), .Y(n_276) );
AND2x2_ASAP7_75t_L g364 ( .A(n_259), .B(n_365), .Y(n_364) );
AOI32xp33_ASAP7_75t_L g403 ( .A1(n_259), .A2(n_289), .A3(n_404), .B1(n_405), .B2(n_408), .Y(n_403) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND3xp33_ASAP7_75t_L g337 ( .A(n_260), .B(n_296), .C(n_319), .Y(n_337) );
AND2x2_ASAP7_75t_L g363 ( .A(n_260), .B(n_356), .Y(n_363) );
INVxp67_ASAP7_75t_L g343 ( .A(n_261), .Y(n_343) );
BUFx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_264), .B(n_316), .Y(n_372) );
INVx2_ASAP7_75t_L g382 ( .A(n_264), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_264), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g351 ( .A(n_267), .Y(n_351) );
OR2x2_ASAP7_75t_L g277 ( .A(n_268), .B(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_270), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_274), .Y(n_270) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_273), .Y(n_356) );
AND2x2_ASAP7_75t_L g315 ( .A(n_274), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g361 ( .A(n_274), .Y(n_361) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_274), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
AOI21xp33_ASAP7_75t_SL g300 ( .A1(n_276), .A2(n_301), .B(n_303), .Y(n_300) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g394 ( .A(n_279), .B(n_304), .Y(n_394) );
AOI211xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_283), .B(n_293), .C(n_300), .Y(n_280) );
AND2x2_ASAP7_75t_L g324 ( .A(n_282), .B(n_292), .Y(n_324) );
INVx2_ASAP7_75t_L g339 ( .A(n_282), .Y(n_339) );
OR2x2_ASAP7_75t_L g377 ( .A(n_282), .B(n_340), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_282), .B(n_420), .Y(n_419) );
AOI211xp5_ASAP7_75t_SL g283 ( .A1(n_284), .A2(n_285), .B(n_287), .C(n_290), .Y(n_283) );
INVxp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_286), .B(n_324), .Y(n_323) );
OAI211xp5_ASAP7_75t_L g405 ( .A1(n_287), .A2(n_382), .B(n_406), .C(n_407), .Y(n_405) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2x1p5_ASAP7_75t_L g303 ( .A(n_288), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g345 ( .A(n_289), .B(n_335), .Y(n_345) );
INVx1_ASAP7_75t_L g350 ( .A(n_289), .Y(n_350) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_294), .B(n_297), .Y(n_293) );
INVxp33_ASAP7_75t_L g401 ( .A(n_295), .Y(n_401) );
AND2x2_ASAP7_75t_L g380 ( .A(n_296), .B(n_359), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_301), .A2(n_363), .B(n_364), .Y(n_362) );
OAI322xp33_ASAP7_75t_L g381 ( .A1(n_303), .A2(n_382), .A3(n_383), .B1(n_384), .B2(n_385), .C1(n_387), .C2(n_391), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B1(n_313), .B2(n_317), .C(n_320), .Y(n_306) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g358 ( .A(n_311), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g402 ( .A(n_315), .Y(n_402) );
INVxp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_318), .B(n_338), .Y(n_404) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g367 ( .A(n_327), .B(n_335), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .B1(n_333), .B2(n_335), .C(n_336), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_331), .A2(n_348), .B1(n_352), .B2(n_353), .C(n_354), .Y(n_347) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVxp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_335), .B(n_350), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B1(n_341), .B2(n_344), .Y(n_336) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx2_ASAP7_75t_SL g365 ( .A(n_340), .Y(n_365) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND5xp2_ASAP7_75t_L g346 ( .A(n_347), .B(n_368), .C(n_393), .D(n_403), .E(n_413), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_349), .B(n_351), .Y(n_348) );
NOR4xp25_ASAP7_75t_L g421 ( .A(n_350), .B(n_356), .C(n_422), .D(n_423), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_353), .A2(n_414), .B1(n_416), .B2(n_418), .C(n_421), .Y(n_413) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g412 ( .A(n_359), .Y(n_412) );
OAI322xp33_ASAP7_75t_L g369 ( .A1(n_363), .A2(n_370), .A3(n_371), .B1(n_372), .B2(n_373), .C1(n_375), .C2(n_379), .Y(n_369) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_369), .B(n_381), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g414 ( .A(n_389), .B(n_415), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B1(n_401), .B2(n_402), .Y(n_397) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g729 ( .A(n_426), .Y(n_729) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g724 ( .A(n_428), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g734 ( .A(n_428), .Y(n_734) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_SL g432 ( .A(n_433), .B(n_677), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_612), .Y(n_433) );
NAND4xp25_ASAP7_75t_SL g434 ( .A(n_435), .B(n_557), .C(n_581), .D(n_604), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_499), .B1(n_529), .B2(n_541), .C(n_544), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_472), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_438), .A2(n_458), .B1(n_500), .B2(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_438), .B(n_473), .Y(n_615) );
AND2x2_ASAP7_75t_L g634 ( .A(n_438), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_438), .B(n_618), .Y(n_704) );
AND2x4_ASAP7_75t_L g438 ( .A(n_439), .B(n_458), .Y(n_438) );
AND2x2_ASAP7_75t_L g572 ( .A(n_439), .B(n_473), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_439), .B(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g595 ( .A(n_439), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g600 ( .A(n_439), .B(n_459), .Y(n_600) );
INVx2_ASAP7_75t_L g632 ( .A(n_439), .Y(n_632) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_439), .Y(n_676) );
AND2x2_ASAP7_75t_L g693 ( .A(n_439), .B(n_570), .Y(n_693) );
INVx5_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g611 ( .A(n_440), .B(n_570), .Y(n_611) );
AND2x4_ASAP7_75t_L g625 ( .A(n_440), .B(n_458), .Y(n_625) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_440), .Y(n_629) );
AND2x2_ASAP7_75t_L g649 ( .A(n_440), .B(n_564), .Y(n_649) );
AND2x2_ASAP7_75t_L g699 ( .A(n_440), .B(n_474), .Y(n_699) );
AND2x2_ASAP7_75t_L g709 ( .A(n_440), .B(n_459), .Y(n_709) );
OR2x6_ASAP7_75t_L g440 ( .A(n_441), .B(n_455), .Y(n_440) );
AOI21xp5_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_446), .B(n_454), .Y(n_441) );
BUFx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx5_ASAP7_75t_L g464 ( .A(n_447), .Y(n_464) );
INVx2_ASAP7_75t_L g453 ( .A(n_451), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_453), .A2(n_480), .B(n_481), .C(n_482), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_453), .A2(n_482), .B(n_506), .C(n_507), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
AND2x2_ASAP7_75t_L g565 ( .A(n_458), .B(n_473), .Y(n_565) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_458), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_458), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g655 ( .A(n_458), .Y(n_655) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g543 ( .A(n_459), .B(n_488), .Y(n_543) );
AND2x2_ASAP7_75t_L g570 ( .A(n_459), .B(n_489), .Y(n_570) );
OA21x2_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B(n_471), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_464), .B(n_465), .C(n_470), .Y(n_462) );
INVx2_ASAP7_75t_L g478 ( .A(n_464), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_464), .A2(n_470), .B(n_515), .C(n_516), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVx1_ASAP7_75t_L g483 ( .A(n_470), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_472), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_486), .Y(n_472) );
OR2x2_ASAP7_75t_L g596 ( .A(n_473), .B(n_487), .Y(n_596) );
AND2x2_ASAP7_75t_L g633 ( .A(n_473), .B(n_543), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_473), .B(n_564), .Y(n_644) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_473), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_473), .B(n_600), .Y(n_717) );
INVx5_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g542 ( .A(n_474), .Y(n_542) );
AND2x2_ASAP7_75t_L g551 ( .A(n_474), .B(n_487), .Y(n_551) );
AND2x2_ASAP7_75t_L g667 ( .A(n_474), .B(n_562), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_474), .B(n_600), .Y(n_689) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_487), .Y(n_635) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_488), .Y(n_587) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g564 ( .A(n_489), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_496), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_509), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_500), .B(n_577), .Y(n_696) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_501), .B(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g548 ( .A(n_501), .B(n_549), .Y(n_548) );
INVx5_ASAP7_75t_SL g556 ( .A(n_501), .Y(n_556) );
OR2x2_ASAP7_75t_L g579 ( .A(n_501), .B(n_549), .Y(n_579) );
OR2x2_ASAP7_75t_L g589 ( .A(n_501), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g652 ( .A(n_501), .B(n_511), .Y(n_652) );
AND2x2_ASAP7_75t_SL g690 ( .A(n_501), .B(n_510), .Y(n_690) );
NOR4xp25_ASAP7_75t_L g711 ( .A(n_501), .B(n_632), .C(n_712), .D(n_713), .Y(n_711) );
AND2x2_ASAP7_75t_L g721 ( .A(n_501), .B(n_553), .Y(n_721) );
OR2x6_ASAP7_75t_L g501 ( .A(n_502), .B(n_508), .Y(n_501) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g546 ( .A(n_510), .B(n_542), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_510), .B(n_548), .Y(n_715) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_520), .Y(n_510) );
OR2x2_ASAP7_75t_L g555 ( .A(n_511), .B(n_556), .Y(n_555) );
INVx3_ASAP7_75t_L g562 ( .A(n_511), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_511), .B(n_531), .Y(n_574) );
INVxp67_ASAP7_75t_L g577 ( .A(n_511), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_511), .B(n_549), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_511), .B(n_521), .Y(n_643) );
AND2x2_ASAP7_75t_L g658 ( .A(n_511), .B(n_553), .Y(n_658) );
OR2x2_ASAP7_75t_L g687 ( .A(n_511), .B(n_521), .Y(n_687) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_519), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_520), .B(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_520), .B(n_556), .Y(n_695) );
OR2x2_ASAP7_75t_L g716 ( .A(n_520), .B(n_593), .Y(n_716) );
INVx1_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
OR2x2_ASAP7_75t_L g530 ( .A(n_521), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g553 ( .A(n_521), .B(n_549), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_521), .B(n_531), .Y(n_568) );
AND2x2_ASAP7_75t_L g638 ( .A(n_521), .B(n_562), .Y(n_638) );
AND2x2_ASAP7_75t_L g672 ( .A(n_521), .B(n_556), .Y(n_672) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_522), .B(n_556), .Y(n_575) );
AND2x2_ASAP7_75t_L g603 ( .A(n_522), .B(n_531), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_529), .B(n_611), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_530), .A2(n_618), .B1(n_654), .B2(n_671), .C(n_673), .Y(n_670) );
INVx5_ASAP7_75t_SL g549 ( .A(n_531), .Y(n_549) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B(n_535), .Y(n_532) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
OAI33xp33_ASAP7_75t_L g569 ( .A1(n_542), .A2(n_570), .A3(n_571), .B1(n_573), .B2(n_576), .B3(n_580), .Y(n_569) );
OR2x2_ASAP7_75t_L g585 ( .A(n_542), .B(n_586), .Y(n_585) );
AOI322xp5_ASAP7_75t_L g694 ( .A1(n_542), .A2(n_611), .A3(n_618), .B1(n_695), .B2(n_696), .C1(n_697), .C2(n_700), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_542), .B(n_570), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_SL g718 ( .A1(n_542), .A2(n_570), .B(n_719), .C(n_721), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g557 ( .A1(n_543), .A2(n_558), .B1(n_563), .B2(n_566), .C(n_569), .Y(n_557) );
INVx1_ASAP7_75t_L g650 ( .A(n_543), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_543), .B(n_699), .Y(n_698) );
OAI22xp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_547), .B1(n_550), .B2(n_552), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g627 ( .A(n_548), .B(n_562), .Y(n_627) );
AND2x2_ASAP7_75t_L g685 ( .A(n_548), .B(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g593 ( .A(n_549), .B(n_556), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_549), .B(n_562), .Y(n_621) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_551), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_551), .B(n_629), .Y(n_683) );
OAI321xp33_ASAP7_75t_L g702 ( .A1(n_551), .A2(n_624), .A3(n_703), .B1(n_704), .B2(n_705), .C(n_706), .Y(n_702) );
INVx1_ASAP7_75t_L g669 ( .A(n_552), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_553), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g608 ( .A(n_553), .B(n_556), .Y(n_608) );
AOI321xp33_ASAP7_75t_L g666 ( .A1(n_553), .A2(n_570), .A3(n_667), .B1(n_668), .B2(n_669), .C(n_670), .Y(n_666) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g583 ( .A(n_555), .B(n_568), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_556), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_556), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_556), .B(n_642), .Y(n_679) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_L g602 ( .A(n_560), .B(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g567 ( .A(n_561), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g675 ( .A(n_562), .Y(n_675) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_565), .B(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g598 ( .A(n_570), .Y(n_598) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_572), .B(n_607), .Y(n_656) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
OR2x2_ASAP7_75t_L g620 ( .A(n_575), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g665 ( .A(n_575), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_576), .A2(n_623), .B1(n_626), .B2(n_628), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g720 ( .A(n_579), .B(n_643), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_584), .B1(n_588), .B2(n_594), .C(n_597), .Y(n_581) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
BUFx2_ASAP7_75t_L g618 ( .A(n_587), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
INVx1_ASAP7_75t_SL g664 ( .A(n_590), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_592), .B(n_642), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_592), .A2(n_660), .B(n_662), .Y(n_659) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g705 ( .A(n_593), .B(n_687), .Y(n_705) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_SL g607 ( .A(n_596), .Y(n_607) );
AOI21xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B(n_601), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g651 ( .A(n_603), .B(n_652), .Y(n_651) );
INVxp67_ASAP7_75t_L g713 ( .A(n_603), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_608), .B(n_609), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_607), .B(n_625), .Y(n_661) );
INVxp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g682 ( .A(n_611), .Y(n_682) );
NAND5xp2_ASAP7_75t_L g612 ( .A(n_613), .B(n_630), .C(n_639), .D(n_659), .E(n_666), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .B(n_619), .C(n_622), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g654 ( .A(n_618), .Y(n_654) );
CKINVDCx16_ASAP7_75t_R g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_626), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g668 ( .A(n_628), .Y(n_668) );
OAI21xp5_ASAP7_75t_SL g630 ( .A1(n_631), .A2(n_634), .B(n_636), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_631), .A2(n_685), .B1(n_688), .B2(n_690), .C(n_691), .Y(n_684) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
AOI321xp33_ASAP7_75t_L g639 ( .A1(n_632), .A2(n_640), .A3(n_644), .B1(n_645), .B2(n_651), .C(n_653), .Y(n_639) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g710 ( .A(n_644), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_646), .B(n_650), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g662 ( .A(n_647), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
NOR2xp67_ASAP7_75t_SL g674 ( .A(n_648), .B(n_655), .Y(n_674) );
AOI321xp33_ASAP7_75t_SL g706 ( .A1(n_651), .A2(n_707), .A3(n_708), .B1(n_709), .B2(n_710), .C(n_711), .Y(n_706) );
O2A1O1Ixp33_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B(n_656), .C(n_657), .Y(n_653) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_664), .B(n_672), .Y(n_701) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND3xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .C(n_676), .Y(n_673) );
NOR3xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_702), .C(n_714), .Y(n_677) );
OAI211xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_680), .B(n_684), .C(n_694), .Y(n_678) );
INVxp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_682), .B(n_683), .Y(n_681) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_683), .A2(n_715), .B1(n_716), .B2(n_717), .C(n_718), .Y(n_714) );
INVx1_ASAP7_75t_L g703 ( .A(n_685), .Y(n_703) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g707 ( .A(n_705), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
CKINVDCx14_ASAP7_75t_R g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NOR2x2_ASAP7_75t_L g733 ( .A(n_725), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx3_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
NAND2xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_741), .Y(n_736) );
NOR2xp33_ASAP7_75t_SL g737 ( .A(n_738), .B(n_740), .Y(n_737) );
INVx1_ASAP7_75t_SL g762 ( .A(n_738), .Y(n_762) );
INVx1_ASAP7_75t_L g761 ( .A(n_740), .Y(n_761) );
OA21x2_ASAP7_75t_L g765 ( .A1(n_740), .A2(n_762), .B(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
NOR3xp33_ASAP7_75t_L g749 ( .A(n_742), .B(n_750), .C(n_755), .Y(n_749) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g746 ( .A(n_743), .Y(n_746) );
BUFx2_ASAP7_75t_L g766 ( .A(n_743), .Y(n_766) );
A2O1A1Ixp33_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_747), .B(n_758), .C(n_763), .Y(n_744) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g757 ( .A(n_751), .Y(n_757) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_759), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_762), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
endmodule