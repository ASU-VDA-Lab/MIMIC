module fake_jpeg_8979_n_226 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_30),
.A2(n_23),
.B1(n_17),
.B2(n_22),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

NOR4xp25_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_7),
.C(n_12),
.D(n_11),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_37),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_40),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_17),
.B1(n_22),
.B2(n_25),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_15),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_49),
.B1(n_15),
.B2(n_16),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_30),
.A2(n_23),
.B1(n_25),
.B2(n_27),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_14),
.B1(n_27),
.B2(n_24),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_33),
.C(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_39),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_23),
.B1(n_29),
.B2(n_24),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_31),
.A2(n_29),
.B1(n_14),
.B2(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_59),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_67),
.B1(n_74),
.B2(n_49),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_64),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_62),
.B(n_77),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_33),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_70),
.Y(n_91)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

OR2x2_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_26),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_16),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_39),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_69),
.A2(n_53),
.B(n_43),
.C(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_39),
.Y(n_70)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_19),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_94),
.C(n_97),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_67),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_81),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_59),
.B1(n_69),
.B2(n_61),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_72),
.B1(n_60),
.B2(n_34),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_85),
.A2(n_95),
.B(n_98),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_26),
.B(n_9),
.Y(n_114)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_100),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_70),
.B(n_52),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_41),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_54),
.C(n_34),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_64),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_45),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_9),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_62),
.B(n_10),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_58),
.B1(n_45),
.B2(n_65),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_102),
.A2(n_104),
.B1(n_118),
.B2(n_119),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_58),
.B1(n_65),
.B2(n_72),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_107),
.B1(n_111),
.B2(n_124),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_75),
.B1(n_36),
.B2(n_31),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_75),
.B1(n_38),
.B2(n_26),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_0),
.Y(n_113)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_118),
.B(n_119),
.Y(n_136)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_0),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_76),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_123),
.B1(n_98),
.B2(n_94),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_124),
.A2(n_80),
.B(n_97),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_140),
.B1(n_38),
.B2(n_56),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_85),
.B1(n_80),
.B2(n_81),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_146),
.B1(n_93),
.B2(n_76),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_114),
.B(n_79),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_134),
.B(n_139),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_143),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_142),
.B(n_125),
.Y(n_161)
);

AND2x4_ASAP7_75t_SL g139 ( 
.A(n_120),
.B(n_79),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_111),
.A2(n_94),
.B(n_83),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_88),
.B(n_83),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_147),
.B(n_11),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_96),
.C(n_38),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_105),
.C(n_116),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_104),
.A2(n_93),
.B1(n_86),
.B2(n_76),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_112),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_151),
.C(n_153),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_102),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_109),
.B(n_110),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_152),
.A2(n_156),
.B(n_161),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_107),
.C(n_96),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_96),
.C(n_115),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_162),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_155),
.B(n_158),
.Y(n_168)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_159),
.B(n_160),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_103),
.C(n_92),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_134),
.A2(n_92),
.B(n_1),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_5),
.Y(n_182)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_148),
.A2(n_131),
.B1(n_137),
.B2(n_147),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_166),
.A2(n_167),
.B1(n_132),
.B2(n_136),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_126),
.A2(n_138),
.B1(n_148),
.B2(n_142),
.Y(n_167)
);

AOI321xp33_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_144),
.A3(n_127),
.B1(n_136),
.B2(n_130),
.C(n_135),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_172),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_167),
.A2(n_143),
.B1(n_135),
.B2(n_130),
.Y(n_173)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

AO22x2_ASAP7_75t_L g174 ( 
.A1(n_161),
.A2(n_133),
.B1(n_129),
.B2(n_132),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_174),
.A2(n_175),
.B1(n_182),
.B2(n_162),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_164),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_157),
.Y(n_185)
);

BUFx24_ASAP7_75t_SL g178 ( 
.A(n_158),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_181),
.B(n_163),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_191),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_153),
.Y(n_188)
);

INVxp67_ASAP7_75t_SL g197 ( 
.A(n_188),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_170),
.B1(n_150),
.B2(n_171),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_175),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_192),
.A2(n_193),
.B(n_194),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_168),
.B(n_151),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_182),
.Y(n_196)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_172),
.B1(n_189),
.B2(n_186),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_198),
.B(n_201),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_169),
.C(n_171),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_154),
.C(n_150),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_191),
.A2(n_180),
.B1(n_176),
.B2(n_169),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_204),
.B(n_0),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_207),
.C(n_211),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_193),
.C(n_6),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_202),
.B(n_199),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_3),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_198),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_3),
.B(n_8),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_207),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_215),
.Y(n_219)
);

NOR2xp67_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_197),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_203),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_218),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_201),
.Y(n_220)
);

AOI321xp33_ASAP7_75t_L g222 ( 
.A1(n_220),
.A2(n_212),
.A3(n_206),
.B1(n_196),
.B2(n_13),
.C(n_8),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_219),
.C(n_8),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_223),
.A2(n_221),
.B(n_13),
.Y(n_224)
);

AOI221xp5_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_1),
.B1(n_2),
.B2(n_13),
.C(n_218),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_2),
.Y(n_226)
);


endmodule