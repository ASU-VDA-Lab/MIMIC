module fake_jpeg_14289_n_586 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_586);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_586;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_17),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_36),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g145 ( 
.A(n_61),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_62),
.Y(n_191)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_65),
.B(n_83),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_66),
.B(n_74),
.Y(n_127)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_69),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_19),
.B(n_17),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_70),
.B(n_85),
.Y(n_140)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_1),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_75),
.Y(n_154)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_79),
.Y(n_202)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_80),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_81),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_3),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_82),
.B(n_122),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_18),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_19),
.B(n_3),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_92),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_35),
.B(n_4),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_93),
.B(n_116),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_4),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_59),
.Y(n_166)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_97),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_18),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_104),
.Y(n_168)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx6_ASAP7_75t_SL g104 ( 
.A(n_20),
.Y(n_104)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_35),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_106),
.B(n_108),
.Y(n_171)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_37),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_37),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_110),
.B(n_113),
.Y(n_180)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_26),
.Y(n_111)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_27),
.B(n_4),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_23),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_114),
.B(n_115),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_21),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_27),
.B(n_40),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_41),
.Y(n_117)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_117),
.Y(n_177)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

INVx11_ASAP7_75t_SL g119 ( 
.A(n_58),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_119),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

BUFx24_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_121),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_29),
.B(n_4),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_42),
.Y(n_123)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_29),
.B(n_5),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_125),
.B(n_38),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_44),
.Y(n_126)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_126),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_132),
.B(n_139),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_62),
.A2(n_55),
.B1(n_42),
.B2(n_56),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_134),
.A2(n_197),
.B(n_186),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_66),
.A2(n_52),
.B(n_51),
.C(n_45),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g213 ( 
.A1(n_136),
.A2(n_51),
.B1(n_28),
.B2(n_45),
.Y(n_213)
);

AOI21xp33_ASAP7_75t_L g139 ( 
.A1(n_74),
.A2(n_40),
.B(n_48),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_141),
.B(n_170),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_82),
.A2(n_53),
.B1(n_56),
.B2(n_42),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_142),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_63),
.A2(n_75),
.B1(n_67),
.B2(n_91),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_159),
.A2(n_193),
.B1(n_8),
.B2(n_9),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_95),
.B(n_38),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_161),
.B(n_184),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_166),
.B(n_129),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_121),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_96),
.B(n_44),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_173),
.B(n_186),
.C(n_202),
.Y(n_272)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_71),
.Y(n_178)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_61),
.B(n_32),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_185),
.Y(n_215)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_79),
.Y(n_183)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_69),
.B(n_32),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_102),
.B(n_31),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_68),
.A2(n_53),
.B1(n_55),
.B2(n_60),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_76),
.Y(n_194)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_194),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_118),
.B(n_49),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_204),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_62),
.A2(n_50),
.B1(n_49),
.B2(n_44),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_101),
.B(n_48),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_104),
.C(n_105),
.Y(n_209)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_73),
.Y(n_201)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_201),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_94),
.B(n_49),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_97),
.B(n_31),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_126),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_209),
.B(n_216),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_153),
.B(n_60),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_210),
.B(n_213),
.Y(n_290)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_211),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_127),
.A2(n_99),
.B1(n_84),
.B2(n_89),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_212),
.A2(n_235),
.B1(n_255),
.B2(n_247),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_136),
.B(n_52),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_214),
.B(n_233),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_171),
.Y(n_216)
);

AOI32xp33_ASAP7_75t_L g217 ( 
.A1(n_140),
.A2(n_78),
.A3(n_49),
.B1(n_44),
.B2(n_30),
.Y(n_217)
);

AOI32xp33_ASAP7_75t_L g288 ( 
.A1(n_217),
.A2(n_175),
.A3(n_207),
.B1(n_133),
.B2(n_151),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_80),
.B1(n_88),
.B2(n_92),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_218),
.A2(n_245),
.B1(n_256),
.B2(n_260),
.Y(n_316)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_219),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_221),
.B(n_239),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_128),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_223),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_166),
.A2(n_50),
.B1(n_117),
.B2(n_98),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_224),
.A2(n_265),
.B(n_253),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_195),
.A2(n_28),
.B1(n_30),
.B2(n_124),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_225),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_189),
.A2(n_120),
.B1(n_112),
.B2(n_109),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_226),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_149),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_228),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_137),
.A2(n_50),
.B1(n_119),
.B2(n_81),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_229),
.Y(n_330)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_158),
.Y(n_231)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_231),
.Y(n_280)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_138),
.Y(n_232)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_232),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_148),
.B(n_6),
.Y(n_233)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_128),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_234),
.Y(n_321)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_8),
.Y(n_239)
);

INVx13_ASAP7_75t_L g240 ( 
.A(n_131),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_240),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_146),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_242),
.B(n_249),
.Y(n_308)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_165),
.Y(n_243)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

NAND2xp33_ASAP7_75t_SL g306 ( 
.A(n_244),
.B(n_277),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_173),
.A2(n_147),
.B1(n_154),
.B2(n_159),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_246),
.A2(n_262),
.B1(n_278),
.B2(n_245),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_152),
.B(n_10),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_255),
.Y(n_286)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_157),
.Y(n_248)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_168),
.Y(n_249)
);

BUFx4f_ASAP7_75t_L g252 ( 
.A(n_169),
.Y(n_252)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_252),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_149),
.Y(n_253)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_158),
.Y(n_254)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_156),
.B(n_11),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_169),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_256)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_176),
.Y(n_257)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_257),
.Y(n_319)
);

NAND2x1_ASAP7_75t_SL g258 ( 
.A(n_145),
.B(n_12),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_258),
.A2(n_214),
.B(n_241),
.Y(n_305)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_177),
.Y(n_259)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_203),
.A2(n_14),
.B1(n_15),
.B2(n_167),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_162),
.B(n_14),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_261),
.B(n_268),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_203),
.A2(n_15),
.B1(n_150),
.B2(n_151),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_130),
.A2(n_135),
.B1(n_191),
.B2(n_134),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_263),
.A2(n_264),
.B1(n_143),
.B2(n_192),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_191),
.A2(n_164),
.B1(n_143),
.B2(n_192),
.Y(n_264)
);

OR2x4_ASAP7_75t_L g265 ( 
.A(n_172),
.B(n_145),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g266 ( 
.A1(n_197),
.A2(n_176),
.B1(n_205),
.B2(n_155),
.Y(n_266)
);

OA22x2_ASAP7_75t_L g289 ( 
.A1(n_266),
.A2(n_175),
.B1(n_144),
.B2(n_150),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_181),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_267),
.B(n_274),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_180),
.B(n_160),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_198),
.B(n_204),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_275),
.Y(n_310)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_164),
.Y(n_270)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_270),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_271),
.A2(n_258),
.B(n_253),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_277),
.C(n_224),
.Y(n_297)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_174),
.Y(n_273)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_273),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_187),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_129),
.B(n_202),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_174),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_276),
.Y(n_323)
);

INVx3_ASAP7_75t_SL g278 ( 
.A(n_205),
.Y(n_278)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_278),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_144),
.Y(n_279)
);

BUFx5_ASAP7_75t_L g331 ( 
.A(n_279),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_281),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_240),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_283),
.B(n_295),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_288),
.A2(n_301),
.B1(n_315),
.B2(n_297),
.Y(n_339)
);

AO21x2_ASAP7_75t_SL g361 ( 
.A1(n_289),
.A2(n_294),
.B(n_332),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_244),
.A2(n_207),
.B1(n_133),
.B2(n_163),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_292),
.Y(n_345)
);

AO21x2_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_155),
.B(n_163),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_208),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_297),
.B(n_324),
.C(n_326),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_268),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_299),
.B(n_314),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_305),
.B(n_336),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_309),
.A2(n_325),
.B1(n_316),
.B2(n_312),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_233),
.B(n_261),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_212),
.A2(n_272),
.B1(n_246),
.B2(n_266),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_210),
.B(n_215),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_320),
.B(n_317),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_269),
.B(n_220),
.C(n_251),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_271),
.A2(n_213),
.B1(n_262),
.B2(n_266),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_230),
.B(n_237),
.C(n_222),
.Y(n_326)
);

OAI32xp33_ASAP7_75t_L g332 ( 
.A1(n_265),
.A2(n_266),
.A3(n_232),
.B1(n_248),
.B2(n_238),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_332),
.B(n_334),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_333),
.A2(n_330),
.B(n_300),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_227),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_312),
.A2(n_228),
.B1(n_243),
.B2(n_211),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_338),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_339),
.A2(n_342),
.B1(n_346),
.B2(n_347),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_308),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_340),
.B(n_357),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_236),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_341),
.B(n_355),
.C(n_376),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_315),
.A2(n_250),
.B1(n_234),
.B2(n_257),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_331),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_343),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_285),
.B(n_270),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_344),
.B(n_378),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_301),
.A2(n_279),
.B1(n_223),
.B2(n_276),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_310),
.A2(n_273),
.B1(n_259),
.B2(n_231),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_286),
.B(n_219),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_349),
.B(n_350),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_286),
.B(n_252),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_252),
.C(n_310),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_352),
.B(n_291),
.C(n_303),
.Y(n_416)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_293),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_353),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_314),
.B(n_298),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_354),
.B(n_366),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_298),
.B(n_305),
.C(n_333),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_356),
.A2(n_361),
.B1(n_289),
.B2(n_328),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_287),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_311),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_358),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_359),
.B(n_360),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_336),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_327),
.Y(n_362)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_362),
.Y(n_384)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_321),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_363),
.Y(n_411)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_327),
.Y(n_364)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_364),
.Y(n_387)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_321),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_365),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_285),
.A2(n_294),
.B1(n_290),
.B2(n_300),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_326),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_367),
.B(n_368),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_304),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_284),
.Y(n_370)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_370),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_313),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_371),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_372),
.A2(n_296),
.B(n_280),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_284),
.B(n_294),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_374),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_294),
.A2(n_289),
.B1(n_309),
.B2(n_330),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_307),
.B(n_282),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_294),
.B(n_307),
.Y(n_378)
);

INVx8_ASAP7_75t_L g379 ( 
.A(n_331),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_379),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_335),
.A2(n_289),
.B(n_304),
.Y(n_380)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_380),
.A2(n_329),
.B(n_293),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_381),
.A2(n_385),
.B1(n_404),
.B2(n_412),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_375),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_382),
.B(n_392),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_356),
.A2(n_361),
.B1(n_369),
.B2(n_380),
.Y(n_385)
);

XOR2x1_ASAP7_75t_SL g386 ( 
.A(n_372),
.B(n_323),
.Y(n_386)
);

OAI21xp33_ASAP7_75t_L g423 ( 
.A1(n_386),
.A2(n_348),
.B(n_378),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_355),
.B(n_282),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_388),
.B(n_391),
.C(n_416),
.Y(n_438)
);

MAJx2_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_302),
.C(n_322),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_373),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_394),
.A2(n_409),
.B(n_348),
.Y(n_433)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_347),
.Y(n_396)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_396),
.Y(n_419)
);

AO21x1_ASAP7_75t_L g397 ( 
.A1(n_348),
.A2(n_328),
.B(n_329),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_397),
.Y(n_426)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_368),
.Y(n_399)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_399),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_360),
.A2(n_322),
.B(n_302),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_402),
.A2(n_351),
.B(n_345),
.Y(n_446)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_376),
.Y(n_403)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_403),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_361),
.A2(n_296),
.B1(n_319),
.B2(n_280),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_361),
.A2(n_319),
.B1(n_318),
.B2(n_323),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_398),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_418),
.B(n_421),
.Y(n_464)
);

BUFx5_ASAP7_75t_L g420 ( 
.A(n_399),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_420),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_408),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_423),
.A2(n_433),
.B(n_390),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_414),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_429),
.Y(n_457)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_384),
.Y(n_427)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_427),
.Y(n_452)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_384),
.Y(n_428)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_428),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_402),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_410),
.A2(n_377),
.B1(n_354),
.B2(n_349),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_430),
.A2(n_434),
.B1(n_440),
.B2(n_447),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_397),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_432),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_410),
.A2(n_350),
.B1(n_337),
.B2(n_374),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_387),
.Y(n_435)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_435),
.Y(n_455)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_387),
.Y(n_436)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_436),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_413),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_445),
.Y(n_462)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_393),
.Y(n_439)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_439),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_400),
.A2(n_352),
.B1(n_337),
.B2(n_366),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_400),
.B(n_383),
.Y(n_441)
);

CKINVDCx14_ASAP7_75t_R g450 ( 
.A(n_441),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_389),
.B(n_341),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_442),
.B(n_411),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_385),
.A2(n_342),
.B1(n_346),
.B2(n_345),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_443),
.A2(n_396),
.B1(n_397),
.B2(n_406),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_392),
.B(n_383),
.Y(n_444)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_444),
.Y(n_468)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_393),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_446),
.A2(n_409),
.B(n_405),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_401),
.A2(n_344),
.B1(n_353),
.B2(n_363),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_401),
.A2(n_365),
.B1(n_318),
.B2(n_379),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_448),
.A2(n_407),
.B1(n_411),
.B2(n_415),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_451),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_438),
.B(n_388),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_453),
.B(n_461),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_456),
.A2(n_460),
.B1(n_465),
.B2(n_477),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_431),
.A2(n_406),
.B1(n_389),
.B2(n_394),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_438),
.B(n_405),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_404),
.Y(n_463)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_463),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_431),
.A2(n_386),
.B1(n_390),
.B2(n_403),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_469),
.A2(n_422),
.B1(n_419),
.B2(n_421),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_416),
.Y(n_470)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_470),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_441),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_471),
.B(n_472),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_434),
.Y(n_472)
);

XNOR2x1_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_391),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_453),
.C(n_461),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_475),
.A2(n_429),
.B(n_426),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_430),
.B(n_407),
.Y(n_476)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_476),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_443),
.A2(n_411),
.B1(n_415),
.B2(n_395),
.Y(n_477)
);

CKINVDCx14_ASAP7_75t_R g494 ( 
.A(n_478),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_475),
.A2(n_433),
.B(n_426),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_479),
.B(n_460),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_480),
.B(n_485),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_473),
.B(n_446),
.C(n_425),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_482),
.B(n_486),
.C(n_492),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_425),
.C(n_447),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_474),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_487),
.Y(n_511)
);

INVxp33_ASAP7_75t_L g488 ( 
.A(n_464),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_488),
.B(n_491),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_464),
.B(n_418),
.Y(n_489)
);

CKINVDCx14_ASAP7_75t_R g504 ( 
.A(n_489),
.Y(n_504)
);

OA21x2_ASAP7_75t_L g491 ( 
.A1(n_467),
.A2(n_432),
.B(n_457),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_451),
.B(n_424),
.C(n_422),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_493),
.A2(n_497),
.B1(n_477),
.B2(n_456),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_472),
.A2(n_419),
.B1(n_442),
.B2(n_448),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_457),
.B(n_445),
.C(n_439),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_498),
.B(n_455),
.C(n_459),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_462),
.B(n_420),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_499),
.B(n_500),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_417),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_467),
.B(n_436),
.Y(n_501)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_501),
.Y(n_507)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_452),
.Y(n_503)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_503),
.Y(n_513)
);

AOI21xp33_ASAP7_75t_L g509 ( 
.A1(n_489),
.A2(n_478),
.B(n_471),
.Y(n_509)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_509),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_492),
.B(n_466),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_510),
.B(n_518),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_512),
.A2(n_494),
.B(n_496),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_484),
.A2(n_466),
.B1(n_476),
.B2(n_468),
.Y(n_514)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_514),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_484),
.A2(n_481),
.B1(n_450),
.B2(n_463),
.Y(n_515)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_515),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_516),
.B(n_520),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_490),
.B(n_465),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_523),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_486),
.B(n_468),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_519),
.B(n_524),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_495),
.A2(n_469),
.B1(n_459),
.B2(n_458),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_495),
.A2(n_458),
.B1(n_455),
.B2(n_454),
.Y(n_522)
);

NOR2xp67_ASAP7_75t_SL g539 ( 
.A(n_522),
.B(n_503),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_497),
.A2(n_454),
.B1(n_452),
.B2(n_435),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_481),
.A2(n_427),
.B1(n_428),
.B2(n_395),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_490),
.C(n_480),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_526),
.B(n_530),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_508),
.B(n_483),
.C(n_502),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_519),
.B(n_483),
.C(n_502),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_531),
.B(n_522),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_521),
.A2(n_479),
.B(n_485),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_532),
.A2(n_534),
.B(n_535),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_533),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_521),
.A2(n_496),
.B(n_491),
.Y(n_534)
);

AO21x1_ASAP7_75t_L g535 ( 
.A1(n_507),
.A2(n_491),
.B(n_501),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_504),
.A2(n_501),
.B(n_498),
.Y(n_538)
);

AND2x2_ASAP7_75t_SL g544 ( 
.A(n_538),
.B(n_507),
.Y(n_544)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_539),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_505),
.C(n_518),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_541),
.B(n_550),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_536),
.A2(n_516),
.B1(n_523),
.B2(n_506),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_542),
.B(n_545),
.Y(n_560)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_544),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_530),
.B(n_531),
.C(n_525),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_528),
.B(n_511),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_547),
.B(n_551),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_525),
.B(n_505),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_548),
.B(n_534),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_527),
.B(n_517),
.C(n_514),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_538),
.B(n_511),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_540),
.B(n_482),
.C(n_520),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_553),
.B(n_527),
.C(n_529),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_554),
.A2(n_546),
.B(n_550),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_549),
.A2(n_532),
.B(n_533),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_557),
.B(n_559),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_545),
.B(n_529),
.C(n_537),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_561),
.B(n_564),
.Y(n_569)
);

OAI21xp33_ASAP7_75t_L g562 ( 
.A1(n_552),
.A2(n_537),
.B(n_535),
.Y(n_562)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_562),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_563),
.B(n_543),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_544),
.B(n_524),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_565),
.A2(n_543),
.B1(n_546),
.B2(n_544),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_567),
.B(n_563),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_556),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_568),
.B(n_570),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_560),
.A2(n_555),
.B(n_565),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g575 ( 
.A1(n_571),
.A2(n_558),
.B(n_562),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_559),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_573),
.B(n_548),
.Y(n_578)
);

A2O1A1O1Ixp25_ASAP7_75t_L g579 ( 
.A1(n_575),
.A2(n_577),
.B(n_578),
.C(n_568),
.D(n_573),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_576),
.Y(n_580)
);

NOR3xp33_ASAP7_75t_L g577 ( 
.A(n_572),
.B(n_566),
.C(n_569),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_SL g582 ( 
.A1(n_579),
.A2(n_581),
.B(n_513),
.Y(n_582)
);

OAI31xp33_ASAP7_75t_SL g581 ( 
.A1(n_574),
.A2(n_513),
.A3(n_493),
.B(n_417),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_582),
.B(n_583),
.C(n_291),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_580),
.B(n_343),
.C(n_303),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_584),
.B(n_358),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_585),
.B(n_311),
.Y(n_586)
);


endmodule