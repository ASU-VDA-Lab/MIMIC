module real_jpeg_25138_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_292;
wire n_215;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_105;
wire n_197;
wire n_299;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_297;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_209;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_273;
wire n_96;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_1),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_1),
.B(n_79),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_163),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_1),
.A2(n_28),
.B(n_48),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_1),
.B(n_120),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_1),
.A2(n_92),
.B1(n_248),
.B2(n_253),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_1),
.A2(n_61),
.B(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_2),
.A2(n_70),
.B1(n_71),
.B2(n_174),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_2),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_174),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_174),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_2),
.A2(n_28),
.B1(n_30),
.B2(n_174),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_4),
.A2(n_66),
.B1(n_70),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_4),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_115),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_115),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_4),
.A2(n_28),
.B1(n_30),
.B2(n_115),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g60 ( 
.A(n_6),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_7),
.A2(n_28),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_7),
.A2(n_36),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_7),
.A2(n_36),
.B1(n_61),
.B2(n_62),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_7),
.A2(n_36),
.B1(n_41),
.B2(n_42),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_8),
.A2(n_27),
.B1(n_61),
.B2(n_62),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_8),
.A2(n_27),
.B1(n_41),
.B2(n_42),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_8),
.A2(n_27),
.B1(n_70),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_9),
.A2(n_28),
.B1(n_30),
.B2(n_53),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_9),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_11),
.B(n_163),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_13),
.A2(n_44),
.B1(n_61),
.B2(n_62),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_13),
.A2(n_28),
.B1(n_30),
.B2(n_44),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_14),
.A2(n_68),
.B1(n_70),
.B2(n_73),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_14),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_14),
.A2(n_61),
.B1(n_62),
.B2(n_73),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_14),
.A2(n_28),
.B1(n_30),
.B2(n_73),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_73),
.Y(n_268)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_15),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_148),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_146),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_20),
.B(n_121),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_90),
.C(n_101),
.Y(n_20)
);

FAx1_ASAP7_75t_L g177 ( 
.A(n_21),
.B(n_90),
.CI(n_101),
.CON(n_177),
.SN(n_177)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_54),
.B2(n_89),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_22),
.B(n_55),
.C(n_80),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_24),
.B(n_39),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_25),
.A2(n_93),
.B(n_168),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_26),
.B(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_30),
.B1(n_48),
.B2(n_50),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_30),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_31),
.A2(n_106),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_31),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_33),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_33),
.B(n_163),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_34),
.A2(n_92),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_45),
.B1(n_51),
.B2(n_52),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_40),
.A2(n_51),
.B(n_111),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_42),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_41),
.A2(n_42),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_41),
.B(n_83),
.Y(n_273)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_42),
.A2(n_50),
.B(n_163),
.C(n_224),
.Y(n_223)
);

OAI32xp33_ASAP7_75t_L g272 ( 
.A1(n_42),
.A2(n_61),
.A3(n_82),
.B1(n_266),
.B2(n_273),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_45),
.A2(n_52),
.B(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_45),
.A2(n_51),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_45),
.A2(n_128),
.B(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_46),
.B(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_46),
.A2(n_98),
.B(n_129),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_46),
.A2(n_130),
.B1(n_222),
.B2(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_46),
.A2(n_130),
.B1(n_230),
.B2(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_51),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_51),
.B(n_163),
.Y(n_246)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_80),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_69),
.B(n_74),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_56),
.A2(n_57),
.B1(n_69),
.B2(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_56),
.A2(n_138),
.B(n_139),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_56),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_65),
.Y(n_56)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_59),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

OAI32xp33_ASAP7_75t_L g161 ( 
.A1(n_58),
.A2(n_62),
.A3(n_77),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_59),
.B(n_61),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_62),
.B1(n_82),
.B2(n_83),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_62),
.B(n_163),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_70),
.A2(n_162),
.B(n_163),
.Y(n_189)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_75),
.Y(n_138)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_79),
.B(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_79),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_79),
.A2(n_173),
.B1(n_175),
.B2(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B(n_85),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_81),
.B(n_118),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_81),
.A2(n_117),
.B1(n_206),
.B2(n_264),
.Y(n_263)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_84),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_86),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_86),
.A2(n_120),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_86),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_86),
.A2(n_120),
.B1(n_158),
.B2(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_86),
.A2(n_120),
.B1(n_191),
.B2(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_95),
.B1(n_96),
.B2(n_100),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_91),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_96),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_91),
.A2(n_100),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B(n_94),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_105),
.B(n_107),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_92),
.A2(n_238),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_92),
.A2(n_94),
.B(n_107),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_113),
.C(n_116),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_102),
.A2(n_103),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_110),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_104),
.B(n_110),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_113),
.B(n_116),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B(n_119),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_145),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_132),
.B1(n_143),
.B2(n_144),
.Y(n_122)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_127),
.B(n_131),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_124),
.B(n_127),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_142),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_178),
.B(n_301),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_177),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_150),
.B(n_177),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_151),
.B(n_182),
.Y(n_210)
);

FAx1_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_155),
.CI(n_156),
.CON(n_151),
.SN(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_172),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_172),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_165),
.B1(n_166),
.B2(n_201),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_161),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_177),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_211),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_193),
.B(n_210),
.Y(n_180)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_181),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.C(n_192),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_184),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_186),
.B(n_192),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.C(n_190),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_190),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_194),
.B(n_197),
.Y(n_300)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.C(n_202),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_198),
.B(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_200),
.A2(n_202),
.B1(n_203),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_200),
.Y(n_297)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.C(n_208),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_204),
.B(n_283),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_284),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_207),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_299),
.C(n_300),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_293),
.B(n_298),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_278),
.B(n_292),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_259),
.B(n_277),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_234),
.B(n_258),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_225),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_217),
.B(n_225),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_223),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_218),
.A2(n_219),
.B1(n_223),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_223),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_232),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_231),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_231),
.C(n_232),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_229),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_233),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_244),
.B(n_257),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_242),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_236),
.B(n_242),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_251),
.B(n_256),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_246),
.B(n_247),
.Y(n_256)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_260),
.B(n_261),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_271),
.B1(n_275),
.B2(n_276),
.Y(n_261)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_262)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_270),
.C(n_275),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_268),
.Y(n_289)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_271),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_274),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_280),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_285),
.B2(n_286),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_288),
.C(n_290),
.Y(n_294)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_288),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);


endmodule