module real_jpeg_6499_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_0),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_1),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_2),
.A2(n_27),
.B1(n_209),
.B2(n_212),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_3),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_3),
.A2(n_49),
.B1(n_83),
.B2(n_85),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_3),
.A2(n_49),
.B1(n_78),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_3),
.A2(n_49),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_4),
.Y(n_172)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_5),
.Y(n_108)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_6),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_6),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_6),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_7),
.A2(n_83),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_7),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_7),
.A2(n_89),
.B1(n_133),
.B2(n_137),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_7),
.A2(n_89),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_7),
.A2(n_89),
.B1(n_293),
.B2(n_295),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_8),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_14)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_11),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_12),
.A2(n_66),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_12),
.A2(n_66),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_12),
.A2(n_66),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_12),
.B(n_77),
.Y(n_239)
);

O2A1O1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_12),
.A2(n_256),
.B(n_257),
.C(n_263),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_12),
.B(n_284),
.C(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_12),
.B(n_148),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_12),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_12),
.B(n_165),
.Y(n_325)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_13),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_13),
.Y(n_161)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_13),
.Y(n_168)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_226),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_224),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_193),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_22),
.B(n_193),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_138),
.C(n_180),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_23),
.B(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_74),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_24),
.B(n_75),
.C(n_101),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_52),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_25),
.B(n_52),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_36),
.B(n_40),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_26),
.A2(n_182),
.B(n_183),
.Y(n_181)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_30),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_30),
.Y(n_295)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_35),
.Y(n_205)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_37),
.B(n_46),
.Y(n_183)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_39),
.Y(n_310)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_40),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_46),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_41),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_41),
.B(n_201),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_41),
.A2(n_201),
.B(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_41),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_51),
.Y(n_285)
);

AOI32xp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_57),
.A3(n_59),
.B1(n_62),
.B2(n_67),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AO22x1_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_77)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_63),
.A2(n_66),
.B(n_83),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_66),
.A2(n_258),
.B(n_260),
.Y(n_257)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_68),
.Y(n_263)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_71),
.Y(n_95)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_101),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_87),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_82),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_77),
.B(n_88),
.Y(n_152)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_82),
.B(n_92),
.Y(n_221)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_92),
.B(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_99),
.Y(n_93)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_121),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_116),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_109),
.B1(n_112),
.B2(n_114),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_114),
.Y(n_259)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_SL g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_117),
.A2(n_122),
.B(n_148),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_117),
.B(n_122),
.Y(n_336)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_121),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_132),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_130),
.Y(n_124)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_128),
.Y(n_256)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_132),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_138),
.B(n_180),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_149),
.C(n_153),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_139),
.A2(n_153),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_139),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_147),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_143),
.B(n_148),
.Y(n_237)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_147),
.B(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_149),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_152),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_153),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_173),
.B(n_174),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_175),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_155),
.B(n_187),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_155),
.B(n_272),
.Y(n_271)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_165),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

AO22x1_ASAP7_75t_SL g165 ( 
.A1(n_158),
.A2(n_166),
.B1(n_169),
.B2(n_171),
.Y(n_165)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_160),
.Y(n_284)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_164),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_164),
.Y(n_275)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_165),
.B(n_272),
.Y(n_287)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

BUFx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_172),
.Y(n_294)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_172),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_173),
.A2(n_208),
.B(n_215),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_173),
.B(n_174),
.Y(n_270)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_184),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_183),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_183),
.B(n_291),
.Y(n_324)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_185),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_186),
.B(n_271),
.Y(n_297)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_216),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_207),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_206),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_198),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_206),
.B(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_215),
.B(n_287),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_244),
.B(n_348),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_242),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_228),
.B(n_242),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_233),
.C(n_235),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.C(n_240),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_252),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_240),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_241),
.B(n_307),
.Y(n_322)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_276),
.B(n_347),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_247),
.B(n_250),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.C(n_267),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_251),
.B(n_343),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_254),
.A2(n_267),
.B1(n_268),
.B2(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_254),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_264),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_255),
.A2(n_264),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_255),
.Y(n_339)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_283),
.Y(n_282)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_264),
.Y(n_338)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_341),
.B(n_346),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_329),
.B(n_340),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_301),
.B(n_328),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_288),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_288),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_286),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_282),
.B1(n_286),
.B2(n_304),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_296),
.Y(n_288)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_289),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_308),
.Y(n_307)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_297),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_298),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_299),
.C(n_331),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_311),
.B(n_327),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_305),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_323),
.B(n_326),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_322),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_320),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_325),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_332),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_332),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_337),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_335),
.C(n_337),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_345),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_342),
.B(n_345),
.Y(n_346)
);


endmodule