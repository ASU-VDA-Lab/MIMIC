module fake_jpeg_2057_n_632 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_632);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_632;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_18),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_59),
.Y(n_153)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_60),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_10),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_64),
.B(n_71),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_65),
.Y(n_151)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_66),
.Y(n_181)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_67),
.Y(n_164)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_68),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_69),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_70),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_57),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_74),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_75),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_78),
.Y(n_192)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_20),
.B(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_80),
.B(n_81),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_20),
.B(n_10),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_84),
.Y(n_155)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_40),
.Y(n_85)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_86),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_27),
.B(n_8),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_87),
.B(n_95),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_91),
.Y(n_190)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_54),
.B(n_8),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_97),
.Y(n_188)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_98),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_45),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_99),
.B(n_100),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_32),
.B(n_41),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_101),
.Y(n_201)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_27),
.B(n_8),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_107),
.B(n_111),
.Y(n_197)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_109),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

BUFx12f_ASAP7_75t_SL g111 ( 
.A(n_22),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_22),
.Y(n_112)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_38),
.Y(n_113)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_115),
.Y(n_211)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_12),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_5),
.Y(n_152)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_22),
.Y(n_118)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_118),
.Y(n_224)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_26),
.Y(n_120)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_121),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_26),
.Y(n_123)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_123),
.Y(n_206)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_28),
.Y(n_124)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_26),
.Y(n_126)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_126),
.Y(n_213)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_26),
.Y(n_127)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_127),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_46),
.Y(n_128)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_128),
.Y(n_208)
);

BUFx8_ASAP7_75t_L g129 ( 
.A(n_39),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_129),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_71),
.B(n_57),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_132),
.B(n_162),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_95),
.A2(n_46),
.B1(n_28),
.B2(n_37),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_138),
.A2(n_63),
.B1(n_65),
.B2(n_2),
.Y(n_248)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_37),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_141),
.B(n_0),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_64),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_149),
.A2(n_42),
.B1(n_44),
.B2(n_47),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_152),
.B(n_177),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_80),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_112),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_174),
.B(n_218),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_81),
.A2(n_39),
.B1(n_37),
.B2(n_53),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_175),
.A2(n_94),
.B1(n_88),
.B2(n_86),
.Y(n_243)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_85),
.Y(n_176)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_87),
.B(n_41),
.Y(n_177)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_67),
.Y(n_179)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_183),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_110),
.B(n_37),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_SL g237 ( 
.A1(n_185),
.A2(n_46),
.B(n_1),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_122),
.B(n_35),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_186),
.B(n_202),
.Y(n_270)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_194),
.Y(n_239)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_114),
.Y(n_198)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_66),
.Y(n_199)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_199),
.Y(n_275)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_61),
.B(n_34),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_123),
.B(n_55),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_216),
.Y(n_240)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_118),
.Y(n_209)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_209),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_62),
.B(n_33),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_212),
.B(n_222),
.Y(n_276)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_120),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_110),
.B(n_55),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_119),
.Y(n_217)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_217),
.Y(n_304)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_128),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_74),
.B(n_51),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_219),
.B(n_223),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_90),
.B(n_51),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_101),
.B(n_49),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_42),
.B1(n_44),
.B2(n_47),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_225),
.A2(n_261),
.B1(n_188),
.B2(n_151),
.Y(n_340)
);

BUFx2_ASAP7_75t_SL g226 ( 
.A(n_139),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_226),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_227),
.B(n_221),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_181),
.Y(n_228)
);

NAND3xp33_ASAP7_75t_L g322 ( 
.A(n_228),
.B(n_232),
.C(n_235),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_133),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_230),
.Y(n_341)
);

AO22x1_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_129),
.B1(n_39),
.B2(n_37),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_231),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_181),
.Y(n_232)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_234),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_219),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_180),
.B(n_49),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_236),
.B(n_250),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_237),
.Y(n_320)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_173),
.Y(n_238)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_238),
.Y(n_325)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_142),
.Y(n_242)
);

INVx3_ASAP7_75t_SL g357 ( 
.A(n_242),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_243),
.A2(n_255),
.B1(n_280),
.B2(n_283),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_165),
.A2(n_75),
.B1(n_70),
.B2(n_69),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_246),
.A2(n_248),
.B1(n_259),
.B2(n_273),
.Y(n_352)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_142),
.Y(n_247)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_247),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_223),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_249),
.B(n_256),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_180),
.B(n_12),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_135),
.Y(n_251)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_251),
.Y(n_364)
);

INVx11_ASAP7_75t_L g253 ( 
.A(n_171),
.Y(n_253)
);

BUFx2_ASAP7_75t_SL g356 ( 
.A(n_253),
.Y(n_356)
);

INVx3_ASAP7_75t_SL g254 ( 
.A(n_192),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_254),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_165),
.A2(n_12),
.B1(n_17),
.B2(n_16),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_216),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_161),
.Y(n_257)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_257),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_175),
.A2(n_6),
.B1(n_16),
.B2(n_15),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_160),
.A2(n_6),
.B1(n_15),
.B2(n_14),
.Y(n_261)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_262),
.Y(n_334)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_172),
.Y(n_263)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_264),
.Y(n_342)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_178),
.Y(n_266)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_266),
.Y(n_310)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_131),
.Y(n_267)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_267),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_153),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_269),
.Y(n_360)
);

BUFx12f_ASAP7_75t_L g271 ( 
.A(n_224),
.Y(n_271)
);

INVx5_ASAP7_75t_L g358 ( 
.A(n_271),
.Y(n_358)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_134),
.Y(n_272)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_L g273 ( 
.A1(n_157),
.A2(n_184),
.B1(n_207),
.B2(n_208),
.Y(n_273)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_133),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_274),
.Y(n_316)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_164),
.Y(n_277)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_277),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_145),
.B(n_0),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_285),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_145),
.B(n_4),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_279),
.B(n_289),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_158),
.A2(n_4),
.B1(n_14),
.B2(n_13),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_213),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_281),
.Y(n_354)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_190),
.Y(n_282)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_282),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_158),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_163),
.B(n_6),
.C(n_18),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_284),
.B(n_168),
.C(n_206),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_166),
.B(n_0),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_224),
.Y(n_286)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_286),
.Y(n_351)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_167),
.Y(n_287)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_287),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_205),
.B(n_1),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_288),
.B(n_294),
.Y(n_350)
);

AOI21xp33_ASAP7_75t_L g289 ( 
.A1(n_185),
.A2(n_18),
.B(n_2),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_137),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_290),
.A2(n_295),
.B1(n_221),
.B2(n_189),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_192),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_291),
.B(n_303),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_136),
.Y(n_292)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_292),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_191),
.Y(n_293)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_140),
.B(n_3),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_146),
.A2(n_3),
.B1(n_150),
.B2(n_147),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_141),
.B(n_3),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_296),
.B(n_299),
.Y(n_355)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_164),
.Y(n_297)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

BUFx4f_ASAP7_75t_SL g298 ( 
.A(n_203),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_148),
.B(n_3),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_191),
.Y(n_300)
);

INVxp33_ASAP7_75t_L g362 ( 
.A(n_300),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_154),
.A2(n_195),
.B1(n_155),
.B2(n_193),
.Y(n_302)
);

OAI22x1_ASAP7_75t_L g363 ( 
.A1(n_302),
.A2(n_169),
.B1(n_220),
.B2(n_203),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_156),
.B(n_159),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_203),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_305),
.B(n_171),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_248),
.A2(n_211),
.B1(n_182),
.B2(n_215),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_313),
.A2(n_318),
.B1(n_273),
.B2(n_231),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_317),
.A2(n_326),
.B1(n_253),
.B2(n_274),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_270),
.A2(n_182),
.B1(n_136),
.B2(n_215),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_268),
.B(n_241),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_321),
.B(n_331),
.C(n_284),
.Y(n_386)
);

MAJx2_ASAP7_75t_L g331 ( 
.A(n_268),
.B(n_130),
.C(n_143),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_265),
.B(n_170),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_332),
.B(n_344),
.Y(n_368)
);

NAND2xp33_ASAP7_75t_SL g410 ( 
.A(n_337),
.B(n_239),
.Y(n_410)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_233),
.Y(n_338)
);

BUFx2_ASAP7_75t_SL g380 ( 
.A(n_338),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_340),
.B(n_346),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_260),
.B(n_204),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_276),
.B(n_210),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_345),
.B(n_347),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_240),
.B(n_196),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_245),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_240),
.B(n_287),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_348),
.B(n_229),
.Y(n_404)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_275),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_353),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_359),
.B(n_229),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_363),
.A2(n_254),
.B1(n_300),
.B2(n_282),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_366),
.A2(n_399),
.B1(n_362),
.B2(n_316),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_333),
.A2(n_243),
.B1(n_296),
.B2(n_285),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_367),
.A2(n_373),
.B1(n_408),
.B2(n_363),
.Y(n_423)
);

INVx8_ASAP7_75t_L g369 ( 
.A(n_341),
.Y(n_369)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_369),
.Y(n_411)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_329),
.Y(n_370)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_370),
.Y(n_446)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_314),
.Y(n_371)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_329),
.Y(n_372)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_372),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_307),
.B(n_264),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_374),
.Y(n_440)
);

INVx8_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_375),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_350),
.B(n_288),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_376),
.B(n_391),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_335),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_377),
.B(n_394),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_307),
.A2(n_264),
.B(n_243),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_378),
.A2(n_409),
.B(n_325),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_361),
.Y(n_379)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_379),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_331),
.B(n_303),
.Y(n_381)
);

NOR2x1_ASAP7_75t_L g417 ( 
.A(n_381),
.B(n_355),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_322),
.A2(n_278),
.B(n_283),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_382),
.A2(n_339),
.B(n_306),
.Y(n_429)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_327),
.Y(n_383)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

INVx8_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_384),
.Y(n_431)
);

MAJx2_ASAP7_75t_L g385 ( 
.A(n_321),
.B(n_294),
.C(n_299),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_389),
.C(n_401),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_386),
.B(n_406),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_324),
.A2(n_243),
.B1(n_234),
.B2(n_304),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_SL g447 ( 
.A1(n_387),
.A2(n_396),
.B1(n_325),
.B2(n_311),
.Y(n_447)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_327),
.Y(n_388)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_388),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_342),
.B(n_244),
.C(n_301),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_328),
.Y(n_390)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_390),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_350),
.B(n_257),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_392),
.Y(n_444)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_330),
.Y(n_393)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_393),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_323),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_352),
.A2(n_297),
.B1(n_277),
.B2(n_286),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_395),
.A2(n_400),
.B1(n_316),
.B2(n_314),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_358),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_362),
.Y(n_427)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_309),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_398),
.B(n_404),
.Y(n_416)
);

OAI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_317),
.A2(n_242),
.B1(n_247),
.B2(n_251),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_352),
.A2(n_272),
.B1(n_267),
.B2(n_252),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_359),
.B(n_263),
.C(n_266),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_356),
.A2(n_293),
.B1(n_262),
.B2(n_271),
.Y(n_405)
);

INVxp33_ASAP7_75t_L g433 ( 
.A(n_405),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_312),
.B(n_269),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_407),
.B(n_311),
.Y(n_443)
);

OAI22xp33_ASAP7_75t_L g408 ( 
.A1(n_313),
.A2(n_230),
.B1(n_292),
.B2(n_189),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_320),
.A2(n_298),
.B(n_238),
.Y(n_409)
);

INVxp33_ASAP7_75t_L g439 ( 
.A(n_410),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_414),
.A2(n_423),
.B1(n_426),
.B2(n_383),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_417),
.B(n_393),
.Y(n_475)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_422),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_378),
.A2(n_381),
.B1(n_395),
.B2(n_367),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_424),
.A2(n_435),
.B1(n_437),
.B2(n_374),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_381),
.A2(n_400),
.B1(n_373),
.B2(n_365),
.Y(n_426)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_427),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_428),
.A2(n_374),
.B(n_397),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_429),
.B(n_443),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_386),
.C(n_401),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_432),
.B(n_442),
.C(n_445),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_391),
.A2(n_306),
.B1(n_355),
.B2(n_318),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_368),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_436),
.B(n_438),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_377),
.A2(n_316),
.B1(n_351),
.B2(n_361),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_402),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_385),
.B(n_354),
.C(n_336),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_376),
.B(n_351),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_447),
.A2(n_357),
.B1(n_371),
.B2(n_343),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_423),
.A2(n_409),
.B1(n_396),
.B2(n_402),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_449),
.A2(n_451),
.B1(n_461),
.B2(n_462),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_450),
.A2(n_454),
.B(n_481),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_425),
.B(n_370),
.Y(n_452)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_452),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_428),
.A2(n_382),
.B(n_394),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_425),
.B(n_372),
.Y(n_456)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_456),
.Y(n_497)
);

MAJx2_ASAP7_75t_L g457 ( 
.A(n_421),
.B(n_389),
.C(n_407),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_457),
.B(n_475),
.Y(n_492)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_418),
.Y(n_458)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_458),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_404),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_459),
.B(n_469),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_413),
.B(n_388),
.Y(n_460)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_460),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_424),
.A2(n_408),
.B1(n_403),
.B2(n_380),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_427),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_463),
.B(n_470),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_390),
.Y(n_464)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_464),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_421),
.B(n_403),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_465),
.B(n_310),
.Y(n_513)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_411),
.Y(n_467)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_467),
.Y(n_511)
);

OAI22x1_ASAP7_75t_L g498 ( 
.A1(n_468),
.A2(n_480),
.B1(n_411),
.B2(n_271),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_417),
.B(n_364),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_418),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_426),
.A2(n_375),
.B1(n_369),
.B2(n_398),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_471),
.A2(n_476),
.B1(n_441),
.B2(n_444),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_417),
.B(n_364),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_472),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_416),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_474),
.B(n_477),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_435),
.A2(n_392),
.B1(n_379),
.B2(n_384),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_430),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_416),
.B(n_379),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_478),
.B(n_431),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_432),
.B(n_336),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_479),
.B(n_483),
.C(n_448),
.Y(n_496)
);

OAI21x1_ASAP7_75t_R g480 ( 
.A1(n_439),
.A2(n_308),
.B(n_358),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_440),
.A2(n_357),
.B(n_349),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_412),
.B(n_309),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_445),
.A2(n_343),
.B1(n_334),
.B2(n_144),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_484),
.A2(n_422),
.B1(n_437),
.B2(n_431),
.Y(n_486)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_485),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_486),
.A2(n_494),
.B1(n_495),
.B2(n_462),
.Y(n_528)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_488),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_451),
.A2(n_429),
.B1(n_430),
.B2(n_434),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_490),
.A2(n_463),
.B1(n_474),
.B2(n_449),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_482),
.B(n_412),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_491),
.B(n_504),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_453),
.A2(n_434),
.B1(n_443),
.B2(n_433),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_453),
.A2(n_442),
.B1(n_441),
.B2(n_444),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_496),
.B(n_505),
.C(n_517),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_498),
.B(n_468),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_450),
.A2(n_448),
.B(n_446),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_500),
.A2(n_493),
.B(n_515),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_479),
.B(n_446),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_512),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_334),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_483),
.B(n_415),
.C(n_419),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_482),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_514),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_466),
.B(n_415),
.Y(n_509)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_509),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_465),
.B(n_310),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_516),
.Y(n_529)
);

AOI21xp33_ASAP7_75t_L g514 ( 
.A1(n_454),
.A2(n_419),
.B(n_420),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_473),
.B(n_319),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_473),
.B(n_319),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_516),
.B(n_457),
.C(n_475),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_521),
.B(n_525),
.C(n_536),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_455),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_522),
.B(n_534),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_523),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_496),
.B(n_455),
.C(n_456),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_515),
.Y(n_526)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_526),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_528),
.A2(n_531),
.B1(n_537),
.B2(n_542),
.Y(n_562)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_507),
.Y(n_530)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_530),
.Y(n_555)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_507),
.Y(n_533)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_533),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_505),
.B(n_460),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_501),
.B(n_513),
.C(n_492),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_502),
.A2(n_471),
.B1(n_452),
.B2(n_478),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_510),
.A2(n_497),
.B1(n_489),
.B2(n_486),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_538),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_492),
.B(n_464),
.C(n_476),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_539),
.B(n_544),
.C(n_499),
.Y(n_554)
);

A2O1A1Ixp33_ASAP7_75t_SL g553 ( 
.A1(n_540),
.A2(n_485),
.B(n_498),
.C(n_494),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_510),
.B(n_484),
.Y(n_541)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_541),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_497),
.A2(n_477),
.B1(n_470),
.B2(n_458),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_489),
.A2(n_481),
.B1(n_467),
.B2(n_480),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_543),
.B(n_493),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_512),
.B(n_495),
.C(n_490),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_SL g545 ( 
.A(n_506),
.B(n_480),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_545),
.B(n_500),
.Y(n_549)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_546),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_549),
.B(n_554),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_532),
.B(n_487),
.Y(n_552)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_552),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_553),
.A2(n_540),
.B1(n_543),
.B2(n_527),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_519),
.B(n_506),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_556),
.B(n_557),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_519),
.B(n_503),
.C(n_511),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_536),
.B(n_503),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_558),
.B(n_539),
.C(n_544),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_534),
.B(n_511),
.Y(n_559)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_559),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_525),
.B(n_298),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_560),
.B(n_561),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_521),
.B(n_529),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_529),
.B(n_420),
.C(n_315),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_563),
.B(n_518),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_557),
.B(n_524),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_567),
.B(n_570),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_554),
.B(n_520),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_548),
.A2(n_531),
.B1(n_537),
.B2(n_535),
.Y(n_572)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_572),
.Y(n_593)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_555),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_574),
.B(n_575),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_550),
.A2(n_527),
.B1(n_541),
.B2(n_523),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_576),
.A2(n_553),
.B1(n_545),
.B2(n_565),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_562),
.B(n_538),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_577),
.B(n_582),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g595 ( 
.A(n_579),
.B(n_580),
.Y(n_595)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_564),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_558),
.B(n_518),
.C(n_522),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_583),
.B(n_584),
.C(n_551),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_563),
.B(n_551),
.C(n_565),
.Y(n_584)
);

NOR2xp67_ASAP7_75t_R g585 ( 
.A(n_568),
.B(n_566),
.Y(n_585)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_585),
.Y(n_601)
);

INVx6_ASAP7_75t_L g586 ( 
.A(n_571),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_586),
.B(n_581),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g587 ( 
.A1(n_568),
.A2(n_547),
.B(n_553),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_587),
.A2(n_588),
.B(n_591),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_575),
.A2(n_549),
.B(n_553),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_589),
.A2(n_577),
.B1(n_580),
.B2(n_583),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_SL g591 ( 
.A1(n_576),
.A2(n_577),
.B(n_569),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_592),
.B(n_597),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g597 ( 
.A(n_584),
.B(n_542),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_578),
.B(n_349),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_598),
.B(n_239),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_578),
.B(n_315),
.C(n_360),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_599),
.A2(n_258),
.B(n_592),
.Y(n_610)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_600),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_603),
.B(n_604),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_SL g604 ( 
.A1(n_593),
.A2(n_574),
.B1(n_582),
.B2(n_573),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_596),
.A2(n_360),
.B1(n_151),
.B2(n_144),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_605),
.B(n_606),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_590),
.B(n_258),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_608),
.B(n_609),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_595),
.B(n_252),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_610),
.A2(n_598),
.B(n_595),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_612),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_SL g614 ( 
.A1(n_602),
.A2(n_594),
.B(n_591),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g620 ( 
.A1(n_614),
.A2(n_617),
.B(n_588),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_600),
.A2(n_587),
.B(n_586),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_609),
.B(n_596),
.C(n_594),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_618),
.B(n_604),
.Y(n_621)
);

AO21x1_ASAP7_75t_L g619 ( 
.A1(n_613),
.A2(n_601),
.B(n_607),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_619),
.B(n_621),
.Y(n_626)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_620),
.Y(n_624)
);

NAND3xp33_ASAP7_75t_L g622 ( 
.A(n_611),
.B(n_585),
.C(n_599),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_622),
.B(n_618),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_625),
.B(n_623),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_627),
.A2(n_628),
.B(n_624),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_626),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_629),
.A2(n_615),
.B(n_616),
.Y(n_630)
);

INVxp67_ASAP7_75t_SL g631 ( 
.A(n_630),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_631),
.A2(n_589),
.B(n_608),
.Y(n_632)
);


endmodule