module fake_jpeg_10356_n_141 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_33),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_30),
.Y(n_43)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_29),
.A2(n_19),
.B1(n_22),
.B2(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_1),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_15),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_41),
.B1(n_19),
.B2(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_38),
.Y(n_48)
);

INVx5_ASAP7_75t_SL g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_39),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_19),
.B1(n_22),
.B2(n_20),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_51),
.B1(n_54),
.B2(n_61),
.Y(n_74)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_47),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_50),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_29),
.B1(n_17),
.B2(n_21),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_29),
.B1(n_16),
.B2(n_21),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_27),
.B1(n_12),
.B2(n_26),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_66),
.B1(n_43),
.B2(n_14),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_28),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_34),
.A2(n_18),
.B1(n_17),
.B2(n_15),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_13),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_14),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_26),
.C(n_23),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_38),
.B1(n_35),
.B2(n_45),
.Y(n_76)
);

OAI22x1_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_41),
.B1(n_26),
.B2(n_12),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_72),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_23),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_77),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_18),
.B1(n_38),
.B2(n_12),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_56),
.A2(n_14),
.B1(n_23),
.B2(n_5),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_48),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_89),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_61),
.B1(n_49),
.B2(n_67),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_98),
.B1(n_99),
.B2(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_59),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_55),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_52),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_74),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_58),
.B(n_57),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_84),
.B(n_73),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_57),
.B1(n_47),
.B2(n_23),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_39),
.B1(n_63),
.B2(n_5),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_2),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_69),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_103),
.A2(n_104),
.B1(n_96),
.B2(n_98),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_88),
.C(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_108),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_110),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_102),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_93),
.B1(n_103),
.B2(n_85),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_118),
.B(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_120),
.A2(n_121),
.B(n_119),
.Y(n_128)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_108),
.C(n_104),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_103),
.C(n_99),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_114),
.C(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_86),
.B1(n_79),
.B2(n_77),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_125),
.B(n_114),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_121),
.C(n_86),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_123),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_128),
.A2(n_130),
.B(n_86),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_119),
.B(n_86),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_132),
.B(n_133),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_85),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_2),
.B(n_4),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_8),
.Y(n_138)
);

AOI21x1_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_8),
.B(n_4),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.C(n_2),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_6),
.C(n_136),
.Y(n_141)
);


endmodule