module fake_jpeg_6716_n_158 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_158);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_22),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_33),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_34),
.B(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_6),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_36),
.B(n_38),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_39),
.B(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_14),
.Y(n_60)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_31),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_26),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_66),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_52),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_23),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_60),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_18),
.B1(n_20),
.B2(n_27),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_56),
.B(n_26),
.C(n_30),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_18),
.B1(n_20),
.B2(n_27),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_20),
.B1(n_18),
.B2(n_28),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_74),
.B(n_31),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_69),
.B(n_71),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_18),
.B1(n_21),
.B2(n_23),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_73),
.Y(n_88)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_28),
.B1(n_16),
.B2(n_14),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_16),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_16),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_81),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_71),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_93),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_26),
.B(n_17),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_68),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_70),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_62),
.B1(n_66),
.B2(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_0),
.Y(n_93)
);

AND2x6_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_17),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_SL g111 ( 
.A(n_94),
.B(n_98),
.C(n_54),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_17),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_1),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_2),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_17),
.C(n_31),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_78),
.C(n_63),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_31),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_53),
.B1(n_61),
.B2(n_65),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_107),
.B1(n_105),
.B2(n_122),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_51),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_112),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_113),
.B1(n_87),
.B2(n_97),
.Y(n_126)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

OAI32xp33_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_76),
.A3(n_58),
.B1(n_55),
.B2(n_49),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_117),
.B(n_118),
.Y(n_124)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_84),
.B(n_3),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_122),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_5),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_5),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_107),
.A2(n_87),
.B1(n_83),
.B2(n_90),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_120),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_83),
.B1(n_97),
.B2(n_101),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_128),
.B(n_129),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_82),
.B1(n_89),
.B2(n_93),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_102),
.C(n_92),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_137),
.A2(n_133),
.B1(n_132),
.B2(n_136),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_123),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_143),
.Y(n_148)
);

OA21x2_ASAP7_75t_SL g142 ( 
.A1(n_127),
.A2(n_111),
.B(n_116),
.Y(n_142)
);

XOR2x2_ASAP7_75t_L g145 ( 
.A(n_142),
.B(n_135),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_131),
.B1(n_125),
.B2(n_134),
.Y(n_144)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_130),
.C(n_100),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_146),
.A2(n_141),
.B(n_133),
.Y(n_149)
);

OR2x2_ASAP7_75t_SL g152 ( 
.A(n_150),
.B(n_148),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_146),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_147),
.C(n_144),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_150),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_154),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_9),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g157 ( 
.A(n_156),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_157),
.Y(n_158)
);


endmodule