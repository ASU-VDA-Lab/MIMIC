module real_jpeg_30089_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_0),
.Y(n_80)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_3),
.A2(n_24),
.B1(n_26),
.B2(n_34),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_3),
.A2(n_4),
.B1(n_34),
.B2(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_3),
.A2(n_34),
.B1(n_42),
.B2(n_43),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_SL g127 ( 
.A1(n_3),
.A2(n_28),
.B(n_72),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_3),
.B(n_70),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_SL g159 ( 
.A1(n_3),
.A2(n_10),
.B(n_24),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g179 ( 
.A1(n_3),
.A2(n_39),
.B(n_43),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_3),
.B(n_23),
.Y(n_182)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_4),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_4),
.A2(n_8),
.B1(n_31),
.B2(n_68),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_4),
.A2(n_34),
.B(n_71),
.C(n_127),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_5),
.A2(n_24),
.B1(n_26),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.Y(n_79)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_6),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_7),
.A2(n_24),
.B1(n_26),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_48),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_8),
.A2(n_24),
.B1(n_26),
.B2(n_31),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_8),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_129)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_10),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_10),
.Y(n_158)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_11),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_117),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_116),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_90),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_16),
.B(n_90),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_76),
.B2(n_89),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_50),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_36),
.B(n_49),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_36),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_20),
.A2(n_83),
.B1(n_94),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_20),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_20),
.B(n_148),
.C(n_149),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_20),
.A2(n_123),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_22),
.B(n_33),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_22),
.B(n_23),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_27),
.Y(n_22)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_26),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_24),
.A2(n_34),
.B(n_40),
.C(n_179),
.Y(n_178)
);

INVx5_ASAP7_75t_SL g29 ( 
.A(n_28),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_28),
.A2(n_29),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_28),
.A2(n_34),
.B(n_158),
.C(n_159),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_30),
.A2(n_35),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_32),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_34),
.B(n_80),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_34),
.B(n_41),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_45),
.B2(n_47),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_37),
.A2(n_41),
.B1(n_62),
.B2(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_37),
.B(n_41),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_45),
.B(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_42),
.B(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_57),
.Y(n_56)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_63),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_59),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_64),
.B1(n_65),
.B2(n_75),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_52),
.A2(n_59),
.B1(n_75),
.B2(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_56),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_55),
.B(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_56),
.A2(n_80),
.B1(n_104),
.B2(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_57),
.A2(n_101),
.B(n_129),
.Y(n_148)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_59),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_61),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_70),
.B1(n_73),
.B2(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_73),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_83),
.C(n_86),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_78),
.A2(n_81),
.B1(n_173),
.B2(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_78),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_81),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_81),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_81),
.A2(n_173),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_81),
.B(n_128),
.C(n_183),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_81),
.B(n_164),
.C(n_172),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_86),
.B1(n_87),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_83),
.B(n_123),
.C(n_124),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_86),
.A2(n_87),
.B1(n_133),
.B2(n_134),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_86),
.B(n_106),
.C(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_86),
.A2(n_87),
.B1(n_105),
.B2(n_106),
.Y(n_201)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_113),
.C(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.C(n_97),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_95),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_97),
.B(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_109),
.C(n_112),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_98),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_105),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_99),
.A2(n_105),
.B1(n_106),
.B2(n_139),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_99),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_105),
.A2(n_106),
.B1(n_178),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_106),
.B(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_113),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_223),
.B(n_228),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_151),
.B(n_211),
.C(n_222),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_140),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_120),
.B(n_140),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_130),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_121),
.B(n_131),
.C(n_138),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_128),
.A2(n_146),
.B1(n_181),
.B2(n_184),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_128),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_128),
.B(n_194),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_137),
.B2(n_138),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_147),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_141),
.B(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_142),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_147),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_148),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_210),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_204),
.B(n_209),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_174),
.B(n_203),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_163),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_163),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_157),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_162),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_169),
.B2(n_170),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_166),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_167),
.B(n_187),
.Y(n_196)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_171),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_198),
.B(n_202),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_185),
.B(n_197),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_180),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_178),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_181),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_182),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_189),
.B(n_196),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_193),
.B(n_195),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_206),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_213),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_220),
.B2(n_221),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_218),
.C(n_221),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_220),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_224),
.B(n_225),
.Y(n_228)
);


endmodule