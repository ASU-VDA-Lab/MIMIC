module fake_jpeg_8487_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_8),
.B(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_41),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_0),
.B(n_1),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_22),
.B1(n_20),
.B2(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_31),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_23),
.B1(n_19),
.B2(n_18),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_60),
.B1(n_29),
.B2(n_38),
.Y(n_81)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_18),
.B1(n_23),
.B2(n_19),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_63),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_23),
.B1(n_19),
.B2(n_18),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_80),
.B1(n_22),
.B2(n_20),
.Y(n_113)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_72),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_62),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_71),
.A2(n_89),
.B(n_30),
.Y(n_115)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_74),
.B(n_27),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_42),
.CI(n_53),
.CON(n_104),
.SN(n_104)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_29),
.B1(n_21),
.B2(n_16),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_77),
.A2(n_81),
.B1(n_86),
.B2(n_30),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_83),
.Y(n_93)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_37),
.B1(n_21),
.B2(n_30),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_51),
.B1(n_43),
.B2(n_44),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_44),
.A2(n_21),
.B1(n_16),
.B2(n_20),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_16),
.B(n_37),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_71),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_101),
.B1(n_105),
.B2(n_110),
.Y(n_131)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_92),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_71),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_95),
.B(n_99),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_96),
.A2(n_83),
.B1(n_88),
.B2(n_90),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_50),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_66),
.B(n_48),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_114),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_15),
.C(n_14),
.Y(n_137)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_48),
.B(n_30),
.C(n_21),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_107),
.A2(n_36),
.B(n_87),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_68),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_113),
.B(n_115),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_63),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_30),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_22),
.C(n_28),
.Y(n_134)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_57),
.B1(n_56),
.B2(n_69),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_119),
.A2(n_92),
.B1(n_106),
.B2(n_116),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_43),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_134),
.Y(n_166)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_143),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_82),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_133),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_78),
.B(n_84),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_137),
.B(n_139),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_34),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_91),
.B1(n_96),
.B2(n_104),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_146),
.B1(n_103),
.B2(n_28),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_136),
.A2(n_147),
.B1(n_110),
.B2(n_101),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_36),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_140),
.Y(n_155)
);

NOR2x1p5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_36),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_25),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_108),
.B(n_109),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_142),
.A2(n_32),
.B(n_10),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_93),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_25),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_145),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_25),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_105),
.A2(n_64),
.B1(n_88),
.B2(n_28),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_149),
.A2(n_159),
.B1(n_167),
.B2(n_124),
.Y(n_201)
);

HAxp5_ASAP7_75t_SL g150 ( 
.A(n_129),
.B(n_27),
.CON(n_150),
.SN(n_150)
);

NAND2xp33_ASAP7_75t_SL g203 ( 
.A(n_150),
.B(n_26),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_123),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_153),
.Y(n_186)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_152),
.B(n_154),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_106),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_146),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_160),
.Y(n_195)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_168),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_162),
.A2(n_172),
.B(n_173),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_32),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_136),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_127),
.A2(n_98),
.B1(n_100),
.B2(n_33),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_122),
.A2(n_17),
.B1(n_32),
.B2(n_33),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_177),
.B(n_180),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_103),
.B1(n_98),
.B2(n_33),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_145),
.B1(n_124),
.B2(n_132),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_25),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_131),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_120),
.B(n_98),
.Y(n_174)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_140),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_175),
.A2(n_176),
.B(n_178),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_130),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g178 ( 
.A1(n_120),
.A2(n_137),
.B(n_128),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_125),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_179),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_142),
.A2(n_25),
.B(n_26),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_158),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_181),
.B(n_194),
.Y(n_219)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_185),
.Y(n_210)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_175),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_126),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_207),
.C(n_208),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_166),
.B(n_138),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_190),
.B(n_206),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_198),
.B1(n_167),
.B2(n_179),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_148),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_143),
.B(n_139),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_196),
.A2(n_200),
.B(n_170),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_139),
.B1(n_125),
.B2(n_121),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_159),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_199),
.B(n_205),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_124),
.B(n_141),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_169),
.B1(n_160),
.B2(n_173),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_203),
.A2(n_161),
.B1(n_152),
.B2(n_162),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_148),
.Y(n_205)
);

XOR2x1_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_134),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_121),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_25),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_186),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_214),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_155),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_213),
.C(n_233),
.Y(n_239)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_215),
.A2(n_226),
.B1(n_228),
.B2(n_17),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_196),
.B1(n_195),
.B2(n_156),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_184),
.A2(n_163),
.B(n_164),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_218),
.A2(n_232),
.B(n_184),
.Y(n_237)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_151),
.Y(n_221)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_225),
.Y(n_247)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_197),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_154),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_227),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_209),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_189),
.B(n_180),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_230),
.B(n_207),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_182),
.B(n_164),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_0),
.B(n_1),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_200),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_177),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_33),
.B1(n_24),
.B2(n_17),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_188),
.B1(n_202),
.B2(n_185),
.Y(n_235)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_225),
.A2(n_182),
.B1(n_191),
.B2(n_206),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_236),
.A2(n_242),
.B1(n_243),
.B2(n_250),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_237),
.A2(n_26),
.B(n_15),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_238),
.B(n_244),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_209),
.B1(n_193),
.B2(n_202),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_230),
.B1(n_217),
.B2(n_220),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_208),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_238),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_217),
.B(n_193),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_246),
.B(n_244),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_194),
.C(n_24),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_210),
.C(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_219),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_213),
.B1(n_210),
.B2(n_221),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_255),
.A2(n_269),
.B1(n_236),
.B2(n_242),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_240),
.B(n_229),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_256),
.B(n_257),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_212),
.C(n_227),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_261),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_231),
.C(n_218),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_262),
.B(n_246),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_247),
.Y(n_265)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_265),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_267),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_233),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_269)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_270),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_274),
.B(n_26),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_255),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_279),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_278),
.B1(n_282),
.B2(n_284),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_253),
.B1(n_254),
.B2(n_248),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_245),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_249),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_13),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_263),
.A2(n_24),
.B1(n_14),
.B2(n_13),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_259),
.B(n_267),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_266),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_264),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_285),
.B(n_26),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_268),
.B(n_262),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_280),
.Y(n_297)
);

XNOR2x1_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_258),
.Y(n_288)
);

MAJx2_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_292),
.C(n_296),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_273),
.A2(n_269),
.B(n_258),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_290),
.A2(n_293),
.B(n_295),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_291),
.B(n_9),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_271),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_10),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_292),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_278),
.A2(n_277),
.B(n_281),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_297),
.B(n_300),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_284),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_301),
.B(n_302),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_305),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_288),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_5),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_307),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_286),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_299),
.B(n_293),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_310),
.A2(n_309),
.B(n_308),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_314),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_299),
.B(n_296),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_315),
.A2(n_313),
.B(n_6),
.Y(n_316)
);

OA21x2_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_5),
.B(n_6),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_7),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_7),
.B(n_8),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_319),
.Y(n_320)
);


endmodule