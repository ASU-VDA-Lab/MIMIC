module fake_netlist_5_2469_n_1917 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1917);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1917;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_196;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_783;
wire n_555;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1835;
wire n_1726;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g183 ( 
.A(n_2),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_130),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_179),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_63),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_62),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_95),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_126),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_166),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_96),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_77),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_26),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_6),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_101),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_128),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_134),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_48),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_72),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_38),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_36),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_45),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_20),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_135),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_154),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_3),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_11),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_97),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_129),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_1),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_20),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_113),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_54),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_54),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_149),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_169),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_40),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_70),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_100),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_115),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_50),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_75),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_143),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_165),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_112),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_107),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_147),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_61),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_79),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_85),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_42),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_38),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_46),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_93),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_87),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_42),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_63),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_119),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_174),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_14),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_0),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_74),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_32),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_81),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_167),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_8),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_178),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_88),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_53),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_144),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_89),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_16),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_90),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_35),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_67),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_51),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_73),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_155),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_48),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_164),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_5),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_86),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_111),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_109),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_5),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_1),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_104),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_0),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_14),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_56),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_121),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_133),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_53),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_127),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_25),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_36),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_30),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_76),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_50),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_153),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_59),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_2),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_162),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_64),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_158),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_8),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_40),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_78),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_83),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_181),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_10),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_175),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_31),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_35),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_142),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_15),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_16),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_177),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_105),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_3),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_170),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_32),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_18),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_125),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_159),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_71),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_140),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_25),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_47),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_91),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_43),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_114),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_139),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_27),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_45),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_66),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_156),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_120),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_116),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_34),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_168),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_150),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_92),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_173),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_56),
.Y(n_332)
);

INVx4_ASAP7_75t_R g333 ( 
.A(n_94),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_37),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_148),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_62),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_65),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_27),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_46),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_17),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_9),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_24),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_99),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_52),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_6),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_41),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_69),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_52),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_43),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_84),
.Y(n_350)
);

BUFx5_ASAP7_75t_L g351 ( 
.A(n_102),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_47),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_39),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_34),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_132),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_61),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_106),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_10),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_26),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_131),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_33),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_17),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_9),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_12),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_223),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_184),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_190),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_212),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_351),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_212),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_191),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_212),
.Y(n_372)
);

INVxp33_ASAP7_75t_L g373 ( 
.A(n_340),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_192),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_270),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_212),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_193),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_245),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_198),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_316),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_351),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_218),
.B(n_4),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_316),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_218),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g385 ( 
.A(n_336),
.B(n_4),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_306),
.B(n_7),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_336),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_199),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_340),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_320),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_201),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_205),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_277),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_277),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_253),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_295),
.Y(n_396)
);

INVxp33_ASAP7_75t_SL g397 ( 
.A(n_200),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_277),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_183),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_306),
.B(n_7),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_319),
.B(n_11),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_185),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_209),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_295),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_185),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_183),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_210),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_214),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_255),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_351),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_215),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_197),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_186),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_255),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_253),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_219),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_248),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_351),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_319),
.B(n_188),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_L g420 ( 
.A(n_186),
.B(n_12),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_197),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_194),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_222),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_225),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_227),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_226),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_194),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_195),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_195),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_206),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_206),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_229),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_232),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_228),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_234),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_228),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_259),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_241),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_242),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_308),
.Y(n_440)
);

NOR2xp67_ASAP7_75t_L g441 ( 
.A(n_259),
.B(n_13),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_263),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_263),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_246),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_283),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_249),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_268),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_251),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_252),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_254),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_268),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_273),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_188),
.B(n_13),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_262),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_264),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_351),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_369),
.Y(n_457)
);

BUFx8_ASAP7_75t_L g458 ( 
.A(n_417),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_369),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_399),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_396),
.B(n_267),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_L g462 ( 
.A(n_401),
.B(n_260),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_399),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_406),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_406),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_396),
.B(n_271),
.Y(n_466)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_369),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_413),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_413),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_381),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_422),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_381),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_381),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_410),
.Y(n_475)
);

OAI21x1_ASAP7_75t_L g476 ( 
.A1(n_410),
.A2(n_233),
.B(n_196),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_422),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_396),
.B(n_274),
.Y(n_478)
);

AND2x6_ASAP7_75t_L g479 ( 
.A(n_404),
.B(n_260),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_410),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_418),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_427),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_427),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_418),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_428),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_428),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_418),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_429),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_429),
.Y(n_489)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_404),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_431),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_456),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_431),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_404),
.B(n_278),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_456),
.Y(n_495)
);

BUFx8_ASAP7_75t_L g496 ( 
.A(n_417),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_456),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_434),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_419),
.B(n_189),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_L g500 ( 
.A(n_401),
.B(n_260),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_434),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_368),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_436),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_368),
.Y(n_504)
);

BUFx8_ASAP7_75t_L g505 ( 
.A(n_409),
.Y(n_505)
);

INVx5_ASAP7_75t_L g506 ( 
.A(n_404),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_393),
.B(n_295),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_436),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_442),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_370),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_382),
.A2(n_363),
.B1(n_235),
.B2(n_341),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_386),
.B(n_207),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_442),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_393),
.B(n_308),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_443),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_370),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_443),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_447),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_372),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_394),
.B(n_398),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_447),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_372),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_394),
.B(n_248),
.Y(n_523)
);

AND3x2_ASAP7_75t_L g524 ( 
.A(n_400),
.B(n_233),
.C(n_196),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_451),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_425),
.B(n_207),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_451),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_452),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_398),
.B(n_189),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_452),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_414),
.B(n_440),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_376),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_395),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_376),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_380),
.Y(n_535)
);

INVxp33_ASAP7_75t_SL g536 ( 
.A(n_511),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_520),
.B(n_409),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_520),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_461),
.B(n_366),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_520),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_460),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_512),
.B(n_237),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_512),
.B(n_237),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_505),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_457),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_460),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_490),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_463),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_526),
.A2(n_384),
.B1(n_454),
.B2(n_426),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_457),
.Y(n_550)
);

OR2x6_ASAP7_75t_L g551 ( 
.A(n_526),
.B(n_420),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_461),
.B(n_367),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_466),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_457),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_459),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_467),
.B(n_297),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_457),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_459),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_463),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_531),
.B(n_415),
.Y(n_560)
);

OAI22xp33_ASAP7_75t_SL g561 ( 
.A1(n_499),
.A2(n_378),
.B1(n_445),
.B2(n_397),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_459),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_464),
.Y(n_563)
);

INVx5_ASAP7_75t_L g564 ( 
.A(n_479),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_466),
.B(n_371),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_457),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_505),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_464),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_465),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_499),
.A2(n_453),
.B1(n_441),
.B2(n_420),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_529),
.B(n_409),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_478),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_457),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_457),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_459),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_465),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_473),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_469),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_469),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_473),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_505),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_473),
.Y(n_582)
);

AND2x6_ASAP7_75t_L g583 ( 
.A(n_529),
.B(n_260),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_478),
.B(n_494),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_470),
.Y(n_585)
);

BUFx4f_ASAP7_75t_L g586 ( 
.A(n_479),
.Y(n_586)
);

CKINVDCx16_ASAP7_75t_R g587 ( 
.A(n_533),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_529),
.B(n_380),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_507),
.B(n_260),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_458),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_470),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_531),
.B(n_441),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_494),
.B(n_374),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_472),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_473),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_474),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_467),
.B(n_297),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_505),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_474),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_524),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_457),
.Y(n_601)
);

CKINVDCx14_ASAP7_75t_R g602 ( 
.A(n_533),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_523),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_467),
.B(n_311),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_474),
.Y(n_605)
);

NAND3xp33_ASAP7_75t_L g606 ( 
.A(n_511),
.B(n_379),
.C(n_377),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_462),
.A2(n_389),
.B1(n_373),
.B2(n_385),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_467),
.B(n_388),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_467),
.B(n_391),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_475),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_505),
.B(n_311),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_514),
.B(n_392),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_475),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_523),
.B(n_445),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_475),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_514),
.B(n_403),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_523),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_472),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_477),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_477),
.Y(n_620)
);

INVx4_ASAP7_75t_SL g621 ( 
.A(n_479),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_471),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_514),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_490),
.B(n_314),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_524),
.B(n_407),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_SL g626 ( 
.A(n_507),
.B(n_239),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_484),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_507),
.B(n_408),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_482),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_504),
.B(n_411),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_482),
.B(n_430),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_504),
.B(n_416),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_490),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_483),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_483),
.B(n_423),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_485),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_504),
.B(n_424),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_484),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_458),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_462),
.A2(n_455),
.B1(n_450),
.B2(n_449),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_485),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_SL g642 ( 
.A1(n_458),
.A2(n_402),
.B1(n_405),
.B2(n_421),
.Y(n_642)
);

INVx4_ASAP7_75t_SL g643 ( 
.A(n_479),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_484),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_476),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_471),
.Y(n_646)
);

AND2x6_ASAP7_75t_L g647 ( 
.A(n_504),
.B(n_260),
.Y(n_647)
);

CKINVDCx6p67_ASAP7_75t_R g648 ( 
.A(n_458),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_495),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_486),
.B(n_425),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_476),
.Y(n_651)
);

NAND2x1_ASAP7_75t_L g652 ( 
.A(n_479),
.B(n_333),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_458),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_476),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_495),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_490),
.B(n_314),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_486),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_490),
.B(n_317),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_500),
.A2(n_448),
.B1(n_446),
.B2(n_444),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_495),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_488),
.Y(n_661)
);

OAI22x1_ASAP7_75t_L g662 ( 
.A1(n_496),
.A2(n_358),
.B1(n_318),
.B2(n_187),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_488),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_489),
.B(n_432),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_489),
.B(n_433),
.Y(n_665)
);

OR2x6_ASAP7_75t_L g666 ( 
.A(n_491),
.B(n_430),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_SL g667 ( 
.A(n_491),
.B(n_412),
.C(n_289),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_493),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_493),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_504),
.B(n_435),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_498),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_490),
.B(n_317),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_471),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_498),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_501),
.Y(n_675)
);

XNOR2xp5_ASAP7_75t_L g676 ( 
.A(n_496),
.B(n_365),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_490),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_500),
.A2(n_385),
.B1(n_339),
.B2(n_332),
.Y(n_678)
);

XOR2x2_ASAP7_75t_SL g679 ( 
.A(n_496),
.B(n_273),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_519),
.B(n_438),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_497),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_490),
.B(n_328),
.Y(n_682)
);

AND2x6_ASAP7_75t_L g683 ( 
.A(n_519),
.B(n_355),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_471),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_497),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_501),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_497),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_468),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_553),
.B(n_572),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_645),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_650),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_596),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_553),
.B(n_439),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_584),
.A2(n_506),
.B(n_480),
.Y(n_694)
);

O2A1O1Ixp5_ASAP7_75t_L g695 ( 
.A1(n_556),
.A2(n_519),
.B(n_328),
.C(n_502),
.Y(n_695)
);

INVx8_ASAP7_75t_L g696 ( 
.A(n_592),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_572),
.B(n_506),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_539),
.B(n_375),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_560),
.B(n_437),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_596),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_650),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_592),
.A2(n_390),
.B1(n_496),
.B2(n_330),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_657),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_586),
.B(n_506),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_608),
.B(n_519),
.Y(n_705)
);

BUFx5_ASAP7_75t_L g706 ( 
.A(n_645),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_609),
.B(n_519),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_651),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_552),
.B(n_565),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_586),
.B(n_506),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_599),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_599),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_593),
.B(n_496),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_623),
.B(n_471),
.Y(n_714)
);

NAND3xp33_ASAP7_75t_L g715 ( 
.A(n_570),
.B(n_204),
.C(n_203),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_605),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_586),
.B(n_506),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_623),
.B(n_612),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_630),
.A2(n_506),
.B(n_480),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_657),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_538),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_616),
.B(n_471),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_540),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_628),
.B(n_208),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_542),
.A2(n_329),
.B1(n_331),
.B2(n_291),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_605),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_571),
.B(n_471),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_571),
.B(n_471),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_635),
.B(n_487),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_664),
.B(n_487),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_537),
.B(n_487),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_651),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_537),
.B(n_487),
.Y(n_733)
);

INVx2_ASAP7_75t_SL g734 ( 
.A(n_665),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_617),
.B(n_503),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_654),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_610),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_537),
.B(n_487),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_610),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_632),
.B(n_506),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_665),
.B(n_211),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_542),
.A2(n_329),
.B1(n_291),
.B2(n_331),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_560),
.B(n_217),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_617),
.B(n_437),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_541),
.B(n_487),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_606),
.B(n_220),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_637),
.B(n_506),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_614),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_654),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_670),
.B(n_355),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_680),
.B(n_355),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_550),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_564),
.B(n_355),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_564),
.B(n_355),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_546),
.B(n_487),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_548),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_559),
.Y(n_757)
);

INVxp33_ASAP7_75t_L g758 ( 
.A(n_614),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_676),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_564),
.B(n_355),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_563),
.B(n_487),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_L g762 ( 
.A(n_607),
.B(n_224),
.C(n_221),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_550),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_556),
.A2(n_480),
.B(n_468),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_568),
.B(n_492),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_564),
.B(n_516),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_564),
.B(n_516),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_613),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_550),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_592),
.A2(n_290),
.B1(n_279),
.B2(n_281),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_551),
.B(n_238),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_613),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_569),
.Y(n_773)
);

NOR2xp67_ASAP7_75t_L g774 ( 
.A(n_640),
.B(n_503),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_615),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_576),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_578),
.B(n_492),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_615),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_551),
.A2(n_592),
.B1(n_666),
.B2(n_631),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_588),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_659),
.B(n_516),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_587),
.B(n_626),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_579),
.Y(n_783)
);

INVxp67_ASAP7_75t_R g784 ( 
.A(n_653),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_627),
.Y(n_785)
);

NOR3xp33_ASAP7_75t_L g786 ( 
.A(n_667),
.B(n_216),
.C(n_240),
.Y(n_786)
);

NOR2xp67_ASAP7_75t_L g787 ( 
.A(n_549),
.B(n_508),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_588),
.Y(n_788)
);

OAI221xp5_ASAP7_75t_L g789 ( 
.A1(n_603),
.A2(n_334),
.B1(n_348),
.B2(n_327),
.C(n_345),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_627),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_585),
.B(n_492),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_638),
.Y(n_792)
);

AOI221xp5_ASAP7_75t_L g793 ( 
.A1(n_536),
.A2(n_280),
.B1(n_275),
.B2(n_327),
.C(n_332),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_543),
.A2(n_357),
.B1(n_213),
.B2(n_230),
.Y(n_794)
);

AO22x2_ASAP7_75t_L g795 ( 
.A1(n_679),
.A2(n_543),
.B1(n_600),
.B2(n_611),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_600),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_591),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_551),
.B(n_243),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_594),
.B(n_492),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_638),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_618),
.B(n_492),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_631),
.B(n_508),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_619),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_621),
.B(n_516),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_550),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_644),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_620),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_621),
.B(n_516),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_629),
.B(n_492),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_L g810 ( 
.A(n_589),
.B(n_479),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_644),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_L g812 ( 
.A(n_589),
.B(n_479),
.Y(n_812)
);

NAND3xp33_ASAP7_75t_L g813 ( 
.A(n_626),
.B(n_551),
.C(n_631),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_621),
.B(n_516),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_625),
.B(n_244),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_634),
.B(n_492),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_621),
.B(n_643),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_676),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_636),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_550),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_561),
.B(n_247),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_641),
.B(n_492),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_649),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_661),
.B(n_468),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_643),
.B(n_516),
.Y(n_825)
);

AO22x2_ASAP7_75t_L g826 ( 
.A1(n_679),
.A2(n_357),
.B1(n_202),
.B2(n_285),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_663),
.B(n_468),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_631),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_668),
.B(n_468),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_643),
.B(n_516),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_669),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_649),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_671),
.B(n_480),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_674),
.A2(n_305),
.B1(n_285),
.B2(n_269),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_655),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_655),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_675),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_686),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_643),
.B(n_532),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_545),
.B(n_480),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_545),
.B(n_554),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_666),
.B(n_602),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_688),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_684),
.B(n_532),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_545),
.B(n_481),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_666),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_660),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_554),
.B(n_481),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_688),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_554),
.B(n_481),
.Y(n_850)
);

BUFx8_ASAP7_75t_L g851 ( 
.A(n_590),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_611),
.A2(n_305),
.B1(n_269),
.B2(n_265),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_660),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_681),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_666),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_681),
.Y(n_856)
);

NAND2x1_ASAP7_75t_L g857 ( 
.A(n_566),
.B(n_333),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_685),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_685),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_687),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_602),
.B(n_250),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_692),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_722),
.A2(n_652),
.B(n_574),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_709),
.A2(n_536),
.B1(n_678),
.B2(n_598),
.Y(n_864)
);

OAI21xp33_ASAP7_75t_L g865 ( 
.A1(n_743),
.A2(n_662),
.B(n_642),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_729),
.A2(n_574),
.B(n_557),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_689),
.B(n_566),
.Y(n_867)
);

AO21x1_ASAP7_75t_L g868 ( 
.A1(n_781),
.A2(n_604),
.B(n_597),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_793),
.A2(n_334),
.B(n_275),
.C(n_349),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_692),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_748),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_727),
.A2(n_728),
.B(n_695),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_735),
.Y(n_873)
);

OR2x6_ASAP7_75t_L g874 ( 
.A(n_696),
.B(n_544),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_780),
.B(n_566),
.Y(n_875)
);

NOR2xp67_ASAP7_75t_L g876 ( 
.A(n_813),
.B(n_639),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_730),
.A2(n_574),
.B(n_557),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_700),
.Y(n_878)
);

NOR2x1_ASAP7_75t_L g879 ( 
.A(n_713),
.B(n_544),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_735),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_731),
.A2(n_574),
.B(n_557),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_718),
.A2(n_597),
.B(n_604),
.C(n_672),
.Y(n_882)
);

INVx11_ASAP7_75t_L g883 ( 
.A(n_851),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_779),
.B(n_639),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_735),
.B(n_573),
.Y(n_885)
);

NOR2x1_ASAP7_75t_L g886 ( 
.A(n_693),
.B(n_567),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_711),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_690),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_690),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_721),
.Y(n_890)
);

NAND2x1_ASAP7_75t_L g891 ( 
.A(n_690),
.B(n_573),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_733),
.A2(n_622),
.B(n_557),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_744),
.B(n_648),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_724),
.B(n_601),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_758),
.B(n_648),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_738),
.A2(n_673),
.B(n_622),
.Y(n_896)
);

BUFx4f_ASAP7_75t_L g897 ( 
.A(n_696),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_788),
.B(n_601),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_714),
.A2(n_747),
.B(n_740),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_781),
.A2(n_646),
.B(n_601),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_723),
.B(n_646),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_706),
.B(n_684),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_706),
.B(n_684),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_734),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_740),
.A2(n_673),
.B(n_622),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_747),
.A2(n_673),
.B(n_622),
.Y(n_906)
);

AOI21x1_ASAP7_75t_L g907 ( 
.A1(n_697),
.A2(n_656),
.B(n_624),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_756),
.B(n_646),
.Y(n_908)
);

NAND3xp33_ASAP7_75t_L g909 ( 
.A(n_741),
.B(n_261),
.C(n_256),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_711),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_712),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_773),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_776),
.B(n_783),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_705),
.A2(n_558),
.B(n_555),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_707),
.A2(n_841),
.B(n_697),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_694),
.A2(n_558),
.B(n_555),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_763),
.A2(n_673),
.B(n_684),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_706),
.B(n_690),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_699),
.B(n_662),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_763),
.A2(n_481),
.B(n_547),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_706),
.B(n_567),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_763),
.A2(n_633),
.B(n_547),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_757),
.B(n_581),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_803),
.B(n_687),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_769),
.A2(n_633),
.B(n_547),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_807),
.B(n_562),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_819),
.B(n_562),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_769),
.A2(n_677),
.B(n_633),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_691),
.B(n_581),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_840),
.A2(n_577),
.B(n_575),
.Y(n_930)
);

CKINVDCx10_ASAP7_75t_R g931 ( 
.A(n_759),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_736),
.A2(n_598),
.B1(n_265),
.B2(n_213),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_712),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_818),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_831),
.B(n_837),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_838),
.B(n_703),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_802),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_769),
.A2(n_677),
.B(n_656),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_720),
.B(n_575),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_769),
.A2(n_677),
.B(n_658),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_701),
.B(n_758),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_757),
.B(n_797),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_843),
.Y(n_943)
);

AOI21xp33_ASAP7_75t_L g944 ( 
.A1(n_746),
.A2(n_230),
.B(n_202),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_846),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_706),
.B(n_577),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_797),
.B(n_774),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_820),
.A2(n_658),
.B(n_624),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_698),
.B(n_796),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_736),
.A2(n_236),
.B1(n_257),
.B2(n_258),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_828),
.B(n_771),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_846),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_736),
.B(n_580),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_706),
.B(n_580),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_708),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_845),
.A2(n_595),
.B(n_582),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_749),
.B(n_582),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_706),
.B(n_595),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_798),
.B(n_266),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_749),
.B(n_589),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_820),
.A2(n_682),
.B(n_672),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_787),
.B(n_589),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_716),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_789),
.A2(n_682),
.B(n_236),
.C(n_257),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_782),
.B(n_509),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_815),
.B(n_589),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_855),
.B(n_509),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_820),
.A2(n_510),
.B(n_522),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_715),
.B(n_513),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_SL g970 ( 
.A1(n_842),
.A2(n_821),
.B1(n_702),
.B2(n_855),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_716),
.Y(n_971)
);

AOI21x1_ASAP7_75t_L g972 ( 
.A1(n_844),
.A2(n_502),
.B(n_522),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_726),
.B(n_583),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_726),
.B(n_583),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_848),
.A2(n_583),
.B(n_647),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_708),
.Y(n_976)
);

OAI21xp33_ASAP7_75t_SL g977 ( 
.A1(n_852),
.A2(n_751),
.B(n_750),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_737),
.B(n_583),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_737),
.B(n_583),
.Y(n_979)
);

AOI21x1_ASAP7_75t_L g980 ( 
.A1(n_844),
.A2(n_502),
.B(n_522),
.Y(n_980)
);

INVx11_ASAP7_75t_L g981 ( 
.A(n_851),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_820),
.A2(n_522),
.B(n_510),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_850),
.A2(n_510),
.B(n_534),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_745),
.A2(n_510),
.B(n_534),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_739),
.B(n_583),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_708),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_739),
.B(n_258),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_708),
.B(n_532),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_732),
.A2(n_302),
.B1(n_347),
.B2(n_343),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_755),
.A2(n_534),
.B(n_532),
.Y(n_990)
);

BUFx8_ASAP7_75t_SL g991 ( 
.A(n_851),
.Y(n_991)
);

CKINVDCx10_ASAP7_75t_R g992 ( 
.A(n_861),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_761),
.A2(n_534),
.B(n_532),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_696),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_765),
.A2(n_532),
.B(n_515),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_777),
.A2(n_532),
.B(n_515),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_795),
.A2(n_350),
.B1(n_287),
.B2(n_292),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_791),
.A2(n_532),
.B(n_517),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_799),
.A2(n_513),
.B(n_517),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_696),
.A2(n_762),
.B(n_794),
.C(n_742),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_750),
.A2(n_521),
.B(n_518),
.C(n_530),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_801),
.A2(n_518),
.B(n_521),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_809),
.A2(n_683),
.B(n_647),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_768),
.B(n_535),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_751),
.A2(n_525),
.B(n_527),
.C(n_530),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_786),
.B(n_525),
.Y(n_1006)
);

AO21x1_ASAP7_75t_L g1007 ( 
.A1(n_816),
.A2(n_822),
.B(n_857),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_849),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_824),
.A2(n_527),
.B(n_528),
.C(n_349),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_770),
.B(n_272),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_704),
.A2(n_528),
.B(n_535),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_704),
.A2(n_535),
.B(n_326),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_732),
.A2(n_335),
.B1(n_325),
.B2(n_337),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_784),
.B(n_283),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_732),
.B(n_817),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_768),
.B(n_535),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_710),
.A2(n_717),
.B(n_719),
.Y(n_1017)
);

AOI33xp33_ASAP7_75t_L g1018 ( 
.A1(n_834),
.A2(n_339),
.A3(n_345),
.B1(n_344),
.B2(n_338),
.B3(n_348),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_732),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_772),
.B(n_535),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_827),
.B(n_276),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_795),
.A2(n_324),
.B1(n_299),
.B2(n_312),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_829),
.B(n_833),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_853),
.B(n_282),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_764),
.B(n_351),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_710),
.A2(n_323),
.B(n_296),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_772),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_717),
.A2(n_313),
.B(n_360),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_752),
.A2(n_387),
.B(n_383),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_858),
.B(n_284),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_775),
.B(n_683),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_826),
.B(n_283),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_795),
.A2(n_294),
.B1(n_286),
.B2(n_288),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_775),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_778),
.A2(n_683),
.B(n_647),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_SL g1036 ( 
.A(n_859),
.B(n_207),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_785),
.B(n_293),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_826),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_752),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_752),
.A2(n_387),
.B(n_383),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_785),
.B(n_683),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_810),
.A2(n_338),
.B(n_344),
.C(n_207),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_805),
.A2(n_479),
.B(n_683),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_826),
.B(n_283),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_790),
.B(n_792),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_790),
.B(n_647),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_792),
.Y(n_1047)
);

NOR2x1_ASAP7_75t_L g1048 ( 
.A(n_817),
.B(n_231),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_725),
.B(n_298),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_959),
.A2(n_860),
.B(n_856),
.C(n_854),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_931),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_888),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_944),
.A2(n_860),
.B(n_856),
.C(n_854),
.Y(n_1053)
);

NAND2xp33_ASAP7_75t_SL g1054 ( 
.A(n_893),
.B(n_804),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_949),
.B(n_800),
.Y(n_1055)
);

INVx5_ASAP7_75t_L g1056 ( 
.A(n_888),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_864),
.B(n_949),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_942),
.B(n_805),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_959),
.A2(n_847),
.B(n_800),
.C(n_836),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_894),
.A2(n_812),
.B(n_810),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_890),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_873),
.A2(n_847),
.B1(n_806),
.B2(n_836),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_912),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_937),
.B(n_951),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_918),
.A2(n_812),
.B(n_808),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_880),
.B(n_806),
.Y(n_1066)
);

NOR2xp67_ASAP7_75t_L g1067 ( 
.A(n_909),
.B(n_811),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_937),
.B(n_811),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_945),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_913),
.B(n_935),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1021),
.B(n_823),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1021),
.B(n_823),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_971),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_947),
.B(n_832),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_951),
.B(n_300),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_L g1076 ( 
.A(n_865),
.B(n_356),
.C(n_301),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_936),
.B(n_832),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_R g1078 ( 
.A(n_934),
.B(n_68),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_1010),
.A2(n_835),
.B(n_839),
.C(n_830),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_965),
.B(n_835),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_1015),
.B(n_804),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_1010),
.A2(n_839),
.B(n_830),
.C(n_825),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_923),
.B(n_231),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_971),
.Y(n_1084)
);

NAND3xp33_ASAP7_75t_L g1085 ( 
.A(n_869),
.B(n_941),
.C(n_997),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_994),
.B(n_808),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1037),
.B(n_814),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_923),
.B(n_231),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_1038),
.B(n_814),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1015),
.A2(n_825),
.B1(n_760),
.B2(n_754),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_977),
.A2(n_760),
.B(n_754),
.C(n_753),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_952),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_888),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_902),
.A2(n_903),
.B(n_863),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1034),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_862),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_866),
.A2(n_767),
.B(n_766),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1037),
.B(n_766),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_871),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_870),
.Y(n_1100)
);

OA22x2_ASAP7_75t_L g1101 ( 
.A1(n_1032),
.A2(n_303),
.B1(n_304),
.B2(n_307),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_926),
.Y(n_1102)
);

AOI21x1_ASAP7_75t_L g1103 ( 
.A1(n_921),
.A2(n_767),
.B(n_753),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_904),
.B(n_231),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_994),
.B(n_118),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_991),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_919),
.B(n_309),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1044),
.B(n_310),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_927),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1024),
.B(n_352),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_991),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_871),
.B(n_315),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_877),
.A2(n_479),
.B(n_108),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_897),
.A2(n_364),
.B1(n_362),
.B2(n_361),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1022),
.A2(n_882),
.B(n_969),
.C(n_1000),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1000),
.A2(n_359),
.B(n_354),
.C(n_353),
.Y(n_1116)
);

AO32x1_ASAP7_75t_L g1117 ( 
.A1(n_950),
.A2(n_351),
.A3(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1014),
.B(n_321),
.Y(n_1118)
);

AOI21x1_ASAP7_75t_L g1119 ( 
.A1(n_921),
.A2(n_351),
.B(n_80),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1006),
.B(n_322),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1024),
.B(n_346),
.Y(n_1121)
);

HB1xp67_ASAP7_75t_L g1122 ( 
.A(n_888),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_878),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_889),
.B(n_351),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1030),
.B(n_342),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_884),
.B(n_15),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_915),
.A2(n_182),
.B(n_176),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_967),
.Y(n_1128)
);

BUFx12f_ASAP7_75t_L g1129 ( 
.A(n_967),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_SL g1130 ( 
.A(n_897),
.B(n_172),
.Y(n_1130)
);

CKINVDCx10_ASAP7_75t_R g1131 ( 
.A(n_883),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_929),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_872),
.A2(n_163),
.B(n_157),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_889),
.B(n_152),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_869),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_884),
.B(n_22),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_924),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_887),
.Y(n_1138)
);

AOI22x1_ASAP7_75t_L g1139 ( 
.A1(n_1017),
.A2(n_146),
.B1(n_145),
.B2(n_141),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_899),
.A2(n_138),
.B(n_137),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_970),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_867),
.B(n_23),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_992),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_889),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_SL g1145 ( 
.A1(n_895),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_895),
.B(n_28),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1049),
.B(n_29),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_881),
.A2(n_136),
.B(n_124),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_972),
.A2(n_117),
.B(n_110),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_876),
.A2(n_30),
.B(n_31),
.C(n_33),
.Y(n_1150)
);

INVxp67_ASAP7_75t_SL g1151 ( 
.A(n_889),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_955),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_955),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_966),
.A2(n_37),
.B(n_39),
.C(n_41),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1033),
.B(n_44),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_910),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_955),
.B(n_103),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_911),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_933),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_943),
.B(n_44),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_963),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1008),
.B(n_49),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_892),
.A2(n_98),
.B(n_82),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1042),
.A2(n_49),
.B(n_51),
.C(n_55),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_1019),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1036),
.B(n_55),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_964),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_1167)
);

OR2x6_ASAP7_75t_L g1168 ( 
.A(n_874),
.B(n_57),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_896),
.A2(n_58),
.B(n_60),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_955),
.B(n_60),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1011),
.A2(n_962),
.B(n_1002),
.C(n_999),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_976),
.B(n_886),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1027),
.B(n_1047),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_953),
.A2(n_957),
.B(n_960),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_932),
.A2(n_1009),
.B(n_1005),
.C(n_1001),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_885),
.A2(n_900),
.B(n_875),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_868),
.A2(n_987),
.B1(n_939),
.B2(n_901),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1045),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1018),
.B(n_1048),
.Y(n_1179)
);

NAND2xp33_ASAP7_75t_SL g1180 ( 
.A(n_976),
.B(n_1019),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_989),
.A2(n_1013),
.B(n_898),
.C(n_908),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_986),
.B(n_976),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_976),
.B(n_1018),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_879),
.B(n_1039),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_981),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_874),
.A2(n_1039),
.B1(n_974),
.B2(n_973),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1023),
.A2(n_1025),
.B(n_1040),
.C(n_1029),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_946),
.A2(n_958),
.B(n_954),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1004),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1023),
.B(n_1016),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_874),
.Y(n_1191)
);

BUFx4f_ASAP7_75t_L g1192 ( 
.A(n_891),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_954),
.A2(n_917),
.B(n_906),
.Y(n_1193)
);

AO21x2_ASAP7_75t_L g1194 ( 
.A1(n_1007),
.A2(n_916),
.B(n_914),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_1025),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1020),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_980),
.A2(n_905),
.B(n_956),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_907),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_995),
.B(n_996),
.Y(n_1199)
);

NOR2x1_ASAP7_75t_L g1200 ( 
.A(n_988),
.B(n_1026),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_998),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_988),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1031),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_948),
.B(n_961),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_938),
.A2(n_940),
.B(n_922),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1041),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1028),
.A2(n_985),
.B1(n_979),
.B2(n_978),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1046),
.A2(n_975),
.B1(n_1003),
.B2(n_930),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1043),
.Y(n_1209)
);

OA21x2_ASAP7_75t_L g1210 ( 
.A1(n_1177),
.A2(n_990),
.B(n_993),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1095),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1069),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1205),
.A2(n_1072),
.B(n_1071),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_1092),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1070),
.B(n_984),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1094),
.A2(n_925),
.B(n_928),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1061),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1115),
.A2(n_1171),
.A3(n_1116),
.B(n_1198),
.Y(n_1218)
);

AOI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_1057),
.A2(n_983),
.B(n_1035),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1057),
.A2(n_968),
.B(n_982),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1075),
.B(n_1012),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1084),
.Y(n_1222)
);

INVx1_ASAP7_75t_SL g1223 ( 
.A(n_1099),
.Y(n_1223)
);

INVx8_ASAP7_75t_L g1224 ( 
.A(n_1056),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1050),
.A2(n_920),
.A3(n_1059),
.B(n_1091),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1137),
.B(n_1102),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1063),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1199),
.A2(n_1204),
.B(n_1087),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1098),
.A2(n_1174),
.B(n_1194),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1082),
.A2(n_1079),
.A3(n_1186),
.B(n_1193),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1099),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1120),
.A2(n_1146),
.B(n_1076),
.C(n_1126),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1194),
.A2(n_1176),
.B(n_1060),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1112),
.Y(n_1234)
);

INVx5_ASAP7_75t_L g1235 ( 
.A(n_1052),
.Y(n_1235)
);

A2O1A1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1120),
.A2(n_1146),
.B(n_1076),
.C(n_1136),
.Y(n_1236)
);

AO21x2_ASAP7_75t_L g1237 ( 
.A1(n_1133),
.A2(n_1142),
.B(n_1188),
.Y(n_1237)
);

OAI221xp5_ASAP7_75t_L g1238 ( 
.A1(n_1141),
.A2(n_1110),
.B1(n_1125),
.B2(n_1121),
.C(n_1136),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1096),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1159),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1201),
.A2(n_1062),
.A3(n_1164),
.B(n_1154),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1155),
.A2(n_1126),
.B(n_1150),
.C(n_1104),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1108),
.B(n_1118),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1064),
.B(n_1080),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1100),
.Y(n_1245)
);

NOR2xp67_ASAP7_75t_L g1246 ( 
.A(n_1056),
.B(n_1085),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1181),
.A2(n_1177),
.B(n_1190),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1064),
.B(n_1080),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1123),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1149),
.A2(n_1103),
.B(n_1097),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1109),
.B(n_1178),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1132),
.B(n_1112),
.Y(n_1252)
);

AO31x2_ASAP7_75t_L g1253 ( 
.A1(n_1155),
.A2(n_1127),
.A3(n_1090),
.B(n_1169),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1208),
.A2(n_1207),
.B(n_1187),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1119),
.A2(n_1065),
.B(n_1200),
.Y(n_1255)
);

AO31x2_ASAP7_75t_L g1256 ( 
.A1(n_1089),
.A2(n_1140),
.A3(n_1183),
.B(n_1074),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1208),
.A2(n_1054),
.B(n_1077),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1052),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1055),
.B(n_1147),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1191),
.B(n_1128),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1058),
.A2(n_1053),
.B(n_1151),
.Y(n_1261)
);

OAI21xp33_ASAP7_75t_L g1262 ( 
.A1(n_1160),
.A2(n_1162),
.B(n_1166),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1151),
.A2(n_1175),
.B(n_1081),
.Y(n_1263)
);

AOI221xp5_ASAP7_75t_L g1264 ( 
.A1(n_1145),
.A2(n_1135),
.B1(n_1107),
.B2(n_1162),
.C(n_1160),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1089),
.A2(n_1067),
.B(n_1179),
.C(n_1167),
.Y(n_1265)
);

AOI221xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1170),
.A2(n_1068),
.B1(n_1195),
.B2(n_1124),
.C(n_1081),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1129),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1068),
.B(n_1196),
.Y(n_1268)
);

INVx3_ASAP7_75t_SL g1269 ( 
.A(n_1051),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1209),
.A2(n_1113),
.B(n_1189),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1111),
.Y(n_1271)
);

AOI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1172),
.A2(n_1184),
.B(n_1124),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1114),
.B(n_1088),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1138),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1185),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1139),
.A2(n_1148),
.B(n_1163),
.Y(n_1276)
);

AOI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1066),
.A2(n_1134),
.B(n_1157),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1156),
.B(n_1158),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1052),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1122),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1105),
.Y(n_1281)
);

AOI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1170),
.A2(n_1101),
.B1(n_1130),
.B2(n_1202),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1105),
.B(n_1086),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1101),
.B(n_1078),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1056),
.Y(n_1285)
);

INVx4_ASAP7_75t_L g1286 ( 
.A(n_1056),
.Y(n_1286)
);

AO21x1_ASAP7_75t_L g1287 ( 
.A1(n_1134),
.A2(n_1157),
.B(n_1182),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1168),
.A2(n_1078),
.B1(n_1106),
.B2(n_1086),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_1143),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1083),
.A2(n_1192),
.B(n_1203),
.C(n_1182),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1161),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1180),
.A2(n_1192),
.B(n_1173),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1168),
.B(n_1144),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1165),
.Y(n_1294)
);

NAND3x1_ASAP7_75t_L g1295 ( 
.A(n_1131),
.B(n_1168),
.C(n_1165),
.Y(n_1295)
);

AO31x2_ASAP7_75t_L g1296 ( 
.A1(n_1117),
.A2(n_1206),
.A3(n_1122),
.B(n_1093),
.Y(n_1296)
);

OAI22x1_ASAP7_75t_L g1297 ( 
.A1(n_1117),
.A2(n_1206),
.B1(n_1093),
.B2(n_1152),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1052),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1206),
.A2(n_1117),
.B(n_1093),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1153),
.B(n_1093),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1152),
.B(n_1153),
.Y(n_1301)
);

AOI221x1_ASAP7_75t_L g1302 ( 
.A1(n_1152),
.A2(n_1153),
.B1(n_944),
.B2(n_1155),
.C(n_1136),
.Y(n_1302)
);

CKINVDCx11_ASAP7_75t_R g1303 ( 
.A(n_1111),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1061),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1205),
.A2(n_894),
.B(n_1071),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1057),
.A2(n_1126),
.B1(n_1136),
.B2(n_1155),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1057),
.A2(n_709),
.B(n_959),
.C(n_865),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1115),
.A2(n_1057),
.B(n_1116),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1070),
.B(n_709),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1115),
.A2(n_868),
.A3(n_1007),
.B(n_1171),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1205),
.A2(n_894),
.B(n_1071),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1131),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1070),
.B(n_709),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1177),
.A2(n_1115),
.B(n_1197),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1073),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1075),
.B(n_1108),
.Y(n_1316)
);

AO31x2_ASAP7_75t_L g1317 ( 
.A1(n_1115),
.A2(n_868),
.A3(n_1007),
.B(n_1171),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1075),
.B(n_1108),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1064),
.B(n_365),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1070),
.B(n_699),
.Y(n_1320)
);

AO32x2_ASAP7_75t_L g1321 ( 
.A1(n_1145),
.A2(n_1038),
.A3(n_970),
.B1(n_1033),
.B2(n_950),
.Y(n_1321)
);

BUFx8_ASAP7_75t_SL g1322 ( 
.A(n_1051),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1069),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1052),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1056),
.B(n_1019),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1070),
.B(n_709),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1205),
.A2(n_1193),
.B(n_1094),
.Y(n_1327)
);

A2O1A1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1057),
.A2(n_709),
.B(n_959),
.C(n_865),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1205),
.A2(n_1193),
.B(n_1094),
.Y(n_1329)
);

NAND3xp33_ASAP7_75t_L g1330 ( 
.A(n_1057),
.B(n_959),
.C(n_944),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1205),
.A2(n_1193),
.B(n_1094),
.Y(n_1331)
);

BUFx2_ASAP7_75t_SL g1332 ( 
.A(n_1069),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1073),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1205),
.A2(n_894),
.B(n_1071),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1205),
.A2(n_1193),
.B(n_1094),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1205),
.A2(n_1193),
.B(n_1094),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1191),
.B(n_994),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1205),
.A2(n_894),
.B(n_1071),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1115),
.A2(n_1057),
.B(n_1116),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1205),
.A2(n_1193),
.B(n_1094),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1070),
.B(n_709),
.Y(n_1341)
);

NOR3xp33_ASAP7_75t_L g1342 ( 
.A(n_1120),
.B(n_959),
.C(n_698),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1205),
.A2(n_1193),
.B(n_1094),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1061),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1070),
.B(n_709),
.Y(n_1345)
);

AOI31xp67_ASAP7_75t_L g1346 ( 
.A1(n_1057),
.A2(n_750),
.A3(n_751),
.B(n_1199),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_SL g1347 ( 
.A1(n_1115),
.A2(n_1082),
.B(n_1057),
.C(n_1116),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1205),
.A2(n_1193),
.B(n_1094),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1205),
.A2(n_1193),
.B(n_1094),
.Y(n_1349)
);

INVxp67_ASAP7_75t_SL g1350 ( 
.A(n_1099),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1052),
.Y(n_1351)
);

INVx3_ASAP7_75t_SL g1352 ( 
.A(n_1051),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1205),
.A2(n_894),
.B(n_1071),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1205),
.A2(n_894),
.B(n_1071),
.Y(n_1354)
);

NOR2xp67_ASAP7_75t_L g1355 ( 
.A(n_1070),
.B(n_947),
.Y(n_1355)
);

AO31x2_ASAP7_75t_L g1356 ( 
.A1(n_1115),
.A2(n_868),
.A3(n_1007),
.B(n_1171),
.Y(n_1356)
);

AO21x2_ASAP7_75t_L g1357 ( 
.A1(n_1115),
.A2(n_1194),
.B(n_1057),
.Y(n_1357)
);

AO32x2_ASAP7_75t_L g1358 ( 
.A1(n_1145),
.A2(n_1038),
.A3(n_970),
.B1(n_1033),
.B2(n_950),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_1099),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1191),
.B(n_994),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1070),
.B(n_709),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1191),
.B(n_994),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1238),
.A2(n_1330),
.B1(n_1319),
.B2(n_1313),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1212),
.Y(n_1364)
);

OAI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1306),
.A2(n_1361),
.B1(n_1309),
.B2(n_1326),
.Y(n_1365)
);

CKINVDCx11_ASAP7_75t_R g1366 ( 
.A(n_1269),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1342),
.A2(n_1306),
.B1(n_1264),
.B2(n_1262),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1330),
.A2(n_1345),
.B1(n_1341),
.B2(n_1273),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1322),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1214),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1262),
.A2(n_1345),
.B1(n_1341),
.B2(n_1308),
.Y(n_1371)
);

OR2x2_ASAP7_75t_L g1372 ( 
.A(n_1320),
.B(n_1259),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1224),
.Y(n_1373)
);

OAI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1244),
.A2(n_1248),
.B1(n_1282),
.B2(n_1234),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1303),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1308),
.A2(n_1339),
.B1(n_1282),
.B2(n_1254),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1227),
.Y(n_1377)
);

BUFx8_ASAP7_75t_L g1378 ( 
.A(n_1323),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1316),
.B(n_1318),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1232),
.A2(n_1236),
.B1(n_1252),
.B2(n_1307),
.Y(n_1380)
);

INVx2_ASAP7_75t_SL g1381 ( 
.A(n_1275),
.Y(n_1381)
);

BUFx4f_ASAP7_75t_SL g1382 ( 
.A(n_1289),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_SL g1383 ( 
.A1(n_1339),
.A2(n_1284),
.B1(n_1254),
.B2(n_1358),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1321),
.A2(n_1358),
.B1(n_1357),
.B2(n_1268),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1304),
.Y(n_1385)
);

INVx6_ASAP7_75t_L g1386 ( 
.A(n_1224),
.Y(n_1386)
);

CKINVDCx11_ASAP7_75t_R g1387 ( 
.A(n_1352),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1283),
.B(n_1281),
.Y(n_1388)
);

OAI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1268),
.A2(n_1226),
.B1(n_1302),
.B2(n_1251),
.Y(n_1389)
);

OAI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1328),
.A2(n_1242),
.B(n_1355),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1355),
.A2(n_1247),
.B1(n_1357),
.B2(n_1226),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_SL g1392 ( 
.A1(n_1288),
.A2(n_1243),
.B(n_1265),
.Y(n_1392)
);

OAI21xp33_ASAP7_75t_L g1393 ( 
.A1(n_1221),
.A2(n_1223),
.B(n_1350),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1283),
.A2(n_1287),
.B1(n_1240),
.B2(n_1344),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1223),
.B(n_1231),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1293),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1245),
.A2(n_1274),
.B1(n_1249),
.B2(n_1263),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1321),
.A2(n_1358),
.B1(n_1314),
.B2(n_1332),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1237),
.A2(n_1215),
.B1(n_1314),
.B2(n_1246),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1267),
.Y(n_1400)
);

BUFx2_ASAP7_75t_L g1401 ( 
.A(n_1359),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1260),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_1260),
.Y(n_1403)
);

CKINVDCx11_ASAP7_75t_R g1404 ( 
.A(n_1271),
.Y(n_1404)
);

CKINVDCx11_ASAP7_75t_R g1405 ( 
.A(n_1337),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1295),
.A2(n_1266),
.B1(n_1246),
.B2(n_1347),
.Y(n_1406)
);

INVx5_ASAP7_75t_L g1407 ( 
.A(n_1285),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1237),
.A2(n_1291),
.B1(n_1257),
.B2(n_1228),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1266),
.B(n_1280),
.Y(n_1409)
);

CKINVDCx11_ASAP7_75t_R g1410 ( 
.A(n_1337),
.Y(n_1410)
);

BUFx8_ASAP7_75t_L g1411 ( 
.A(n_1360),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1321),
.B(n_1360),
.Y(n_1412)
);

INVx4_ASAP7_75t_SL g1413 ( 
.A(n_1258),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1222),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1278),
.B(n_1290),
.Y(n_1415)
);

INVx6_ASAP7_75t_L g1416 ( 
.A(n_1235),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1299),
.A2(n_1210),
.B1(n_1233),
.B2(n_1362),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1211),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1298),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1315),
.Y(n_1420)
);

OAI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1333),
.A2(n_1297),
.B1(n_1294),
.B2(n_1299),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1300),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1312),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1301),
.B(n_1279),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1272),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1258),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1210),
.A2(n_1276),
.B1(n_1286),
.B2(n_1235),
.Y(n_1427)
);

OAI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1261),
.A2(n_1235),
.B1(n_1277),
.B2(n_1292),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1279),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1324),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_SL g1431 ( 
.A1(n_1213),
.A2(n_1229),
.B1(n_1220),
.B2(n_1270),
.Y(n_1431)
);

INVx2_ASAP7_75t_SL g1432 ( 
.A(n_1324),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1218),
.B(n_1351),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1351),
.Y(n_1434)
);

INVx5_ASAP7_75t_L g1435 ( 
.A(n_1351),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1325),
.Y(n_1436)
);

CKINVDCx11_ASAP7_75t_R g1437 ( 
.A(n_1256),
.Y(n_1437)
);

INVx3_ASAP7_75t_SL g1438 ( 
.A(n_1346),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1256),
.B(n_1354),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1241),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_SL g1441 ( 
.A1(n_1270),
.A2(n_1220),
.B1(n_1253),
.B2(n_1241),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1241),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1255),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1310),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1219),
.A2(n_1305),
.B1(n_1353),
.B2(n_1334),
.Y(n_1445)
);

OAI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1311),
.A2(n_1338),
.B1(n_1253),
.B2(n_1216),
.Y(n_1446)
);

BUFx10_ASAP7_75t_L g1447 ( 
.A(n_1253),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1317),
.B(n_1356),
.Y(n_1448)
);

INVx8_ASAP7_75t_L g1449 ( 
.A(n_1327),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1329),
.A2(n_1336),
.B1(n_1340),
.B2(n_1343),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_SL g1451 ( 
.A1(n_1331),
.A2(n_1335),
.B1(n_1349),
.B2(n_1348),
.Y(n_1451)
);

BUFx4f_ASAP7_75t_SL g1452 ( 
.A(n_1317),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1225),
.Y(n_1453)
);

BUFx12f_ASAP7_75t_L g1454 ( 
.A(n_1356),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1250),
.A2(n_1230),
.B1(n_1296),
.B2(n_1225),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1230),
.Y(n_1456)
);

AOI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1230),
.A2(n_1342),
.B1(n_959),
.B2(n_1306),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1342),
.A2(n_1306),
.B1(n_1264),
.B2(n_1262),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1224),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1322),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1342),
.A2(n_1306),
.B1(n_1264),
.B2(n_1262),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1224),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1342),
.A2(n_1306),
.B1(n_1264),
.B2(n_1262),
.Y(n_1463)
);

CKINVDCx20_ASAP7_75t_R g1464 ( 
.A(n_1289),
.Y(n_1464)
);

CKINVDCx6p67_ASAP7_75t_R g1465 ( 
.A(n_1269),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1309),
.B(n_1313),
.Y(n_1466)
);

INVx5_ASAP7_75t_L g1467 ( 
.A(n_1224),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1238),
.A2(n_1141),
.B1(n_1145),
.B2(n_536),
.Y(n_1468)
);

BUFx12f_ASAP7_75t_L g1469 ( 
.A(n_1303),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1309),
.A2(n_1313),
.B1(n_1361),
.B2(n_1326),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1238),
.A2(n_1141),
.B1(n_1145),
.B2(n_536),
.Y(n_1471)
);

INVx6_ASAP7_75t_L g1472 ( 
.A(n_1224),
.Y(n_1472)
);

AND2x2_ASAP7_75t_SL g1473 ( 
.A(n_1342),
.B(n_1306),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1342),
.A2(n_1306),
.B1(n_1264),
.B2(n_1262),
.Y(n_1474)
);

BUFx12f_ASAP7_75t_L g1475 ( 
.A(n_1303),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1212),
.Y(n_1476)
);

BUFx4f_ASAP7_75t_L g1477 ( 
.A(n_1269),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1238),
.A2(n_1141),
.B1(n_1145),
.B2(n_536),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1309),
.A2(n_1313),
.B1(n_1361),
.B2(n_1326),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1239),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1214),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1214),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1217),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1444),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1433),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1453),
.B(n_1443),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1379),
.Y(n_1487)
);

OR2x6_ASAP7_75t_L g1488 ( 
.A(n_1449),
.B(n_1454),
.Y(n_1488)
);

AO21x2_ASAP7_75t_L g1489 ( 
.A1(n_1446),
.A2(n_1428),
.B(n_1457),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1450),
.A2(n_1439),
.B(n_1445),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1470),
.B(n_1479),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1412),
.B(n_1383),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1386),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1440),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1442),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1446),
.A2(n_1380),
.B(n_1431),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1370),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1386),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1383),
.B(n_1384),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1448),
.Y(n_1500)
);

CKINVDCx6p67_ASAP7_75t_R g1501 ( 
.A(n_1404),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1425),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1377),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1395),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1390),
.B(n_1456),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1385),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1416),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1473),
.A2(n_1471),
.B1(n_1468),
.B2(n_1478),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1452),
.Y(n_1509)
);

AOI21xp33_ASAP7_75t_L g1510 ( 
.A1(n_1473),
.A2(n_1458),
.B(n_1461),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1422),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1452),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1409),
.B(n_1376),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1384),
.B(n_1398),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_SL g1515 ( 
.A1(n_1468),
.A2(n_1471),
.B1(n_1478),
.B2(n_1461),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1441),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1372),
.B(n_1365),
.Y(n_1517)
);

AO21x2_ASAP7_75t_L g1518 ( 
.A1(n_1428),
.A2(n_1421),
.B(n_1389),
.Y(n_1518)
);

AO21x1_ASAP7_75t_L g1519 ( 
.A1(n_1374),
.A2(n_1389),
.B(n_1421),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1376),
.B(n_1367),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1408),
.A2(n_1399),
.B(n_1455),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1398),
.B(n_1368),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1394),
.B(n_1467),
.Y(n_1523)
);

NOR2x1_ASAP7_75t_R g1524 ( 
.A(n_1387),
.B(n_1375),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1367),
.B(n_1458),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_1416),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1401),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1404),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1396),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1472),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1483),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1447),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1414),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1447),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1437),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1481),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1394),
.B(n_1467),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1455),
.A2(n_1391),
.B(n_1399),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1368),
.B(n_1417),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1437),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1417),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1482),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1391),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1418),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1472),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1463),
.B(n_1474),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1438),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1420),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1438),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1397),
.A2(n_1371),
.B(n_1415),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1392),
.B(n_1466),
.Y(n_1551)
);

INVx5_ASAP7_75t_L g1552 ( 
.A(n_1416),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1463),
.B(n_1474),
.Y(n_1553)
);

NAND2x1p5_ASAP7_75t_L g1554 ( 
.A(n_1467),
.B(n_1407),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1397),
.A2(n_1371),
.B(n_1406),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1424),
.B(n_1363),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1427),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1480),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1427),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1405),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1393),
.B(n_1365),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1431),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1403),
.B(n_1388),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1429),
.B(n_1434),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1402),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_1464),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1388),
.B(n_1426),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1451),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1451),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1432),
.B(n_1430),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1366),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1373),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1472),
.Y(n_1573)
);

AOI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1381),
.A2(n_1364),
.B(n_1435),
.Y(n_1574)
);

BUFx2_ASAP7_75t_SL g1575 ( 
.A(n_1435),
.Y(n_1575)
);

OR2x6_ASAP7_75t_L g1576 ( 
.A(n_1496),
.B(n_1373),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1489),
.A2(n_1435),
.B(n_1436),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1515),
.A2(n_1465),
.B1(n_1387),
.B2(n_1469),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1556),
.B(n_1419),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1556),
.B(n_1511),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1535),
.B(n_1410),
.Y(n_1581)
);

NAND2xp33_ASAP7_75t_R g1582 ( 
.A(n_1528),
.B(n_1369),
.Y(n_1582)
);

A2O1A1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1510),
.A2(n_1477),
.B(n_1400),
.C(n_1459),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1491),
.B(n_1373),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1504),
.B(n_1378),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1535),
.B(n_1476),
.Y(n_1586)
);

OA21x2_ASAP7_75t_L g1587 ( 
.A1(n_1490),
.A2(n_1413),
.B(n_1462),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1536),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1542),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1513),
.B(n_1462),
.Y(n_1590)
);

OAI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1525),
.A2(n_1477),
.B(n_1460),
.Y(n_1591)
);

OR2x6_ASAP7_75t_L g1592 ( 
.A(n_1523),
.B(n_1462),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1513),
.B(n_1517),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1540),
.B(n_1413),
.Y(n_1594)
);

AOI221xp5_ASAP7_75t_L g1595 ( 
.A1(n_1515),
.A2(n_1423),
.B1(n_1411),
.B2(n_1382),
.C(n_1475),
.Y(n_1595)
);

AND2x4_ASAP7_75t_SL g1596 ( 
.A(n_1501),
.B(n_1382),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_R g1597 ( 
.A(n_1566),
.B(n_1411),
.Y(n_1597)
);

AND2x2_ASAP7_75t_SL g1598 ( 
.A(n_1539),
.B(n_1522),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1527),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1553),
.A2(n_1525),
.B1(n_1546),
.B2(n_1508),
.Y(n_1600)
);

AOI221xp5_ASAP7_75t_L g1601 ( 
.A1(n_1551),
.A2(n_1553),
.B1(n_1519),
.B2(n_1562),
.C(n_1539),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1546),
.A2(n_1520),
.B(n_1555),
.Y(n_1602)
);

A2O1A1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1520),
.A2(n_1555),
.B(n_1561),
.C(n_1516),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1562),
.B(n_1522),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1485),
.B(n_1500),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_1529),
.Y(n_1606)
);

A2O1A1Ixp33_ASAP7_75t_L g1607 ( 
.A1(n_1561),
.A2(n_1516),
.B(n_1550),
.C(n_1523),
.Y(n_1607)
);

NAND2x1p5_ASAP7_75t_L g1608 ( 
.A(n_1552),
.B(n_1523),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1540),
.B(n_1487),
.Y(n_1609)
);

O2A1O1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1519),
.A2(n_1565),
.B(n_1518),
.C(n_1489),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1492),
.B(n_1567),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1497),
.B(n_1563),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1550),
.A2(n_1537),
.B(n_1523),
.C(n_1541),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1503),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1492),
.B(n_1506),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1571),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1506),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1560),
.B(n_1501),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1499),
.A2(n_1514),
.B1(n_1541),
.B2(n_1552),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1499),
.A2(n_1514),
.B1(n_1552),
.B2(n_1543),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1552),
.A2(n_1543),
.B1(n_1557),
.B2(n_1559),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1493),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1509),
.B(n_1512),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_SL g1624 ( 
.A1(n_1518),
.A2(n_1537),
.B1(n_1505),
.B2(n_1557),
.Y(n_1624)
);

INVx4_ASAP7_75t_L g1625 ( 
.A(n_1552),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1512),
.B(n_1486),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1524),
.B(n_1570),
.Y(n_1627)
);

AO21x1_ASAP7_75t_L g1628 ( 
.A1(n_1574),
.A2(n_1549),
.B(n_1547),
.Y(n_1628)
);

OAI21xp33_ASAP7_75t_SL g1629 ( 
.A1(n_1507),
.A2(n_1526),
.B(n_1488),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1486),
.B(n_1488),
.Y(n_1630)
);

OAI221xp5_ASAP7_75t_L g1631 ( 
.A1(n_1559),
.A2(n_1568),
.B1(n_1569),
.B2(n_1534),
.C(n_1532),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1531),
.B(n_1564),
.Y(n_1632)
);

OAI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1568),
.A2(n_1569),
.B1(n_1534),
.B2(n_1532),
.C(n_1547),
.Y(n_1633)
);

NOR2xp67_ASAP7_75t_SL g1634 ( 
.A(n_1552),
.B(n_1575),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1502),
.B(n_1505),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1613),
.B(n_1538),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1615),
.B(n_1538),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1593),
.B(n_1505),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1615),
.B(n_1538),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_SL g1640 ( 
.A(n_1601),
.B(n_1537),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1635),
.B(n_1538),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1593),
.B(n_1505),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1587),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1635),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1629),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1614),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1624),
.B(n_1521),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1611),
.B(n_1521),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1605),
.B(n_1549),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1617),
.Y(n_1650)
);

INVxp67_ASAP7_75t_SL g1651 ( 
.A(n_1628),
.Y(n_1651)
);

NAND2x1p5_ASAP7_75t_L g1652 ( 
.A(n_1634),
.B(n_1537),
.Y(n_1652)
);

BUFx2_ASAP7_75t_L g1653 ( 
.A(n_1587),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1588),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1578),
.A2(n_1518),
.B1(n_1486),
.B2(n_1507),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1600),
.A2(n_1575),
.B1(n_1530),
.B2(n_1545),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_1592),
.Y(n_1657)
);

OAI222xp33_ASAP7_75t_L g1658 ( 
.A1(n_1604),
.A2(n_1488),
.B1(n_1574),
.B2(n_1533),
.C1(n_1548),
.C2(n_1544),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1632),
.Y(n_1659)
);

BUFx6f_ASAP7_75t_L g1660 ( 
.A(n_1625),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1595),
.A2(n_1533),
.B1(n_1558),
.B2(n_1548),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1602),
.B(n_1495),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1608),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1602),
.B(n_1494),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1607),
.B(n_1494),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1603),
.B(n_1484),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1644),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1654),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1650),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1646),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1648),
.B(n_1609),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1646),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1644),
.B(n_1606),
.Y(n_1673)
);

AND2x4_ASAP7_75t_SL g1674 ( 
.A(n_1660),
.B(n_1576),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1646),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1640),
.A2(n_1598),
.B1(n_1576),
.B2(n_1619),
.Y(n_1676)
);

NOR2xp67_ASAP7_75t_L g1677 ( 
.A(n_1643),
.B(n_1633),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1650),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1642),
.Y(n_1679)
);

OAI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1655),
.A2(n_1591),
.B1(n_1583),
.B2(n_1610),
.C(n_1584),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1648),
.B(n_1580),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1649),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1640),
.A2(n_1619),
.B1(n_1620),
.B2(n_1576),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1648),
.B(n_1589),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1649),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1643),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1663),
.B(n_1630),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1655),
.A2(n_1591),
.B1(n_1584),
.B2(n_1631),
.Y(n_1688)
);

OAI31xp33_ASAP7_75t_L g1689 ( 
.A1(n_1656),
.A2(n_1620),
.A3(n_1636),
.B(n_1661),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1653),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1649),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1642),
.B(n_1599),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1659),
.B(n_1626),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1643),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1643),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1659),
.B(n_1626),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1641),
.B(n_1590),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1638),
.B(n_1590),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1641),
.B(n_1621),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1654),
.B(n_1627),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1672),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1690),
.B(n_1645),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1682),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1680),
.A2(n_1689),
.B1(n_1688),
.B2(n_1676),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1672),
.Y(n_1705)
);

AND2x4_ASAP7_75t_SL g1706 ( 
.A(n_1683),
.B(n_1660),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1686),
.B(n_1643),
.Y(n_1707)
);

NAND2x1p5_ASAP7_75t_L g1708 ( 
.A(n_1690),
.B(n_1653),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1675),
.Y(n_1709)
);

NAND3xp33_ASAP7_75t_L g1710 ( 
.A(n_1689),
.B(n_1651),
.C(n_1666),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1679),
.B(n_1645),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1686),
.B(n_1653),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1681),
.B(n_1645),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1697),
.B(n_1651),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1670),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1697),
.B(n_1637),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1670),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1681),
.B(n_1636),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1686),
.B(n_1636),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1694),
.B(n_1641),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1670),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1667),
.B(n_1637),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1694),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1694),
.B(n_1647),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1695),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1695),
.Y(n_1726)
);

INVx4_ASAP7_75t_L g1727 ( 
.A(n_1674),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1678),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1695),
.B(n_1647),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1693),
.B(n_1647),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1693),
.B(n_1637),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1699),
.B(n_1639),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1669),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1696),
.B(n_1639),
.Y(n_1734)
);

INVx2_ASAP7_75t_SL g1735 ( 
.A(n_1669),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1685),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1736),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1711),
.B(n_1671),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1736),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1714),
.B(n_1699),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1703),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1711),
.B(n_1671),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1713),
.B(n_1684),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1703),
.Y(n_1744)
);

NOR2x1p5_ASAP7_75t_L g1745 ( 
.A(n_1727),
.B(n_1668),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1701),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1713),
.B(n_1684),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1714),
.B(n_1673),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1713),
.B(n_1687),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1702),
.B(n_1687),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1701),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1708),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1701),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1705),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1702),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1702),
.Y(n_1756)
);

NAND2x1p5_ASAP7_75t_L g1757 ( 
.A(n_1727),
.B(n_1677),
.Y(n_1757)
);

NAND3xp33_ASAP7_75t_SL g1758 ( 
.A(n_1704),
.B(n_1683),
.C(n_1700),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1727),
.B(n_1677),
.Y(n_1759)
);

OAI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1710),
.A2(n_1666),
.B1(n_1652),
.B2(n_1656),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1704),
.A2(n_1524),
.B(n_1665),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1705),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1710),
.B(n_1692),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1708),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1705),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_SL g1766 ( 
.A(n_1727),
.B(n_1658),
.Y(n_1766)
);

AOI32xp33_ASAP7_75t_L g1767 ( 
.A1(n_1706),
.A2(n_1665),
.A3(n_1674),
.B1(n_1662),
.B2(n_1664),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1714),
.B(n_1673),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1732),
.B(n_1691),
.Y(n_1769)
);

XNOR2x1_ASAP7_75t_L g1770 ( 
.A(n_1730),
.B(n_1581),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1730),
.B(n_1687),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1708),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1708),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1706),
.A2(n_1674),
.B1(n_1687),
.B2(n_1623),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1732),
.B(n_1698),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1709),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1709),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1706),
.B(n_1665),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1706),
.B(n_1662),
.Y(n_1779)
);

INVxp67_ASAP7_75t_SL g1780 ( 
.A(n_1770),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1746),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1745),
.B(n_1727),
.Y(n_1782)
);

INVx1_ASAP7_75t_SL g1783 ( 
.A(n_1770),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1769),
.Y(n_1784)
);

NAND2x1_ASAP7_75t_L g1785 ( 
.A(n_1759),
.B(n_1735),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1759),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1763),
.B(n_1730),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1758),
.B(n_1718),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1751),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1750),
.B(n_1718),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1761),
.B(n_1616),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1753),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1760),
.B(n_1718),
.Y(n_1793)
);

INVxp67_ASAP7_75t_SL g1794 ( 
.A(n_1757),
.Y(n_1794)
);

AND4x1_ASAP7_75t_L g1795 ( 
.A(n_1766),
.B(n_1618),
.C(n_1661),
.D(n_1577),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1754),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1750),
.B(n_1731),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1739),
.B(n_1731),
.Y(n_1798)
);

INVxp67_ASAP7_75t_SL g1799 ( 
.A(n_1757),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1738),
.B(n_1731),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1742),
.B(n_1734),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1769),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1749),
.B(n_1759),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1762),
.Y(n_1804)
);

NOR2x1_ASAP7_75t_L g1805 ( 
.A(n_1737),
.B(n_1712),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1755),
.Y(n_1806)
);

AOI32xp33_ASAP7_75t_L g1807 ( 
.A1(n_1778),
.A2(n_1596),
.A3(n_1724),
.B1(n_1729),
.B2(n_1719),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1756),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1749),
.B(n_1734),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1765),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1776),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1777),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1737),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1740),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1774),
.B(n_1585),
.Y(n_1815)
);

OAI21xp33_ASAP7_75t_L g1816 ( 
.A1(n_1780),
.A2(n_1788),
.B(n_1783),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1785),
.Y(n_1817)
);

O2A1O1Ixp33_ASAP7_75t_SL g1818 ( 
.A1(n_1785),
.A2(n_1773),
.B(n_1779),
.C(n_1740),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1806),
.Y(n_1819)
);

AOI221xp5_ASAP7_75t_SL g1820 ( 
.A1(n_1793),
.A2(n_1744),
.B1(n_1741),
.B2(n_1764),
.C(n_1772),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1808),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1808),
.Y(n_1822)
);

INVxp67_ASAP7_75t_SL g1823 ( 
.A(n_1808),
.Y(n_1823)
);

AOI222xp33_ASAP7_75t_L g1824 ( 
.A1(n_1787),
.A2(n_1664),
.B1(n_1662),
.B2(n_1719),
.C1(n_1729),
.C2(n_1724),
.Y(n_1824)
);

OAI321xp33_ASAP7_75t_L g1825 ( 
.A1(n_1807),
.A2(n_1767),
.A3(n_1757),
.B1(n_1708),
.B2(n_1764),
.C(n_1772),
.Y(n_1825)
);

OAI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1795),
.A2(n_1775),
.B1(n_1748),
.B2(n_1768),
.Y(n_1826)
);

AOI221x1_ASAP7_75t_L g1827 ( 
.A1(n_1813),
.A2(n_1752),
.B1(n_1712),
.B2(n_1733),
.C(n_1747),
.Y(n_1827)
);

AOI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1782),
.A2(n_1743),
.B1(n_1747),
.B2(n_1771),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1786),
.B(n_1743),
.Y(n_1829)
);

NAND4xp25_ASAP7_75t_L g1830 ( 
.A(n_1807),
.B(n_1612),
.C(n_1752),
.D(n_1586),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1781),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1786),
.B(n_1775),
.Y(n_1832)
);

INVx2_ASAP7_75t_SL g1833 ( 
.A(n_1803),
.Y(n_1833)
);

AOI31xp33_ASAP7_75t_L g1834 ( 
.A1(n_1782),
.A2(n_1582),
.A3(n_1768),
.B(n_1748),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1781),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1789),
.Y(n_1836)
);

AOI21xp33_ASAP7_75t_L g1837 ( 
.A1(n_1794),
.A2(n_1712),
.B(n_1719),
.Y(n_1837)
);

OAI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1795),
.A2(n_1652),
.B1(n_1732),
.B2(n_1657),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1803),
.B(n_1790),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1789),
.Y(n_1840)
);

NAND3xp33_ASAP7_75t_SL g1841 ( 
.A(n_1814),
.B(n_1597),
.C(n_1622),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_SL g1842 ( 
.A1(n_1826),
.A2(n_1799),
.B1(n_1815),
.B2(n_1791),
.Y(n_1842)
);

AOI21xp5_ASAP7_75t_SL g1843 ( 
.A1(n_1826),
.A2(n_1813),
.B(n_1802),
.Y(n_1843)
);

OAI21xp33_ASAP7_75t_L g1844 ( 
.A1(n_1816),
.A2(n_1798),
.B(n_1784),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1823),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1819),
.B(n_1784),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1838),
.A2(n_1805),
.B(n_1802),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1823),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1821),
.Y(n_1849)
);

INVxp67_ASAP7_75t_L g1850 ( 
.A(n_1841),
.Y(n_1850)
);

INVxp67_ASAP7_75t_L g1851 ( 
.A(n_1841),
.Y(n_1851)
);

INVx2_ASAP7_75t_SL g1852 ( 
.A(n_1839),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1822),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1831),
.Y(n_1854)
);

AOI31xp33_ASAP7_75t_L g1855 ( 
.A1(n_1838),
.A2(n_1805),
.A3(n_1784),
.B(n_1802),
.Y(n_1855)
);

AND2x2_ASAP7_75t_SL g1856 ( 
.A(n_1832),
.B(n_1790),
.Y(n_1856)
);

INVx2_ASAP7_75t_SL g1857 ( 
.A(n_1817),
.Y(n_1857)
);

OAI322xp33_ASAP7_75t_L g1858 ( 
.A1(n_1829),
.A2(n_1792),
.A3(n_1811),
.B1(n_1810),
.B2(n_1796),
.C1(n_1804),
.C2(n_1812),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1834),
.A2(n_1800),
.B1(n_1801),
.B2(n_1797),
.Y(n_1859)
);

INVxp67_ASAP7_75t_L g1860 ( 
.A(n_1833),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1820),
.B(n_1797),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1835),
.Y(n_1862)
);

OAI21xp5_ASAP7_75t_SL g1863 ( 
.A1(n_1842),
.A2(n_1830),
.B(n_1828),
.Y(n_1863)
);

OAI21xp5_ASAP7_75t_SL g1864 ( 
.A1(n_1850),
.A2(n_1827),
.B(n_1837),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1845),
.Y(n_1865)
);

OAI22xp5_ASAP7_75t_L g1866 ( 
.A1(n_1843),
.A2(n_1809),
.B1(n_1836),
.B2(n_1840),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1851),
.A2(n_1809),
.B1(n_1771),
.B2(n_1825),
.Y(n_1867)
);

OAI211xp5_ASAP7_75t_L g1868 ( 
.A1(n_1847),
.A2(n_1818),
.B(n_1824),
.C(n_1812),
.Y(n_1868)
);

INVx1_ASAP7_75t_SL g1869 ( 
.A(n_1856),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1848),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1852),
.B(n_1792),
.Y(n_1871)
);

XNOR2x1_ASAP7_75t_L g1872 ( 
.A(n_1859),
.B(n_1594),
.Y(n_1872)
);

OA21x2_ASAP7_75t_L g1873 ( 
.A1(n_1855),
.A2(n_1810),
.B(n_1804),
.Y(n_1873)
);

INVxp67_ASAP7_75t_L g1874 ( 
.A(n_1857),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1865),
.Y(n_1875)
);

INVx1_ASAP7_75t_SL g1876 ( 
.A(n_1869),
.Y(n_1876)
);

INVx1_ASAP7_75t_SL g1877 ( 
.A(n_1873),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1874),
.B(n_1860),
.Y(n_1878)
);

AOI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1866),
.A2(n_1855),
.B1(n_1844),
.B2(n_1859),
.C(n_1858),
.Y(n_1879)
);

NAND3xp33_ASAP7_75t_L g1880 ( 
.A(n_1873),
.B(n_1846),
.C(n_1849),
.Y(n_1880)
);

AOI211x1_ASAP7_75t_SL g1881 ( 
.A1(n_1867),
.A2(n_1861),
.B(n_1853),
.C(n_1854),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1863),
.B(n_1862),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1870),
.B(n_1796),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1871),
.Y(n_1884)
);

AOI222xp33_ASAP7_75t_L g1885 ( 
.A1(n_1879),
.A2(n_1864),
.B1(n_1868),
.B2(n_1811),
.C1(n_1872),
.C2(n_1712),
.Y(n_1885)
);

AOI221x1_ASAP7_75t_L g1886 ( 
.A1(n_1880),
.A2(n_1878),
.B1(n_1875),
.B2(n_1882),
.C(n_1884),
.Y(n_1886)
);

NAND3xp33_ASAP7_75t_SL g1887 ( 
.A(n_1881),
.B(n_1877),
.C(n_1876),
.Y(n_1887)
);

AOI211x1_ASAP7_75t_L g1888 ( 
.A1(n_1883),
.A2(n_1724),
.B(n_1729),
.C(n_1722),
.Y(n_1888)
);

AOI211x1_ASAP7_75t_SL g1889 ( 
.A1(n_1880),
.A2(n_1733),
.B(n_1726),
.C(n_1723),
.Y(n_1889)
);

OAI221xp5_ASAP7_75t_L g1890 ( 
.A1(n_1879),
.A2(n_1722),
.B1(n_1735),
.B2(n_1652),
.C(n_1716),
.Y(n_1890)
);

OAI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1887),
.A2(n_1712),
.B(n_1707),
.Y(n_1891)
);

INVxp33_ASAP7_75t_L g1892 ( 
.A(n_1886),
.Y(n_1892)
);

A2O1A1Ixp33_ASAP7_75t_L g1893 ( 
.A1(n_1890),
.A2(n_1712),
.B(n_1735),
.C(n_1707),
.Y(n_1893)
);

AO22x2_ASAP7_75t_L g1894 ( 
.A1(n_1885),
.A2(n_1733),
.B1(n_1707),
.B2(n_1726),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1889),
.A2(n_1707),
.B(n_1723),
.Y(n_1895)
);

NOR3xp33_ASAP7_75t_L g1896 ( 
.A(n_1888),
.B(n_1573),
.C(n_1579),
.Y(n_1896)
);

NAND4xp75_ASAP7_75t_L g1897 ( 
.A(n_1891),
.B(n_1892),
.C(n_1895),
.D(n_1894),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1896),
.Y(n_1898)
);

AOI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1893),
.A2(n_1707),
.B1(n_1720),
.B2(n_1726),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1894),
.Y(n_1900)
);

NAND2x1_ASAP7_75t_SL g1901 ( 
.A(n_1894),
.B(n_1733),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_SL g1902 ( 
.A1(n_1898),
.A2(n_1554),
.B1(n_1498),
.B2(n_1493),
.Y(n_1902)
);

NAND3xp33_ASAP7_75t_SL g1903 ( 
.A(n_1900),
.B(n_1554),
.C(n_1652),
.Y(n_1903)
);

AOI221xp5_ASAP7_75t_L g1904 ( 
.A1(n_1899),
.A2(n_1707),
.B1(n_1723),
.B2(n_1726),
.C(n_1725),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1902),
.A2(n_1897),
.B(n_1901),
.Y(n_1905)
);

OAI22x1_ASAP7_75t_L g1906 ( 
.A1(n_1905),
.A2(n_1903),
.B1(n_1725),
.B2(n_1723),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1906),
.Y(n_1907)
);

INVxp67_ASAP7_75t_L g1908 ( 
.A(n_1906),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1907),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_SL g1910 ( 
.A1(n_1908),
.A2(n_1904),
.B1(n_1725),
.B2(n_1715),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1909),
.A2(n_1725),
.B(n_1721),
.Y(n_1911)
);

OAI21x1_ASAP7_75t_SL g1912 ( 
.A1(n_1910),
.A2(n_1717),
.B(n_1715),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1911),
.A2(n_1721),
.B(n_1715),
.Y(n_1913)
);

NOR2xp67_ASAP7_75t_SL g1914 ( 
.A(n_1913),
.B(n_1912),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1914),
.Y(n_1915)
);

AOI221xp5_ASAP7_75t_L g1916 ( 
.A1(n_1915),
.A2(n_1717),
.B1(n_1715),
.B2(n_1721),
.C(n_1728),
.Y(n_1916)
);

AOI211xp5_ASAP7_75t_L g1917 ( 
.A1(n_1916),
.A2(n_1572),
.B(n_1526),
.C(n_1573),
.Y(n_1917)
);


endmodule