module real_jpeg_5090_n_6 (n_46, n_5, n_4, n_0, n_1, n_47, n_2, n_48, n_50, n_3, n_49, n_6);

input n_46;
input n_5;
input n_4;
input n_0;
input n_1;
input n_47;
input n_2;
input n_48;
input n_50;
input n_3;
input n_49;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_40;
wire n_39;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_32),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_1),
.B(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_2),
.B(n_11),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_5),
.B(n_36),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_7),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_17),
.B1(n_43),
.B2(n_44),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_9),
.B(n_15),
.Y(n_8)
);

INVxp67_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_23),
.B(n_42),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_22),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_22),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_21),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_35),
.B(n_41),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_34),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_33),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_46),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_47),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_48),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_49),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_50),
.Y(n_40)
);


endmodule