module real_jpeg_26382_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_0),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_0),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_0),
.B(n_48),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_0),
.B(n_51),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_0),
.B(n_28),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_0),
.B(n_17),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_0),
.B(n_56),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_0),
.B(n_68),
.Y(n_211)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_3),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_3),
.B(n_43),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_3),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_3),
.B(n_65),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_3),
.B(n_68),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_3),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_3),
.B(n_28),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_3),
.B(n_56),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_5),
.B(n_28),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_5),
.B(n_56),
.Y(n_97)
);

INVx8_ASAP7_75t_SL g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_8),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_9),
.B(n_68),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_9),
.B(n_28),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_9),
.B(n_51),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_9),
.B(n_43),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_9),
.B(n_48),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_11),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_11),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_11),
.B(n_68),
.Y(n_96)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_13),
.B(n_56),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_13),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_13),
.B(n_43),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_13),
.B(n_28),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_13),
.B(n_17),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_14),
.B(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_14),
.B(n_68),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_14),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_14),
.B(n_51),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_14),
.B(n_56),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_14),
.B(n_40),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_14),
.B(n_28),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_15),
.B(n_28),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_15),
.B(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_15),
.B(n_51),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_15),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_15),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_16),
.B(n_56),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_16),
.B(n_28),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_16),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_16),
.B(n_68),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_16),
.B(n_51),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_16),
.B(n_43),
.Y(n_234)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_17),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_155),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_130),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_53),
.C(n_60),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_22),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.C(n_46),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_23),
.B(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_33),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_30),
.C(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_27),
.B(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_32),
.Y(n_185)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_38),
.A2(n_39),
.B(n_42),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_38),
.B(n_46),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_41),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.C(n_52),
.Y(n_46)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_47),
.B(n_50),
.CI(n_52),
.CON(n_134),
.SN(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_48),
.Y(n_80)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_53),
.B(n_60),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_55),
.B(n_58),
.C(n_59),
.Y(n_119)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_57),
.B(n_63),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_70),
.C(n_72),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_61),
.B(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.C(n_67),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_62),
.B(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_66),
.B(n_67),
.Y(n_251)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_98),
.B2(n_129),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_88),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_82),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_83),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_84),
.A2(n_86),
.B1(n_90),
.B2(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_90),
.C(n_91),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_92),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx24_ASAP7_75t_SL g269 ( 
.A(n_94),
.Y(n_269)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.CI(n_97),
.CON(n_94),
.SN(n_94)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_98),
.Y(n_273)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_119),
.CI(n_120),
.CON(n_98),
.SN(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.C(n_115),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_100),
.B(n_152),
.Y(n_151)
);

BUFx24_ASAP7_75t_SL g271 ( 
.A(n_100),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_104),
.CI(n_107),
.CON(n_100),
.SN(n_100)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_104),
.C(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_105),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_109),
.B(n_115),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.C(n_113),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_128),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_124),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_151),
.C(n_153),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_131),
.A2(n_132),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_147),
.C(n_149),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_133),
.B(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.C(n_143),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_134),
.B(n_244),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g268 ( 
.A(n_134),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_135),
.A2(n_136),
.B1(n_143),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_143),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.C(n_146),
.Y(n_143)
);

FAx1_ASAP7_75t_SL g230 ( 
.A(n_144),
.B(n_145),
.CI(n_146),
.CON(n_230),
.SN(n_230)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_147),
.B(n_149),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_151),
.B(n_153),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_264),
.C(n_265),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_254),
.C(n_255),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_237),
.C(n_238),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_224),
.C(n_225),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_206),
.C(n_207),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_186),
.C(n_187),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_174),
.C(n_179),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_170),
.B2(n_171),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_172),
.C(n_173),
.Y(n_186)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_165),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_169),
.Y(n_190)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.C(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_197),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_192),
.C(n_197),
.Y(n_206)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_193),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_194),
.B(n_196),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_205),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_198),
.Y(n_205)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_201),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_204),
.C(n_205),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_215),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_210),
.C(n_215),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_213),
.C(n_214),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_218),
.C(n_219),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_223),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_231),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_232),
.C(n_236),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_229),
.C(n_230),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_230),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_232),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_234),
.CI(n_235),
.CON(n_232),
.SN(n_232)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_246),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_242),
.C(n_246),
.Y(n_254)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_250),
.C(n_252),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_249),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_250),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_263),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_260),
.C(n_261),
.Y(n_264)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_259),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_266),
.Y(n_267)
);


endmodule