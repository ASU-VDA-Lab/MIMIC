module real_jpeg_4409_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_1),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_1),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_1),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_1),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_1),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_1),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_1),
.B(n_223),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_1),
.B(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_2),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_2),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_2),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_2),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_2),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_2),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_2),
.B(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_3),
.Y(n_123)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_4),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_4),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_4),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_4),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_4),
.B(n_272),
.Y(n_271)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_6),
.Y(n_125)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_6),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_6),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_7),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_7),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_8),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_8),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_8),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_8),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_8),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_8),
.B(n_197),
.Y(n_196)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_10),
.Y(n_96)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_10),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g195 ( 
.A(n_10),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_11),
.B(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_11),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_11),
.B(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_11),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_12),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_12),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_12),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_12),
.B(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_13),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_14),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_14),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_14),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_14),
.B(n_327),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_15),
.B(n_26),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_15),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_15),
.B(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_205),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_204),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_161),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_19),
.B(n_161),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.C(n_131),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_20),
.A2(n_21),
.B1(n_104),
.B2(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_66),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_22),
.B(n_67),
.C(n_84),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.C(n_54),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_23),
.B(n_54),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_25),
.B(n_30),
.C(n_34),
.Y(n_106)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_29),
.Y(n_143)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_29),
.Y(n_173)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_33),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_38),
.Y(n_197)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_39),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_40),
.B(n_367),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_46),
.C(n_50),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_41),
.B(n_50),
.Y(n_134)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_44),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_45),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_46),
.B(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_49),
.Y(n_333)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.C(n_61),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_55),
.A2(n_166),
.B1(n_167),
.B2(n_174),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_55),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_55),
.A2(n_61),
.B1(n_166),
.B2(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_59),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_60),
.A2(n_346),
.B1(n_347),
.B2(n_349),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_60),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_61),
.Y(n_348)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_64),
.Y(n_130)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_84),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_76),
.C(n_79),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_68),
.B(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_68),
.A2(n_69),
.B(n_71),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_75),
.B(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_76),
.B(n_79),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_80),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_80),
.B(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_80),
.B(n_280),
.Y(n_279)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_97),
.Y(n_84)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_85),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.C(n_95),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_86),
.A2(n_95),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_86),
.A2(n_158),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_90),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

OR2x2_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_91),
.Y(n_230)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_93),
.Y(n_169)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_93),
.Y(n_239)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_110),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_125),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_95),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_98),
.B(n_101),
.C(n_191),
.Y(n_190)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_104),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_117),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_106),
.B(n_107),
.C(n_117),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_116),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_109),
.B(n_201),
.C(n_202),
.Y(n_200)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_114),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_127),
.B2(n_128),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_124),
.B2(n_126),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_120),
.A2(n_121),
.B1(n_136),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_136),
.C(n_139),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_124),
.C(n_128),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_122),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

BUFx8_ASAP7_75t_L g290 ( 
.A(n_123),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_124),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_124),
.A2(n_126),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_124),
.A2(n_126),
.B1(n_236),
.B2(n_237),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_126),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_130),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_131),
.B(n_372),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_153),
.C(n_159),
.Y(n_131)
);

FAx1_ASAP7_75t_L g363 ( 
.A(n_132),
.B(n_153),
.CI(n_159),
.CON(n_363),
.SN(n_363)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.C(n_144),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_133),
.B(n_355),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_135),
.A2(n_144),
.B1(n_145),
.B2(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_135),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_136),
.Y(n_312)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_139),
.B(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_315)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_149),
.Y(n_282)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_158),
.B(n_246),
.Y(n_322)
);

BUFx24_ASAP7_75t_SL g379 ( 
.A(n_161),
.Y(n_379)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_187),
.CI(n_203),
.CON(n_161),
.SN(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_177),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_175),
.B2(n_176),
.Y(n_163)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_173),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_186),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_182),
.A2(n_183),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_183),
.B(n_228),
.C(n_233),
.Y(n_314)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_200),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_193)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_194),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_196),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_359),
.B(n_374),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_337),
.B(n_358),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_305),
.B(n_336),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_260),
.B(n_304),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_251),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_211),
.B(n_251),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_234),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_225),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_213),
.B(n_225),
.C(n_234),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.C(n_221),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_221),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_233),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_240),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_235),
.B(n_319),
.C(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_245),
.Y(n_240)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_241),
.Y(n_319)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_245),
.Y(n_320)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.C(n_259),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_252),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_254),
.A2(n_259),
.B1(n_296),
.B2(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_255),
.Y(n_294)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_257),
.Y(n_295)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_259),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_298),
.B(n_303),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_284),
.B(n_297),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_269),
.B(n_283),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_279),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_279),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_274),
.B(n_278),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_274),
.Y(n_278)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_286),
.B1(n_291),
.B2(n_292),
.Y(n_285)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx8_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_293),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_293),
.Y(n_297)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_286),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_287),
.A2(n_288),
.B(n_291),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_295),
.B(n_296),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_307),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_316),
.B2(n_317),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_308),
.B(n_318),
.C(n_321),
.Y(n_338)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_313),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_310),
.B(n_314),
.C(n_315),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_321),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_324),
.B2(n_335),
.Y(n_321)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_322),
.Y(n_335)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_330),
.B2(n_334),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_334),
.C(n_335),
.Y(n_342)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_338),
.B(n_339),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_341),
.B1(n_352),
.B2(n_357),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_340),
.B(n_353),
.C(n_354),
.Y(n_368)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_345),
.C(n_350),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_350),
.B2(n_351),
.Y(n_343)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_344),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_345),
.Y(n_351)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_347),
.Y(n_349)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_352),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_369),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_368),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_368),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_365),
.C(n_366),
.Y(n_370)
);

BUFx24_ASAP7_75t_SL g378 ( 
.A(n_363),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_369),
.A2(n_376),
.B(n_377),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_370),
.B(n_371),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);


endmodule