module fake_jpeg_13956_n_304 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_304);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_265;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_21),
.B(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_51),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_63),
.Y(n_73)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_47),
.B(n_65),
.Y(n_91)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_48),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_59),
.Y(n_92)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_29),
.B(n_1),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_22),
.B(n_1),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_16),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_29),
.B1(n_19),
.B2(n_43),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_70),
.A2(n_72),
.B1(n_82),
.B2(n_86),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_43),
.B1(n_19),
.B2(n_34),
.Y(n_72)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_32),
.B1(n_24),
.B2(n_40),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_78),
.A2(n_100),
.B1(n_101),
.B2(n_112),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_79),
.B(n_81),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_28),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_55),
.A2(n_43),
.B1(n_19),
.B2(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_85),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_34),
.B1(n_41),
.B2(n_20),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_41),
.B1(n_39),
.B2(n_35),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_33),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_35),
.B1(n_40),
.B2(n_39),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_95),
.B1(n_48),
.B2(n_61),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_42),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_94),
.B(n_102),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_32),
.B1(n_24),
.B2(n_22),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_41),
.B1(n_38),
.B2(n_25),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_51),
.A2(n_41),
.B1(n_38),
.B2(n_25),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_42),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_50),
.B(n_31),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_108),
.B(n_111),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_68),
.A2(n_41),
.B1(n_23),
.B2(n_33),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_66),
.B(n_23),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_61),
.A2(n_33),
.B1(n_3),
.B2(n_4),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_2),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_49),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_114),
.B(n_121),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_115),
.B(n_117),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_125),
.Y(n_151)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_52),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g167 ( 
.A(n_120),
.B(n_10),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_67),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_3),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_123),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_71),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_67),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_127),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_61),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_143),
.B1(n_89),
.B2(n_88),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_48),
.B(n_5),
.C(n_6),
.Y(n_130)
);

OR2x6_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_133),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_74),
.B(n_12),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_131),
.B(n_142),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_69),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_4),
.Y(n_133)
);

BUFx8_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_74),
.B(n_11),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_76),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_85),
.B1(n_77),
.B2(n_84),
.Y(n_154)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_147),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_69),
.B(n_8),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_75),
.B(n_8),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_149),
.B(n_133),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_98),
.B(n_11),
.C(n_10),
.Y(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g199 ( 
.A1(n_150),
.A2(n_161),
.B(n_174),
.C(n_176),
.D(n_169),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_177),
.Y(n_198)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_164),
.B1(n_166),
.B2(n_127),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_141),
.A2(n_104),
.B1(n_99),
.B2(n_107),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_158),
.Y(n_185)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_141),
.A2(n_104),
.B1(n_107),
.B2(n_97),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_172),
.Y(n_200)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_125),
.A2(n_98),
.A3(n_88),
.B1(n_89),
.B2(n_75),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_162),
.B(n_171),
.Y(n_197)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_106),
.B1(n_96),
.B2(n_97),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_146),
.A2(n_109),
.B1(n_96),
.B2(n_10),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_167),
.A2(n_173),
.B(n_168),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_120),
.A2(n_135),
.B1(n_146),
.B2(n_119),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_115),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_116),
.B(n_124),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_175),
.B(n_178),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_114),
.B(n_133),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_121),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

AO22x2_ASAP7_75t_L g184 ( 
.A1(n_173),
.A2(n_130),
.B1(n_119),
.B2(n_120),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_187),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_151),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_129),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_203),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_152),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_192),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_138),
.B1(n_134),
.B2(n_145),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_172),
.B1(n_177),
.B2(n_159),
.Y(n_220)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_121),
.B(n_148),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_207),
.B(n_173),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_199),
.A2(n_179),
.B(n_169),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_160),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_201),
.Y(n_231)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_148),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_181),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_209),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_210),
.B(n_165),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_128),
.C(n_136),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_128),
.C(n_156),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_170),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_173),
.A2(n_138),
.B(n_144),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_203),
.B(n_171),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_216),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_222),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_150),
.B(n_167),
.Y(n_223)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_223),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_199),
.A2(n_168),
.B(n_174),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_227),
.C(n_228),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_200),
.A2(n_155),
.B(n_178),
.Y(n_228)
);

HAxp5_ASAP7_75t_SL g247 ( 
.A(n_229),
.B(n_184),
.CON(n_247),
.SN(n_247)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_200),
.A2(n_165),
.B1(n_170),
.B2(n_118),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_185),
.B1(n_193),
.B2(n_189),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_210),
.A2(n_188),
.B(n_198),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_184),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_220),
.A2(n_197),
.B1(n_232),
.B2(n_185),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_233),
.A2(n_225),
.B1(n_227),
.B2(n_217),
.Y(n_254)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_236),
.A2(n_239),
.B1(n_245),
.B2(n_246),
.Y(n_252)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_241),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_184),
.B1(n_183),
.B2(n_208),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_240),
.B(n_243),
.Y(n_256)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_221),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_218),
.B1(n_224),
.B2(n_223),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_229),
.A2(n_228),
.B1(n_230),
.B2(n_222),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_247),
.A2(n_225),
.B(n_226),
.Y(n_253)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_248),
.B(n_189),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_211),
.C(n_216),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_212),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_242),
.B(n_124),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_234),
.Y(n_266)
);

AO21x1_ASAP7_75t_L g274 ( 
.A1(n_253),
.A2(n_254),
.B(n_247),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_261),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_263),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_221),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_263),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_239),
.A2(n_212),
.B1(n_202),
.B2(n_170),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_243),
.B1(n_241),
.B2(n_250),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_190),
.B1(n_195),
.B2(n_194),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_264),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_266),
.B(n_271),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_267),
.A2(n_269),
.B1(n_273),
.B2(n_236),
.Y(n_284)
);

BUFx24_ASAP7_75t_SL g268 ( 
.A(n_258),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_191),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_250),
.B1(n_237),
.B2(n_242),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_191),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_274),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_258),
.A2(n_250),
.B1(n_244),
.B2(n_234),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_270),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_279),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_260),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_280),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_259),
.C(n_254),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_282),
.B(n_134),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_262),
.C(n_253),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_264),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_284),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_277),
.A2(n_265),
.B1(n_257),
.B2(n_190),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_286),
.B(n_287),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_282),
.A2(n_265),
.B1(n_257),
.B2(n_206),
.Y(n_289)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_289),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_276),
.C(n_281),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_292),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_287),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_295),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_294),
.A2(n_288),
.B(n_276),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_147),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_297),
.A2(n_288),
.B(n_280),
.Y(n_299)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_300),
.B(n_296),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_136),
.C(n_140),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_302),
.B(n_140),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_303),
.B(n_140),
.CI(n_245),
.CON(n_304),
.SN(n_304)
);


endmodule