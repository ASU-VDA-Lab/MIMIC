module fake_jpeg_25419_n_310 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

CKINVDCx9p33_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_42),
.Y(n_61)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_45),
.B(n_46),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_49),
.B(n_60),
.Y(n_83)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_25),
.Y(n_53)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_33),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_63),
.Y(n_87)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_42),
.B(n_28),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_16),
.B1(n_23),
.B2(n_18),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_32),
.B1(n_41),
.B2(n_34),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_34),
.B1(n_53),
.B2(n_49),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_68),
.B1(n_78),
.B2(n_80),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_82),
.Y(n_93)
);

CKINVDCx9p33_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_34),
.B1(n_16),
.B2(n_32),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_30),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_44),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_85),
.Y(n_109)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_90),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_86),
.A2(n_26),
.B1(n_19),
.B2(n_25),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_106),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_61),
.B1(n_65),
.B2(n_34),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_105),
.B1(n_110),
.B2(n_114),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_59),
.B1(n_51),
.B2(n_56),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_61),
.B(n_41),
.C(n_54),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_108),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_54),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_63),
.B1(n_52),
.B2(n_50),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_35),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_50),
.B1(n_64),
.B2(n_22),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_71),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_115),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_56),
.B(n_44),
.C(n_58),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_78),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_118),
.A2(n_119),
.B(n_127),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_79),
.B(n_1),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_45),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_120),
.B(n_121),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_95),
.B(n_45),
.Y(n_124)
);

OAI32xp33_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_126),
.A3(n_135),
.B1(n_121),
.B2(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_46),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_46),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_91),
.B(n_20),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_133),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_116),
.B1(n_85),
.B2(n_69),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_43),
.B(n_31),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_139),
.B(n_98),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_11),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_93),
.B(n_20),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_20),
.Y(n_161)
);

NAND2x1_ASAP7_75t_SL g139 ( 
.A(n_97),
.B(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_74),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_35),
.Y(n_142)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_142),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_152),
.Y(n_176)
);

AOI32xp33_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_66),
.A3(n_107),
.B1(n_44),
.B2(n_112),
.Y(n_145)
);

NOR4xp25_ASAP7_75t_SL g171 ( 
.A(n_145),
.B(n_133),
.C(n_132),
.D(n_127),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_148),
.A2(n_151),
.B(n_155),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_141),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_97),
.B(n_113),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_99),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_122),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_153),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_116),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_124),
.Y(n_185)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_159),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_129),
.A2(n_64),
.B1(n_88),
.B2(n_94),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_160),
.A2(n_163),
.B1(n_139),
.B2(n_130),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_162),
.Y(n_180)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_129),
.A2(n_92),
.B1(n_70),
.B2(n_69),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_126),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_122),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_166),
.Y(n_184)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_183),
.B1(n_192),
.B2(n_195),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_154),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_127),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_186),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_193),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_164),
.A2(n_119),
.B1(n_133),
.B2(n_132),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_176),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_160),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_188),
.B(n_148),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_128),
.B1(n_120),
.B2(n_138),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_190),
.A2(n_194),
.B1(n_155),
.B2(n_143),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_146),
.A2(n_136),
.B1(n_92),
.B2(n_103),
.Y(n_192)
);

AO21x1_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_25),
.B(n_125),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_152),
.A2(n_103),
.B1(n_70),
.B2(n_82),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_146),
.A2(n_75),
.B1(n_125),
.B2(n_37),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_199),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_211),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_192),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_210),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_212),
.B1(n_215),
.B2(n_216),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_177),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_208),
.Y(n_231)
);

AO22x1_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_144),
.B1(n_165),
.B2(n_143),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_209),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_167),
.C(n_157),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_163),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_183),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_213),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_170),
.A2(n_188),
.B1(n_174),
.B2(n_175),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_214),
.A2(n_37),
.B1(n_31),
.B2(n_24),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_194),
.A2(n_168),
.B1(n_158),
.B2(n_149),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_219),
.B1(n_125),
.B2(n_98),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_33),
.C(n_71),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_172),
.C(n_182),
.Y(n_221)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_218),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_190),
.C(n_178),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_234),
.C(n_235),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_191),
.C(n_181),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_204),
.C(n_196),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_29),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_236),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_181),
.C(n_71),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_30),
.C(n_21),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_29),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_238),
.A2(n_239),
.B1(n_219),
.B2(n_215),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_37),
.B1(n_31),
.B2(n_24),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_253),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_243),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_202),
.C(n_204),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_223),
.C(n_230),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_224),
.B(n_209),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_29),
.Y(n_265)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_249),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_250),
.Y(n_259)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_251),
.B(n_252),
.Y(n_264)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_201),
.C(n_24),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_201),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_9),
.B(n_15),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_21),
.C(n_9),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_245),
.A2(n_231),
.B1(n_220),
.B2(n_222),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_265),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_244),
.A2(n_222),
.B1(n_226),
.B2(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_30),
.C(n_24),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_241),
.C(n_21),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_246),
.A2(n_242),
.B(n_241),
.C(n_11),
.Y(n_267)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_5),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_277),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_21),
.C(n_27),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_265),
.C(n_264),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_263),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_273),
.B(n_275),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_259),
.A2(n_6),
.B(n_15),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_27),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_6),
.C(n_14),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_12),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_281),
.B(n_13),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_287),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_276),
.A2(n_262),
.B1(n_257),
.B2(n_267),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_0),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_289),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_274),
.A2(n_260),
.B1(n_10),
.B2(n_12),
.Y(n_287)
);

NAND3xp33_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_5),
.C(n_14),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_5),
.B(n_1),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_4),
.B1(n_13),
.B2(n_10),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_291),
.Y(n_298)
);

AOI31xp67_ASAP7_75t_L g292 ( 
.A1(n_288),
.A2(n_279),
.A3(n_271),
.B(n_270),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_294),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_283),
.A2(n_4),
.B(n_13),
.Y(n_294)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_0),
.B(n_1),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_291),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_286),
.C(n_282),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_301),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_302),
.A2(n_298),
.B(n_293),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_304),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_305),
.B(n_303),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_300),
.B(n_301),
.C(n_27),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_0),
.B(n_2),
.Y(n_308)
);

AOI32xp33_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_0),
.A3(n_2),
.B1(n_3),
.B2(n_27),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_3),
.B(n_303),
.Y(n_310)
);


endmodule