module fake_jpeg_1588_n_691 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_691);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_691;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_60),
.Y(n_152)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_30),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_64),
.B(n_129),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_66),
.Y(n_207)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_68),
.Y(n_224)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_30),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g197 ( 
.A(n_69),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_70),
.B(n_131),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_71),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_74),
.Y(n_176)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_76),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_78),
.Y(n_184)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_80),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_81),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_40),
.B(n_8),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_83),
.B(n_27),
.Y(n_136)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_85),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_86),
.Y(n_198)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_88),
.Y(n_229)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_91),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g171 ( 
.A(n_92),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_26),
.A2(n_46),
.B(n_52),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_94),
.A2(n_33),
.B(n_47),
.C(n_49),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_95),
.Y(n_201)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g199 ( 
.A(n_96),
.Y(n_199)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_97),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_98),
.Y(n_172)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_99),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_50),
.Y(n_101)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_101),
.Y(n_203)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_102),
.Y(n_186)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_21),
.Y(n_103)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_103),
.Y(n_196)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_106),
.Y(n_215)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_107),
.Y(n_227)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_21),
.Y(n_109)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_46),
.Y(n_110)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_34),
.Y(n_111)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_21),
.Y(n_112)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_113),
.B(n_125),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_34),
.Y(n_114)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_115),
.Y(n_194)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_21),
.Y(n_116)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_20),
.Y(n_117)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_117),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_118),
.Y(n_216)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_119),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_120),
.Y(n_223)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_121),
.Y(n_226)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_21),
.Y(n_122)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_122),
.Y(n_230)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_21),
.Y(n_123)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_26),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_126),
.Y(n_219)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_127),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_51),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_130),
.Y(n_160)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_51),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g131 ( 
.A(n_24),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_24),
.B(n_8),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_133),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_20),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_136),
.B(n_169),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_83),
.A2(n_27),
.B1(n_45),
.B2(n_44),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g235 ( 
.A1(n_138),
.A2(n_149),
.B1(n_161),
.B2(n_173),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_65),
.A2(n_78),
.B1(n_92),
.B2(n_71),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_140),
.A2(n_180),
.B1(n_63),
.B2(n_1),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_101),
.A2(n_27),
.B1(n_45),
.B2(n_44),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_72),
.A2(n_45),
.B1(n_44),
.B2(n_41),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_154),
.A2(n_175),
.B1(n_183),
.B2(n_193),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_24),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_158),
.B(n_159),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_69),
.B(n_31),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_85),
.A2(n_41),
.B1(n_31),
.B2(n_59),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_82),
.B(n_31),
.Y(n_169)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_95),
.B(n_74),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_170),
.B(n_206),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_103),
.A2(n_41),
.B1(n_59),
.B2(n_28),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_98),
.B(n_20),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_174),
.B(n_178),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_76),
.A2(n_23),
.B1(n_58),
.B2(n_57),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_100),
.B(n_23),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_80),
.A2(n_23),
.B1(n_58),
.B2(n_57),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_105),
.B(n_39),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_182),
.B(n_192),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_81),
.A2(n_59),
.B1(n_58),
.B2(n_57),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_185),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_133),
.B(n_54),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_187),
.B(n_191),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_88),
.B(n_54),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_111),
.B(n_54),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_91),
.A2(n_49),
.B1(n_28),
.B2(n_42),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_114),
.B(n_37),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_205),
.B(n_211),
.Y(n_256)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_118),
.B(n_37),
.Y(n_206)
);

OA22x2_ASAP7_75t_SL g208 ( 
.A1(n_109),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_208)
);

AO22x1_ASAP7_75t_L g276 ( 
.A1(n_208),
.A2(n_139),
.B1(n_196),
.B2(n_173),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_112),
.A2(n_49),
.B1(n_28),
.B2(n_42),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_210),
.A2(n_218),
.B1(n_231),
.B2(n_33),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_120),
.B(n_37),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_124),
.B(n_36),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_212),
.B(n_221),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_116),
.A2(n_36),
.B1(n_42),
.B2(n_39),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_L g221 ( 
.A(n_123),
.B(n_39),
.C(n_38),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_126),
.A2(n_38),
.B1(n_35),
.B2(n_36),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_135),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_232),
.B(n_247),
.Y(n_316)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_233),
.Y(n_321)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_150),
.Y(n_234)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_234),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_236),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_197),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_238),
.B(n_276),
.Y(n_339)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_239),
.Y(n_367)
);

AND2x2_ASAP7_75t_SL g240 ( 
.A(n_162),
.B(n_47),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_240),
.Y(n_332)
);

INVx13_ASAP7_75t_L g241 ( 
.A(n_166),
.Y(n_241)
);

INVx13_ASAP7_75t_L g329 ( 
.A(n_241),
.Y(n_329)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_242),
.Y(n_343)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_166),
.Y(n_243)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_243),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_208),
.A2(n_149),
.B1(n_185),
.B2(n_193),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_244),
.A2(n_314),
.B1(n_201),
.B2(n_220),
.Y(n_374)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_151),
.Y(n_245)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_245),
.Y(n_371)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_166),
.Y(n_246)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_246),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_222),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_177),
.A2(n_32),
.B1(n_35),
.B2(n_38),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_248),
.A2(n_274),
.B(n_292),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_206),
.B(n_47),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_250),
.B(n_265),
.Y(n_320)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_137),
.Y(n_253)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_253),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_255),
.A2(n_263),
.B1(n_273),
.B2(n_290),
.Y(n_337)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_157),
.Y(n_259)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_259),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_177),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_260),
.B(n_280),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_134),
.B(n_130),
.C(n_128),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_261),
.B(n_172),
.C(n_220),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_35),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_262),
.B(n_279),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_213),
.A2(n_32),
.B1(n_33),
.B2(n_122),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_179),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_264),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_160),
.B(n_32),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_266),
.A2(n_304),
.B1(n_312),
.B2(n_168),
.Y(n_348)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_163),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_267),
.Y(n_377)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_145),
.Y(n_268)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_268),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_221),
.A2(n_8),
.B1(n_17),
.B2(n_15),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_269),
.A2(n_278),
.B1(n_309),
.B2(n_229),
.Y(n_330)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_142),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_270),
.Y(n_326)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_146),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_272),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_214),
.A2(n_7),
.B1(n_17),
.B2(n_14),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_161),
.A2(n_7),
.B(n_17),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_145),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_275),
.Y(n_359)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_148),
.Y(n_277)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_277),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_208),
.A2(n_7),
.B1(n_17),
.B2(n_14),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_164),
.B(n_6),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_224),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_194),
.B(n_0),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g368 ( 
.A(n_281),
.B(n_310),
.Y(n_368)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_156),
.Y(n_282)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_146),
.Y(n_283)
);

INVx5_ASAP7_75t_L g328 ( 
.A(n_283),
.Y(n_328)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_139),
.Y(n_284)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_284),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_167),
.B(n_6),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_285),
.B(n_300),
.Y(n_352)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_207),
.Y(n_286)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_219),
.Y(n_287)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_287),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_228),
.Y(n_288)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_288),
.Y(n_342)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_198),
.Y(n_289)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_289),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_217),
.A2(n_5),
.B1(n_14),
.B2(n_13),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_196),
.Y(n_291)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_291),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_141),
.B(n_0),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_293),
.B(n_301),
.Y(n_327)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_228),
.Y(n_294)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_294),
.Y(n_357)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_207),
.Y(n_295)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_295),
.Y(n_362)
);

INVx4_ASAP7_75t_SL g296 ( 
.A(n_186),
.Y(n_296)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_296),
.Y(n_378)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_195),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_297),
.B(n_298),
.Y(n_356)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_163),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_224),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_299),
.B(n_311),
.Y(n_354)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_199),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_143),
.B(n_0),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_153),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_302),
.B(n_305),
.Y(n_375)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_199),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_303),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_231),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_171),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_226),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_306),
.B(n_307),
.Y(n_366)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_195),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_204),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_308),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_210),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_144),
.B(n_170),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_171),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_218),
.A2(n_2),
.B1(n_3),
.B2(n_10),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_165),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_313),
.A2(n_238),
.B1(n_243),
.B2(n_246),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_209),
.B(n_10),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_186),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_315),
.B(n_186),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_258),
.A2(n_227),
.B1(n_155),
.B2(n_152),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_317),
.A2(n_376),
.B1(n_312),
.B2(n_296),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_251),
.A2(n_230),
.B1(n_189),
.B2(n_200),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_318),
.A2(n_319),
.B1(n_333),
.B2(n_348),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_236),
.A2(n_249),
.B1(n_250),
.B2(n_265),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_330),
.B(n_370),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_249),
.A2(n_229),
.B1(n_202),
.B2(n_147),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_257),
.B(n_155),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_345),
.A2(n_374),
.B(n_286),
.Y(n_413)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_349),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_252),
.B(n_188),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_350),
.B(n_261),
.C(n_248),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_276),
.A2(n_223),
.B1(n_216),
.B2(n_190),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_360),
.A2(n_361),
.B1(n_305),
.B2(n_311),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_266),
.A2(n_172),
.B1(n_215),
.B2(n_152),
.Y(n_361)
);

BUFx24_ASAP7_75t_L g398 ( 
.A(n_363),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_369),
.B(n_298),
.Y(n_418)
);

AND2x2_ASAP7_75t_SL g370 ( 
.A(n_257),
.B(n_201),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_240),
.B(n_181),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_240),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_257),
.A2(n_201),
.B1(n_18),
.B2(n_147),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_375),
.Y(n_379)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_379),
.Y(n_433)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_375),
.Y(n_380)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_380),
.Y(n_438)
);

OA22x2_ASAP7_75t_L g381 ( 
.A1(n_374),
.A2(n_235),
.B1(n_292),
.B2(n_274),
.Y(n_381)
);

OA22x2_ASAP7_75t_L g466 ( 
.A1(n_381),
.A2(n_295),
.B1(n_289),
.B2(n_275),
.Y(n_466)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_375),
.Y(n_382)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_382),
.Y(n_440)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_377),
.Y(n_383)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_383),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_348),
.A2(n_256),
.B1(n_237),
.B2(n_304),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_384),
.A2(n_364),
.B1(n_341),
.B2(n_323),
.Y(n_459)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_377),
.Y(n_385)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_385),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_386),
.B(n_417),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_316),
.B(n_271),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_387),
.B(n_399),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_254),
.Y(n_388)
);

INVxp33_ASAP7_75t_L g444 ( 
.A(n_388),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_SL g432 ( 
.A1(n_389),
.A2(n_404),
.B1(n_420),
.B2(n_427),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_352),
.B(n_308),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_390),
.Y(n_447)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_377),
.Y(n_391)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_391),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_327),
.B(n_301),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_392),
.B(n_396),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_350),
.B(n_306),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_393),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_R g394 ( 
.A(n_339),
.B(n_324),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_394),
.B(n_410),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_339),
.A2(n_235),
.B(n_310),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_395),
.A2(n_378),
.B(n_355),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_327),
.B(n_293),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_320),
.B(n_234),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_320),
.B(n_281),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_400),
.B(n_405),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_339),
.A2(n_235),
.B1(n_310),
.B2(n_281),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_401),
.A2(n_406),
.B1(n_419),
.B2(n_421),
.Y(n_429)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_354),
.Y(n_402)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_402),
.Y(n_452)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_356),
.Y(n_403)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_403),
.Y(n_464)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_357),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_372),
.B(n_235),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_332),
.A2(n_360),
.B1(n_368),
.B2(n_337),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_407),
.B(n_321),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_302),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_408),
.B(n_415),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_368),
.B(n_264),
.C(n_245),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_409),
.B(n_418),
.C(n_346),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_349),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_326),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_414),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_412),
.Y(n_431)
);

NAND2xp33_ASAP7_75t_R g470 ( 
.A(n_413),
.B(n_329),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_356),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_369),
.B(n_302),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_324),
.B(n_259),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_416),
.B(n_423),
.Y(n_456)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_356),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_361),
.A2(n_202),
.B1(n_184),
.B2(n_176),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_328),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_370),
.A2(n_184),
.B1(n_181),
.B2(n_176),
.Y(n_421)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_334),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_422),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_345),
.B(n_291),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_322),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_424),
.B(n_426),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_331),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_357),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_405),
.A2(n_345),
.B1(n_344),
.B2(n_358),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_436),
.A2(n_448),
.B1(n_455),
.B2(n_457),
.Y(n_471)
);

MAJx2_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_370),
.C(n_345),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_443),
.B(n_400),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_406),
.A2(n_322),
.B1(n_342),
.B2(n_347),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_449),
.B(n_407),
.C(n_402),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_454),
.A2(n_470),
.B(n_423),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_401),
.A2(n_342),
.B1(n_347),
.B2(n_362),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_397),
.A2(n_362),
.B1(n_323),
.B2(n_341),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_384),
.A2(n_272),
.B1(n_283),
.B2(n_294),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_458),
.A2(n_389),
.B1(n_419),
.B2(n_421),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_459),
.A2(n_461),
.B1(n_462),
.B2(n_463),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_460),
.B(n_396),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_397),
.A2(n_328),
.B1(n_288),
.B2(n_340),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_397),
.A2(n_340),
.B1(n_284),
.B2(n_378),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_395),
.A2(n_331),
.B1(n_338),
.B2(n_346),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_428),
.A2(n_338),
.B1(n_366),
.B2(n_365),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_465),
.A2(n_468),
.B1(n_469),
.B2(n_385),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_466),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_416),
.A2(n_365),
.B1(n_359),
.B2(n_373),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_425),
.A2(n_359),
.B1(n_371),
.B2(n_373),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_469),
.Y(n_472)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_472),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_474),
.A2(n_482),
.B1(n_496),
.B2(n_436),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_435),
.B(n_392),
.Y(n_475)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_475),
.Y(n_510)
);

OAI21xp33_ASAP7_75t_L g476 ( 
.A1(n_430),
.A2(n_408),
.B(n_413),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_476),
.B(n_489),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_439),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_477),
.B(n_490),
.Y(n_522)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_451),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_478),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_479),
.A2(n_506),
.B(n_466),
.Y(n_537)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_451),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_480),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_481),
.B(n_483),
.C(n_484),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_431),
.A2(n_381),
.B1(n_394),
.B2(n_418),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_409),
.C(n_386),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_439),
.Y(n_485)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_485),
.Y(n_540)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_441),
.Y(n_486)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_486),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_487),
.B(n_438),
.Y(n_526)
);

FAx1_ASAP7_75t_SL g488 ( 
.A(n_443),
.B(n_381),
.CI(n_414),
.CON(n_488),
.SN(n_488)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_488),
.B(n_501),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_446),
.B(n_444),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_437),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_431),
.A2(n_412),
.B1(n_381),
.B2(n_382),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_491),
.A2(n_454),
.B1(n_463),
.B2(n_462),
.Y(n_515)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_492),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_435),
.B(n_380),
.Y(n_493)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_493),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_447),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_494),
.B(n_505),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_449),
.B(n_379),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_495),
.B(n_497),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_446),
.A2(n_403),
.B1(n_417),
.B2(n_411),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g497 ( 
.A(n_453),
.B(n_424),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_453),
.B(n_383),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_498),
.B(n_500),
.C(n_503),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_452),
.B(n_427),
.Y(n_499)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_499),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_443),
.B(n_426),
.C(n_404),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_450),
.B(n_353),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_452),
.B(n_353),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_502),
.B(n_504),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_445),
.B(n_325),
.C(n_336),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_467),
.B(n_325),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_464),
.B(n_391),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_459),
.A2(n_398),
.B1(n_420),
.B2(n_336),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_445),
.B(n_335),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_507),
.B(n_495),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_433),
.B(n_343),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_508),
.B(n_367),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_482),
.A2(n_429),
.B1(n_448),
.B2(n_456),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_511),
.B(n_512),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_509),
.A2(n_429),
.B1(n_456),
.B2(n_434),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_513),
.A2(n_515),
.B1(n_517),
.B2(n_524),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_505),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_514),
.B(n_499),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_509),
.A2(n_458),
.B1(n_434),
.B2(n_465),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_523),
.B(n_526),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_490),
.A2(n_432),
.B1(n_455),
.B2(n_461),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_477),
.A2(n_433),
.B1(n_438),
.B2(n_440),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_525),
.A2(n_528),
.B1(n_486),
.B2(n_474),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_491),
.A2(n_440),
.B1(n_464),
.B2(n_457),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_479),
.A2(n_468),
.B(n_442),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_531),
.A2(n_471),
.B(n_473),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_484),
.B(n_483),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_534),
.B(n_539),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_494),
.A2(n_442),
.B1(n_441),
.B2(n_466),
.Y(n_536)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_536),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_537),
.A2(n_546),
.B(n_488),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_481),
.B(n_466),
.C(n_335),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_538),
.B(n_542),
.C(n_503),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_487),
.B(n_466),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_485),
.A2(n_398),
.B1(n_268),
.B2(n_307),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_541),
.B(n_506),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_500),
.B(n_371),
.C(n_367),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g575 ( 
.A(n_545),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_488),
.A2(n_398),
.B(n_329),
.Y(n_546)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_548),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_549),
.B(n_563),
.Y(n_601)
);

XOR2x2_ASAP7_75t_L g550 ( 
.A(n_519),
.B(n_498),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_550),
.B(n_559),
.Y(n_587)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_522),
.Y(n_551)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_551),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_552),
.B(n_553),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_520),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_522),
.Y(n_554)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_554),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_SL g555 ( 
.A(n_519),
.B(n_497),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_SL g591 ( 
.A(n_555),
.B(n_510),
.Y(n_591)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_525),
.Y(n_557)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_557),
.Y(n_590)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_535),
.Y(n_561)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_561),
.Y(n_594)
);

CKINVDCx16_ASAP7_75t_R g562 ( 
.A(n_543),
.Y(n_562)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_562),
.Y(n_599)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_535),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_518),
.B(n_507),
.C(n_493),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_564),
.B(n_570),
.C(n_576),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g566 ( 
.A(n_533),
.B(n_450),
.Y(n_566)
);

NOR3xp33_ASAP7_75t_L g597 ( 
.A(n_566),
.B(n_567),
.C(n_569),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_531),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_568),
.A2(n_571),
.B1(n_577),
.B2(n_517),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_518),
.B(n_475),
.C(n_480),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_530),
.A2(n_478),
.B1(n_398),
.B2(n_297),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_546),
.A2(n_343),
.B(n_242),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_572),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_537),
.A2(n_539),
.B(n_516),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_574),
.B(n_528),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_534),
.B(n_527),
.C(n_542),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_530),
.A2(n_267),
.B1(n_239),
.B2(n_241),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_540),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_578),
.A2(n_579),
.B1(n_580),
.B2(n_532),
.Y(n_603)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_544),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_547),
.Y(n_580)
);

FAx1_ASAP7_75t_SL g581 ( 
.A(n_564),
.B(n_576),
.CI(n_526),
.CON(n_581),
.SN(n_581)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_581),
.B(n_584),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_570),
.B(n_527),
.C(n_523),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_591),
.B(n_592),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_573),
.B(n_538),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_573),
.B(n_511),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_593),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_595),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_560),
.A2(n_512),
.B1(n_532),
.B2(n_510),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_596),
.A2(n_561),
.B1(n_563),
.B2(n_569),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_565),
.B(n_515),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_598),
.B(n_600),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_565),
.B(n_547),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_602),
.B(n_559),
.C(n_574),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_603),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_SL g604 ( 
.A(n_555),
.B(n_521),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_SL g622 ( 
.A(n_604),
.B(n_541),
.Y(n_622)
);

BUFx24_ASAP7_75t_SL g605 ( 
.A(n_551),
.Y(n_605)
);

CKINVDCx16_ASAP7_75t_R g615 ( 
.A(n_605),
.Y(n_615)
);

CKINVDCx14_ASAP7_75t_R g606 ( 
.A(n_558),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_606),
.B(n_601),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_586),
.A2(n_554),
.B1(n_568),
.B2(n_556),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_607),
.A2(n_617),
.B1(n_595),
.B2(n_585),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_608),
.B(n_594),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_582),
.B(n_550),
.C(n_552),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_610),
.B(n_611),
.C(n_625),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_582),
.B(n_580),
.C(n_558),
.Y(n_611)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_612),
.Y(n_631)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_613),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_583),
.B(n_578),
.Y(n_614)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_614),
.Y(n_634)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_588),
.Y(n_616)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_616),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_596),
.A2(n_549),
.B1(n_572),
.B2(n_571),
.Y(n_617)
);

FAx1_ASAP7_75t_SL g620 ( 
.A(n_591),
.B(n_577),
.CI(n_549),
.CON(n_620),
.SN(n_620)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_620),
.B(n_600),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g629 ( 
.A(n_622),
.B(n_601),
.Y(n_629)
);

INVxp67_ASAP7_75t_SL g623 ( 
.A(n_597),
.Y(n_623)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_623),
.Y(n_641)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_589),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_624),
.B(n_628),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_584),
.B(n_592),
.C(n_593),
.Y(n_625)
);

INVxp33_ASAP7_75t_SL g628 ( 
.A(n_599),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g653 ( 
.A(n_629),
.B(n_622),
.Y(n_653)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_630),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_632),
.B(n_619),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g637 ( 
.A(n_614),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_637),
.B(n_638),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_625),
.B(n_587),
.C(n_598),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_618),
.B(n_602),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_639),
.B(n_642),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_612),
.B(n_590),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_640),
.Y(n_649)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_611),
.B(n_587),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_608),
.B(n_604),
.C(n_581),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_643),
.B(n_646),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_644),
.B(n_647),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_615),
.B(n_553),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_610),
.B(n_575),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_647),
.A2(n_626),
.B(n_609),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_650),
.B(n_653),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_636),
.B(n_627),
.C(n_621),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_652),
.B(n_655),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_654),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_636),
.B(n_619),
.C(n_607),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_641),
.B(n_613),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_656),
.B(n_658),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_644),
.B(n_579),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_642),
.B(n_521),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_661),
.B(n_662),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g662 ( 
.A(n_639),
.B(n_617),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_652),
.B(n_631),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_663),
.B(n_667),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_657),
.A2(n_643),
.B(n_638),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_SL g680 ( 
.A1(n_664),
.A2(n_659),
.B(n_640),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_649),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_651),
.B(n_633),
.C(n_640),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g674 ( 
.A(n_669),
.B(n_673),
.C(n_666),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_655),
.B(n_634),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_670),
.B(n_672),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_648),
.B(n_645),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g684 ( 
.A(n_674),
.B(n_629),
.C(n_529),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_666),
.B(n_660),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_677),
.A2(n_680),
.B(n_681),
.Y(n_682)
);

MAJIxp5_ASAP7_75t_L g678 ( 
.A(n_668),
.B(n_659),
.C(n_662),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_678),
.A2(n_679),
.B(n_665),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_668),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_SL g681 ( 
.A1(n_671),
.A2(n_649),
.B(n_635),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_SL g687 ( 
.A1(n_683),
.A2(n_685),
.B(n_620),
.Y(n_687)
);

MAJIxp5_ASAP7_75t_L g686 ( 
.A(n_684),
.B(n_679),
.C(n_676),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_675),
.A2(n_620),
.B(n_529),
.Y(n_685)
);

OAI21xp5_ASAP7_75t_SL g688 ( 
.A1(n_686),
.A2(n_687),
.B(n_682),
.Y(n_688)
);

AOI21x1_ASAP7_75t_L g689 ( 
.A1(n_688),
.A2(n_303),
.B(n_18),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_SL g690 ( 
.A1(n_689),
.A2(n_18),
.B(n_3),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_690),
.A2(n_3),
.B(n_623),
.Y(n_691)
);


endmodule