module fake_jpeg_10820_n_172 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_172);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_47),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_7),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_19),
.B(n_32),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_4),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_1),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_81),
.Y(n_94)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_1),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_84),
.Y(n_93)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_2),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_2),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_3),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_67),
.B1(n_75),
.B2(n_68),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_68),
.B1(n_67),
.B2(n_57),
.Y(n_103)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_50),
.B(n_68),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_59),
.B(n_53),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_120)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_SL g98 ( 
.A(n_78),
.Y(n_98)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_107),
.B1(n_109),
.B2(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_64),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_14),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_76),
.A3(n_72),
.B1(n_73),
.B2(n_69),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_18),
.C(n_20),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_65),
.B1(n_63),
.B2(n_61),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_120),
.B1(n_48),
.B2(n_23),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_52),
.B1(n_58),
.B2(n_51),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_45),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_56),
.B1(n_49),
.B2(n_50),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_114),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_49),
.B(n_5),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_113),
.C(n_111),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_98),
.C(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_3),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_5),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_115),
.B(n_26),
.Y(n_139)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_12),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_123),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_102),
.B(n_12),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_15),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_17),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_127),
.Y(n_152)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_133),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_44),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_31),
.C(n_35),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_21),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_138),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_140),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_119),
.B(n_27),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_28),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_40),
.Y(n_150)
);

NAND2x1_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_29),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_142),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_144),
.B(n_150),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_153),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_154),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_152),
.B1(n_145),
.B2(n_149),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_161),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_131),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_131),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_136),
.B(n_142),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_159),
.B(n_147),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_163),
.A2(n_143),
.B(n_157),
.Y(n_166)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_163),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_162),
.Y(n_168)
);

AOI31xp67_ASAP7_75t_SL g169 ( 
.A1(n_168),
.A2(n_165),
.A3(n_151),
.B(n_158),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_169),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_160),
.B(n_148),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g172 ( 
.A(n_171),
.Y(n_172)
);


endmodule