module fake_jpeg_11288_n_296 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_296);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_288;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_282;
wire n_258;
wire n_96;

INVxp67_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_33),
.B(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_51),
.Y(n_83)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_0),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_39),
.Y(n_103)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_30),
.B(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_56),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_30),
.B(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_57),
.B(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_31),
.B(n_16),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_70),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_20),
.B(n_14),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_40),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_0),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_27),
.B1(n_19),
.B2(n_38),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_72),
.A2(n_79),
.B1(n_85),
.B2(n_92),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_53),
.A2(n_27),
.B1(n_29),
.B2(n_36),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_87),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_47),
.A2(n_20),
.B1(n_24),
.B2(n_36),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_29),
.B1(n_24),
.B2(n_25),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_35),
.B1(n_19),
.B2(n_38),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_46),
.A2(n_26),
.B1(n_39),
.B2(n_37),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_106),
.Y(n_117)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_65),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_1),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_70),
.A2(n_26),
.B1(n_37),
.B2(n_40),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_7),
.C(n_112),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_55),
.B(n_13),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_107),
.B(n_109),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_51),
.B(n_10),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_45),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_44),
.A2(n_40),
.B1(n_2),
.B2(n_3),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_7),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_119),
.B(n_122),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_1),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_10),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_129),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_8),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_125),
.B(n_126),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_2),
.C(n_5),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_81),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_139),
.Y(n_161)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_7),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_133),
.B(n_91),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_108),
.B1(n_97),
.B2(n_88),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_81),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_136),
.B(n_138),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_94),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_75),
.C(n_102),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_148),
.Y(n_168)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_99),
.Y(n_142)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_77),
.Y(n_145)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_104),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_75),
.B1(n_88),
.B2(n_74),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_SL g204 ( 
.A1(n_149),
.A2(n_132),
.B(n_114),
.Y(n_204)
);

O2A1O1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_142),
.B(n_128),
.C(n_125),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_99),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_162),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_74),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_172),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_159),
.B(n_163),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_91),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_146),
.B(n_76),
.Y(n_163)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_115),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_117),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_176),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_120),
.B(n_108),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_143),
.A2(n_82),
.B1(n_80),
.B2(n_98),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_97),
.B1(n_76),
.B2(n_82),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_175),
.A2(n_177),
.B1(n_159),
.B2(n_164),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_127),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_80),
.B1(n_86),
.B2(n_95),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_179),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_182),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_178),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_183),
.A2(n_123),
.B1(n_150),
.B2(n_114),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_141),
.C(n_134),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_177),
.C(n_172),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_168),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_203),
.Y(n_210)
);

NOR2x1_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_144),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_198),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_170),
.B(n_127),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_192),
.B(n_199),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_171),
.A2(n_145),
.B(n_137),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_153),
.B(n_154),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_137),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_194),
.B(n_175),
.Y(n_211)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_160),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_167),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_204),
.B1(n_160),
.B2(n_152),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_155),
.B(n_116),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_150),
.Y(n_205)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_169),
.B(n_123),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_176),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_217),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_193),
.C(n_181),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_167),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_214),
.B(n_185),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_162),
.B1(n_165),
.B2(n_166),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_218),
.B1(n_186),
.B2(n_195),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_183),
.A2(n_165),
.B1(n_166),
.B2(n_86),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_225),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_187),
.A2(n_154),
.B1(n_197),
.B2(n_184),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_223),
.A2(n_188),
.B1(n_181),
.B2(n_186),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_183),
.B(n_189),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_227),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_231),
.B(n_223),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_202),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_245),
.Y(n_255)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_228),
.B1(n_218),
.B2(n_214),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_196),
.C(n_198),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_209),
.Y(n_254)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_244),
.B1(n_209),
.B2(n_225),
.Y(n_246)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_243),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_207),
.A2(n_185),
.B1(n_200),
.B2(n_190),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_254),
.C(n_238),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_256),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_210),
.B1(n_209),
.B2(n_211),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_252),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_210),
.B1(n_226),
.B2(n_222),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_237),
.Y(n_257)
);

INVx13_ASAP7_75t_L g264 ( 
.A(n_257),
.Y(n_264)
);

OAI21xp33_ASAP7_75t_SL g259 ( 
.A1(n_251),
.A2(n_237),
.B(n_230),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_260),
.Y(n_273)
);

NOR5xp2_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_236),
.C(n_229),
.D(n_231),
.E(n_221),
.Y(n_261)
);

INVx11_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_229),
.C(n_242),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_263),
.C(n_267),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_217),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_230),
.C(n_235),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_246),
.B(n_244),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_276),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_256),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_275),
.Y(n_278)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_267),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_269),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_268),
.B1(n_264),
.B2(n_253),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_234),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_280),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_277),
.A2(n_268),
.B1(n_264),
.B2(n_262),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_282),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_247),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_271),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_274),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_283),
.B(n_273),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_286),
.A2(n_283),
.B(n_278),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_289),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_273),
.B(n_260),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_270),
.A3(n_287),
.B1(n_285),
.B2(n_232),
.C1(n_272),
.C2(n_258),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_272),
.B1(n_235),
.B2(n_239),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_291),
.C(n_243),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_294),
.B(n_212),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_270),
.Y(n_296)
);


endmodule