module fake_netlist_6_2041_n_769 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_769);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_769;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_15),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_107),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_57),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_12),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_27),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_8),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_129),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_30),
.Y(n_168)
);

BUFx8_ASAP7_75t_SL g169 ( 
.A(n_56),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_7),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_61),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_37),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_116),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_97),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_26),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_91),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_112),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_59),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_144),
.Y(n_181)
);

NOR2xp67_ASAP7_75t_L g182 ( 
.A(n_114),
.B(n_15),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_89),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_94),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_54),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_154),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_142),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_6),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_131),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_50),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_120),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_137),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_109),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_48),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_73),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_110),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_49),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_45),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_23),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_103),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_79),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_83),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_88),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_44),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_93),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_75),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_64),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_35),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_68),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_119),
.Y(n_215)
);

OAI22x1_ASAP7_75t_R g216 ( 
.A1(n_166),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_167),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_0),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_175),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_1),
.Y(n_223)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_173),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_159),
.Y(n_226)
);

NOR2x1_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_18),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_177),
.B(n_19),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_172),
.B(n_20),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_172),
.B(n_21),
.Y(n_233)
);

NOR2x1_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_22),
.Y(n_234)
);

AND2x4_ASAP7_75t_L g235 ( 
.A(n_186),
.B(n_24),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_164),
.Y(n_236)
);

OA21x2_ASAP7_75t_L g237 ( 
.A1(n_186),
.A2(n_162),
.B(n_160),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_166),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_163),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_165),
.Y(n_240)
);

OAI22x1_ASAP7_75t_R g241 ( 
.A1(n_161),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_168),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_169),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_161),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_174),
.Y(n_247)
);

OAI21x1_ASAP7_75t_L g248 ( 
.A1(n_176),
.A2(n_80),
.B(n_155),
.Y(n_248)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_180),
.B(n_25),
.Y(n_249)
);

CKINVDCx11_ASAP7_75t_R g250 ( 
.A(n_195),
.Y(n_250)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_181),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

OAI22x1_ASAP7_75t_R g253 ( 
.A1(n_195),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_253)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_183),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_189),
.B(n_8),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_188),
.B(n_9),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_198),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_219),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_225),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_222),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_224),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_222),
.Y(n_267)
);

NAND2xp33_ASAP7_75t_L g268 ( 
.A(n_223),
.B(n_185),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_232),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_228),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_236),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_187),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_207),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_239),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_220),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_220),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g280 ( 
.A1(n_232),
.A2(n_208),
.B(n_214),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_218),
.B(n_209),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_233),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_233),
.Y(n_285)
);

NAND2xp33_ASAP7_75t_SL g286 ( 
.A(n_230),
.B(n_197),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_230),
.B(n_210),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_239),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_251),
.B(n_212),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_220),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_239),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_240),
.Y(n_293)
);

NAND3xp33_ASAP7_75t_L g294 ( 
.A(n_257),
.B(n_215),
.C(n_213),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_245),
.B(n_230),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_229),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_211),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_SL g298 ( 
.A(n_218),
.B(n_197),
.Y(n_298)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_233),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_240),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_220),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_240),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_235),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_231),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_250),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_235),
.Y(n_307)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_244),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_278),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_283),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_288),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_251),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_229),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_269),
.B(n_251),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_278),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_229),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_283),
.A2(n_256),
.B1(n_246),
.B2(n_235),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_273),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_254),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_266),
.B(n_249),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_283),
.B(n_254),
.Y(n_325)
);

NAND3xp33_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_258),
.C(n_249),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_291),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_276),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_292),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_266),
.B(n_249),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_254),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_298),
.A2(n_243),
.B1(n_231),
.B2(n_245),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_273),
.B(n_266),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_285),
.B(n_254),
.Y(n_335)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_262),
.B(n_243),
.Y(n_336)
);

OAI22xp33_ASAP7_75t_L g337 ( 
.A1(n_285),
.A2(n_253),
.B1(n_241),
.B2(n_216),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_266),
.B(n_234),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_293),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_303),
.B(n_221),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_303),
.B(n_307),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_303),
.A2(n_224),
.B1(n_191),
.B2(n_193),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_291),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_276),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_300),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_307),
.B(n_221),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_277),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_301),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_307),
.B(n_221),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_266),
.B(n_221),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_287),
.A2(n_224),
.B1(n_194),
.B2(n_196),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_299),
.B(n_301),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_300),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_276),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_299),
.B(n_244),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_299),
.B(n_237),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_277),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_299),
.B(n_237),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_282),
.B(n_242),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_282),
.B(n_242),
.Y(n_360)
);

NOR3xp33_ASAP7_75t_L g361 ( 
.A(n_263),
.B(n_238),
.C(n_227),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_296),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_299),
.B(n_190),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_299),
.B(n_237),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_282),
.B(n_247),
.Y(n_365)
);

NAND3xp33_ASAP7_75t_L g366 ( 
.A(n_268),
.B(n_247),
.C(n_199),
.Y(n_366)
);

NOR2x1p5_ASAP7_75t_L g367 ( 
.A(n_296),
.B(n_201),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_280),
.B(n_202),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_297),
.B(n_247),
.Y(n_369)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_276),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_302),
.B(n_247),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_302),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_265),
.B(n_238),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_304),
.B(n_203),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_333),
.B(n_268),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_311),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_326),
.A2(n_280),
.B1(n_289),
.B2(n_204),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_304),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_347),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_322),
.A2(n_308),
.B1(n_205),
.B2(n_265),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_373),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_310),
.A2(n_279),
.B(n_274),
.Y(n_382)
);

O2A1O1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_321),
.A2(n_271),
.B(n_272),
.C(n_284),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_336),
.B(n_296),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_313),
.B(n_308),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_356),
.A2(n_364),
.B(n_358),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_313),
.B(n_320),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_314),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_362),
.B(n_305),
.Y(n_389)
);

NAND2x1_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_260),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_357),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_320),
.B(n_305),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_309),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_341),
.A2(n_284),
.B1(n_281),
.B2(n_279),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_369),
.A2(n_274),
.B(n_281),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_368),
.A2(n_260),
.B(n_261),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_261),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_368),
.A2(n_267),
.B(n_264),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_359),
.B(n_360),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_315),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_324),
.A2(n_270),
.B1(n_272),
.B2(n_271),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_355),
.B(n_276),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_337),
.B(n_306),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_351),
.B(n_270),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_372),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_359),
.B(n_264),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_360),
.B(n_367),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_363),
.A2(n_248),
.B1(n_267),
.B2(n_250),
.Y(n_408)
);

O2A1O1Ixp33_ASAP7_75t_L g409 ( 
.A1(n_324),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_319),
.B(n_28),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_327),
.B(n_29),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_330),
.A2(n_306),
.B(n_86),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_330),
.A2(n_85),
.B(n_152),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_316),
.Y(n_414)
);

INVx5_ASAP7_75t_L g415 ( 
.A(n_328),
.Y(n_415)
);

O2A1O1Ixp5_ASAP7_75t_L g416 ( 
.A1(n_338),
.A2(n_363),
.B(n_317),
.C(n_325),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_343),
.B(n_31),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_361),
.B(n_10),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_374),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_342),
.B(n_11),
.Y(n_420)
);

AOI21xp33_ASAP7_75t_L g421 ( 
.A1(n_337),
.A2(n_12),
.B(n_13),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_332),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_348),
.B(n_32),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_318),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_312),
.A2(n_90),
.B(n_151),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_361),
.B(n_13),
.Y(n_426)
);

O2A1O1Ixp33_ASAP7_75t_L g427 ( 
.A1(n_338),
.A2(n_14),
.B(n_16),
.C(n_17),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_323),
.B(n_14),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_329),
.B(n_33),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_334),
.B(n_339),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_345),
.B(n_34),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_353),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_331),
.A2(n_96),
.B(n_150),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_366),
.B(n_16),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_335),
.B(n_328),
.Y(n_435)
);

A2O1A1Ixp33_ASAP7_75t_L g436 ( 
.A1(n_352),
.A2(n_17),
.B(n_36),
.C(n_38),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_340),
.A2(n_39),
.B(n_40),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_346),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_438)
);

O2A1O1Ixp5_ASAP7_75t_L g439 ( 
.A1(n_349),
.A2(n_46),
.B(n_47),
.C(n_51),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_328),
.B(n_52),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_371),
.A2(n_350),
.B(n_370),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_354),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_328),
.B(n_53),
.Y(n_443)
);

NAND2x1p5_ASAP7_75t_L g444 ( 
.A(n_379),
.B(n_354),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_386),
.A2(n_344),
.B(n_354),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_399),
.B(n_354),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_440),
.A2(n_344),
.B(n_58),
.Y(n_447)
);

O2A1O1Ixp5_ASAP7_75t_L g448 ( 
.A1(n_404),
.A2(n_344),
.B(n_60),
.C(n_62),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_381),
.Y(n_449)
);

OA22x2_ASAP7_75t_L g450 ( 
.A1(n_418),
.A2(n_55),
.B1(n_63),
.B2(n_65),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_379),
.B(n_344),
.Y(n_451)
);

BUFx10_ASAP7_75t_L g452 ( 
.A(n_385),
.Y(n_452)
);

AO31x2_ASAP7_75t_L g453 ( 
.A1(n_377),
.A2(n_66),
.A3(n_67),
.B(n_69),
.Y(n_453)
);

A2O1A1Ixp33_ASAP7_75t_L g454 ( 
.A1(n_383),
.A2(n_70),
.B(n_71),
.C(n_72),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_441),
.A2(n_398),
.B(n_396),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_387),
.B(n_74),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_441),
.A2(n_76),
.B(n_77),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_389),
.B(n_78),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_419),
.B(n_81),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_435),
.A2(n_82),
.B(n_84),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_375),
.A2(n_407),
.B1(n_408),
.B2(n_412),
.Y(n_461)
);

OAI21x1_ASAP7_75t_L g462 ( 
.A1(n_396),
.A2(n_87),
.B(n_92),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_406),
.B(n_98),
.Y(n_463)
);

AND3x1_ASAP7_75t_SL g464 ( 
.A(n_421),
.B(n_99),
.C(n_100),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_415),
.A2(n_101),
.B(n_102),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_415),
.A2(n_104),
.B(n_105),
.Y(n_466)
);

O2A1O1Ixp33_ASAP7_75t_L g467 ( 
.A1(n_434),
.A2(n_106),
.B(n_111),
.C(n_113),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_405),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_391),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_415),
.A2(n_115),
.B(n_117),
.Y(n_470)
);

AO31x2_ASAP7_75t_L g471 ( 
.A1(n_398),
.A2(n_436),
.A3(n_394),
.B(n_378),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_382),
.A2(n_118),
.B(n_121),
.Y(n_472)
);

OAI21x1_ASAP7_75t_L g473 ( 
.A1(n_382),
.A2(n_416),
.B(n_395),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_393),
.B(n_397),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_395),
.A2(n_122),
.B(n_123),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_439),
.A2(n_124),
.B(n_126),
.Y(n_476)
);

NOR2x1_ASAP7_75t_SL g477 ( 
.A(n_415),
.B(n_127),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_403),
.Y(n_478)
);

AO31x2_ASAP7_75t_L g479 ( 
.A1(n_401),
.A2(n_130),
.A3(n_132),
.B(n_133),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_376),
.B(n_134),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_402),
.A2(n_136),
.B(n_138),
.Y(n_481)
);

AOI21xp33_ASAP7_75t_L g482 ( 
.A1(n_420),
.A2(n_139),
.B(n_140),
.Y(n_482)
);

NAND2xp33_ASAP7_75t_L g483 ( 
.A(n_410),
.B(n_141),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_388),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_430),
.A2(n_143),
.B(n_145),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_400),
.B(n_146),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_390),
.A2(n_148),
.B(n_149),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_414),
.B(n_157),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_424),
.B(n_432),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_443),
.A2(n_431),
.B(n_429),
.Y(n_490)
);

AO21x2_ASAP7_75t_L g491 ( 
.A1(n_411),
.A2(n_423),
.B(n_417),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_442),
.A2(n_413),
.B(n_433),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_392),
.B(n_426),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_413),
.A2(n_425),
.B(n_433),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_384),
.B(n_428),
.Y(n_495)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_438),
.B(n_380),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_422),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_409),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_427),
.A2(n_425),
.B(n_437),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_387),
.A2(n_399),
.B1(n_419),
.B2(n_407),
.Y(n_500)
);

AOI21xp33_ASAP7_75t_L g501 ( 
.A1(n_385),
.A2(n_321),
.B(n_313),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_450),
.B1(n_496),
.B2(n_461),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_474),
.B(n_500),
.Y(n_503)
);

AO21x2_ASAP7_75t_L g504 ( 
.A1(n_499),
.A2(n_445),
.B(n_494),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_493),
.A2(n_446),
.B1(n_498),
.B2(n_456),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_SL g506 ( 
.A(n_458),
.B(n_459),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_468),
.Y(n_507)
);

AO21x2_ASAP7_75t_L g508 ( 
.A1(n_476),
.A2(n_473),
.B(n_455),
.Y(n_508)
);

AO21x2_ASAP7_75t_L g509 ( 
.A1(n_463),
.A2(n_492),
.B(n_457),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_451),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_469),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_497),
.B(n_452),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_478),
.B(n_449),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_497),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_497),
.A2(n_451),
.B1(n_444),
.B2(n_489),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_462),
.A2(n_472),
.B(n_475),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_487),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_490),
.A2(n_448),
.B(n_486),
.Y(n_518)
);

AO21x1_ASAP7_75t_L g519 ( 
.A1(n_467),
.A2(n_483),
.B(n_482),
.Y(n_519)
);

OA21x2_ASAP7_75t_L g520 ( 
.A1(n_454),
.A2(n_488),
.B(n_480),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_495),
.A2(n_484),
.B1(n_496),
.B2(n_460),
.Y(n_521)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_481),
.A2(n_485),
.B(n_470),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_495),
.B(n_471),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_471),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_477),
.Y(n_525)
);

AO21x2_ASAP7_75t_L g526 ( 
.A1(n_491),
.A2(n_465),
.B(n_466),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_447),
.A2(n_464),
.B(n_479),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_496),
.B(n_479),
.Y(n_528)
);

AOI21x1_ASAP7_75t_L g529 ( 
.A1(n_453),
.A2(n_445),
.B(n_446),
.Y(n_529)
);

INVx6_ASAP7_75t_L g530 ( 
.A(n_479),
.Y(n_530)
);

AOI21x1_ASAP7_75t_L g531 ( 
.A1(n_453),
.A2(n_445),
.B(n_446),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_468),
.B(n_469),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_449),
.Y(n_533)
);

NOR2xp67_ASAP7_75t_L g534 ( 
.A(n_497),
.B(n_362),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_468),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_501),
.A2(n_386),
.B(n_461),
.Y(n_536)
);

OA21x2_ASAP7_75t_L g537 ( 
.A1(n_473),
.A2(n_455),
.B(n_476),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_468),
.Y(n_538)
);

AO21x2_ASAP7_75t_L g539 ( 
.A1(n_499),
.A2(n_445),
.B(n_494),
.Y(n_539)
);

BUFx5_ASAP7_75t_L g540 ( 
.A(n_451),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_449),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_449),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_449),
.Y(n_543)
);

NAND2x1_ASAP7_75t_L g544 ( 
.A(n_525),
.B(n_517),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_502),
.A2(n_536),
.B1(n_532),
.B2(n_523),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_507),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_511),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_535),
.Y(n_548)
);

AO21x2_ASAP7_75t_L g549 ( 
.A1(n_528),
.A2(n_531),
.B(n_529),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_538),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_541),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_510),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_513),
.A2(n_502),
.B1(n_521),
.B2(n_503),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_524),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_524),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_542),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_532),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_540),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_532),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_510),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_510),
.B(n_514),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_510),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_543),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_514),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_543),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_540),
.Y(n_566)
);

OAI21x1_ASAP7_75t_L g567 ( 
.A1(n_516),
.A2(n_517),
.B(n_522),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_540),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_513),
.A2(n_506),
.B1(n_519),
.B2(n_540),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_505),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_540),
.B(n_542),
.Y(n_571)
);

CKINVDCx11_ASAP7_75t_R g572 ( 
.A(n_533),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_515),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_540),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_540),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_539),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_504),
.Y(n_577)
);

OAI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_512),
.A2(n_530),
.B1(n_506),
.B2(n_517),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_539),
.Y(n_579)
);

BUFx4f_ASAP7_75t_L g580 ( 
.A(n_530),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_527),
.B(n_504),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_554),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_554),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_555),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_545),
.B(n_553),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_566),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_559),
.B(n_527),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_546),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_572),
.A2(n_534),
.B1(n_512),
.B2(n_530),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_580),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_555),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_566),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_561),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_559),
.B(n_537),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_576),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_551),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_576),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_571),
.B(n_526),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_580),
.A2(n_520),
.B1(n_508),
.B2(n_526),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_571),
.B(n_520),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_547),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_548),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_550),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_579),
.B(n_509),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_557),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_579),
.B(n_509),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_563),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_570),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_552),
.B(n_522),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_577),
.Y(n_610)
);

NOR2x1_ASAP7_75t_L g611 ( 
.A(n_565),
.B(n_520),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_558),
.B(n_518),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_558),
.B(n_518),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_568),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_556),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_574),
.B(n_552),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_561),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_581),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_573),
.A2(n_569),
.B1(n_572),
.B2(n_581),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_556),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_618),
.B(n_594),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_618),
.B(n_549),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_609),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_596),
.B(n_560),
.Y(n_624)
);

OAI22xp33_ASAP7_75t_L g625 ( 
.A1(n_585),
.A2(n_580),
.B1(n_564),
.B2(n_552),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_593),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_594),
.B(n_549),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_582),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_598),
.B(n_574),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_600),
.B(n_587),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_595),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_607),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_600),
.B(n_575),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_597),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_620),
.B(n_561),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_587),
.B(n_598),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_589),
.A2(n_564),
.B1(n_562),
.B2(n_544),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_598),
.B(n_562),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_614),
.Y(n_639)
);

INVxp67_ASAP7_75t_SL g640 ( 
.A(n_614),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_615),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_597),
.B(n_544),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_610),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_610),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_583),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_609),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_585),
.A2(n_578),
.B1(n_564),
.B2(n_562),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_584),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_591),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_591),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_608),
.B(n_564),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_616),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_604),
.B(n_606),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_619),
.B(n_590),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_630),
.B(n_612),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_631),
.Y(n_656)
);

AND3x1_ASAP7_75t_L g657 ( 
.A(n_635),
.B(n_590),
.C(n_601),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_632),
.B(n_608),
.Y(n_658)
);

NAND2x1_ASAP7_75t_SL g659 ( 
.A(n_623),
.B(n_611),
.Y(n_659)
);

OR2x6_ASAP7_75t_L g660 ( 
.A(n_629),
.B(n_609),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_630),
.B(n_613),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_641),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_631),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_634),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_623),
.B(n_592),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_654),
.B(n_625),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_636),
.B(n_616),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_653),
.B(n_606),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_623),
.B(n_592),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_652),
.B(n_603),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g671 ( 
.A(n_647),
.B(n_605),
.C(n_599),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_634),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_636),
.B(n_617),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_652),
.B(n_588),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_628),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_645),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_628),
.Y(n_677)
);

AND2x2_ASAP7_75t_SL g678 ( 
.A(n_629),
.B(n_586),
.Y(n_678)
);

NOR2x1_ASAP7_75t_L g679 ( 
.A(n_624),
.B(n_602),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_621),
.B(n_612),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_653),
.B(n_604),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_638),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_638),
.B(n_617),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_621),
.B(n_613),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_645),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_656),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_662),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_655),
.B(n_629),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_655),
.B(n_627),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_666),
.B(n_658),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_675),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_668),
.B(n_681),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_682),
.B(n_646),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_675),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_662),
.B(n_633),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_661),
.B(n_627),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_666),
.B(n_679),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_667),
.B(n_633),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_670),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_661),
.B(n_646),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_663),
.Y(n_701)
);

INVxp33_ASAP7_75t_L g702 ( 
.A(n_683),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_664),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_682),
.B(n_622),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_672),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_674),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_676),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_697),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_690),
.B(n_684),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_690),
.B(n_699),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_691),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_689),
.B(n_684),
.Y(n_712)
);

NAND4xp25_ASAP7_75t_L g713 ( 
.A(n_697),
.B(n_671),
.C(n_706),
.D(n_651),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_687),
.A2(n_657),
.B(n_678),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_692),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_696),
.B(n_680),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_688),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_689),
.B(n_680),
.Y(n_718)
);

INVxp67_ASAP7_75t_SL g719 ( 
.A(n_691),
.Y(n_719)
);

OA21x2_ASAP7_75t_L g720 ( 
.A1(n_719),
.A2(n_694),
.B(n_705),
.Y(n_720)
);

AOI21xp33_ASAP7_75t_SL g721 ( 
.A1(n_708),
.A2(n_702),
.B(n_695),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_711),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_713),
.A2(n_710),
.B(n_714),
.C(n_637),
.Y(n_723)
);

OAI22xp33_ASAP7_75t_L g724 ( 
.A1(n_713),
.A2(n_702),
.B1(n_660),
.B2(n_698),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_715),
.B(n_700),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_723),
.B(n_709),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_720),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_L g728 ( 
.A(n_723),
.B(n_590),
.C(n_703),
.Y(n_728)
);

NAND4xp25_ASAP7_75t_L g729 ( 
.A(n_721),
.B(n_707),
.C(n_701),
.D(n_686),
.Y(n_729)
);

AOI22x1_ASAP7_75t_L g730 ( 
.A1(n_722),
.A2(n_694),
.B1(n_693),
.B2(n_718),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_725),
.B(n_712),
.Y(n_731)
);

NAND4xp25_ASAP7_75t_L g732 ( 
.A(n_728),
.B(n_626),
.C(n_593),
.D(n_724),
.Y(n_732)
);

AND4x1_ASAP7_75t_L g733 ( 
.A(n_726),
.B(n_700),
.C(n_673),
.D(n_685),
.Y(n_733)
);

NOR3x1_ASAP7_75t_L g734 ( 
.A(n_729),
.B(n_717),
.C(n_716),
.Y(n_734)
);

AOI221x1_ASAP7_75t_L g735 ( 
.A1(n_727),
.A2(n_693),
.B1(n_643),
.B2(n_644),
.C(n_564),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_731),
.A2(n_693),
.B(n_659),
.C(n_678),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_733),
.B(n_736),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_734),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_738),
.Y(n_739)
);

NOR3xp33_ASAP7_75t_L g740 ( 
.A(n_737),
.B(n_732),
.C(n_646),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_738),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_739),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_741),
.Y(n_743)
);

NOR2x1_ASAP7_75t_L g744 ( 
.A(n_740),
.B(n_720),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_741),
.B(n_735),
.C(n_730),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_741),
.B(n_704),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_743),
.Y(n_747)
);

INVx3_ASAP7_75t_SL g748 ( 
.A(n_742),
.Y(n_748)
);

XNOR2x1_ASAP7_75t_L g749 ( 
.A(n_746),
.B(n_626),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_L g750 ( 
.A(n_745),
.B(n_562),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_744),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_743),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_752),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_747),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_751),
.A2(n_626),
.B(n_677),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_750),
.A2(n_660),
.B1(n_629),
.B2(n_665),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_753),
.A2(n_748),
.B1(n_754),
.B2(n_749),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_755),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_756),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_753),
.Y(n_760)
);

OAI21xp5_ASAP7_75t_L g761 ( 
.A1(n_757),
.A2(n_677),
.B(n_642),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_SL g762 ( 
.A1(n_760),
.A2(n_660),
.B1(n_669),
.B2(n_665),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_758),
.B(n_669),
.Y(n_763)
);

XNOR2xp5_ASAP7_75t_L g764 ( 
.A(n_763),
.B(n_759),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_761),
.A2(n_639),
.B(n_640),
.Y(n_765)
);

OAI21xp5_ASAP7_75t_L g766 ( 
.A1(n_764),
.A2(n_765),
.B(n_762),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_766),
.A2(n_567),
.B(n_650),
.Y(n_767)
);

AOI221xp5_ASAP7_75t_L g768 ( 
.A1(n_767),
.A2(n_648),
.B1(n_649),
.B2(n_650),
.C(n_643),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_768),
.A2(n_648),
.B1(n_649),
.B2(n_665),
.Y(n_769)
);


endmodule