module real_aes_6439_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g536 ( .A1(n_0), .A2(n_186), .B(n_537), .C(n_540), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_1), .B(n_525), .Y(n_541) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
AOI221xp5_ASAP7_75t_L g101 ( .A1(n_3), .A2(n_102), .B1(n_114), .B2(n_739), .C(n_745), .Y(n_101) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_3), .A2(n_750), .B1(n_753), .B2(n_754), .Y(n_749) );
INVx1_ASAP7_75t_L g754 ( .A(n_3), .Y(n_754) );
INVx1_ASAP7_75t_L g204 ( .A(n_4), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_5), .B(n_175), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_6), .A2(n_440), .B(n_519), .Y(n_518) );
AO21x2_ASAP7_75t_L g486 ( .A1(n_7), .A2(n_151), .B(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_8), .A2(n_36), .B1(n_131), .B2(n_140), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_9), .B(n_151), .Y(n_215) );
AND2x6_ASAP7_75t_L g149 ( .A(n_10), .B(n_150), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_11), .A2(n_149), .B(n_443), .C(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_12), .B(n_37), .Y(n_110) );
INVx1_ASAP7_75t_L g147 ( .A(n_13), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_14), .B(n_138), .Y(n_158) );
INVx1_ASAP7_75t_L g196 ( .A(n_15), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_16), .B(n_175), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_17), .B(n_152), .Y(n_220) );
AO32x2_ASAP7_75t_L g183 ( .A1(n_18), .A2(n_148), .A3(n_151), .B1(n_184), .B2(n_188), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_19), .B(n_140), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_20), .B(n_152), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g187 ( .A1(n_21), .A2(n_52), .B1(n_131), .B2(n_140), .Y(n_187) );
AOI22xp33_ASAP7_75t_SL g137 ( .A1(n_22), .A2(n_81), .B1(n_138), .B2(n_140), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_23), .B(n_140), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_24), .A2(n_148), .B(n_443), .C(n_445), .Y(n_442) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_25), .A2(n_148), .B(n_443), .C(n_490), .Y(n_489) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_26), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_27), .B(n_143), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_28), .A2(n_440), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_29), .B(n_143), .Y(n_181) );
INVx2_ASAP7_75t_L g133 ( .A(n_30), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_31), .A2(n_464), .B(n_473), .C(n_475), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_32), .B(n_140), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_33), .B(n_143), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_34), .A2(n_73), .B1(n_116), .B2(n_117), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_34), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_35), .B(n_160), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_38), .B(n_439), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_39), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_40), .B(n_175), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_41), .B(n_440), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_42), .A2(n_464), .B(n_473), .C(n_510), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_43), .A2(n_121), .B1(n_425), .B2(n_426), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_43), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_43), .A2(n_79), .B1(n_425), .B2(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_44), .B(n_140), .Y(n_210) );
INVx1_ASAP7_75t_L g538 ( .A(n_45), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_46), .A2(n_89), .B1(n_131), .B2(n_134), .Y(n_130) );
INVx1_ASAP7_75t_L g511 ( .A(n_47), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_48), .B(n_140), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_49), .B(n_140), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_50), .B(n_440), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_51), .B(n_202), .Y(n_214) );
AOI22xp33_ASAP7_75t_SL g224 ( .A1(n_53), .A2(n_58), .B1(n_138), .B2(n_140), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_54), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_55), .B(n_140), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_56), .B(n_140), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_57), .Y(n_757) );
INVx1_ASAP7_75t_L g150 ( .A(n_59), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_60), .B(n_440), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_61), .B(n_525), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g521 ( .A1(n_62), .A2(n_199), .B(n_202), .C(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_63), .B(n_140), .Y(n_205) );
INVx1_ASAP7_75t_L g146 ( .A(n_64), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_65), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_66), .B(n_175), .Y(n_477) );
AO32x2_ASAP7_75t_L g128 ( .A1(n_67), .A2(n_129), .A3(n_142), .B1(n_148), .B2(n_151), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_68), .B(n_141), .Y(n_501) );
INVx1_ASAP7_75t_L g238 ( .A(n_69), .Y(n_238) );
INVx1_ASAP7_75t_L g173 ( .A(n_70), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g535 ( .A(n_71), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_72), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g117 ( .A(n_73), .Y(n_117) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_74), .A2(n_443), .B(n_460), .C(n_464), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_75), .B(n_138), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g520 ( .A(n_76), .Y(n_520) );
INVx1_ASAP7_75t_L g113 ( .A(n_77), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_78), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_79), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_80), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_82), .B(n_131), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_83), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_84), .B(n_138), .Y(n_178) );
INVx2_ASAP7_75t_L g144 ( .A(n_85), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_86), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_87), .B(n_135), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_88), .B(n_138), .Y(n_211) );
OR2x2_ASAP7_75t_L g106 ( .A(n_90), .B(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g429 ( .A(n_90), .B(n_108), .Y(n_429) );
INVx2_ASAP7_75t_L g726 ( .A(n_90), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_91), .A2(n_100), .B1(n_138), .B2(n_139), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_92), .B(n_440), .Y(n_471) );
INVx1_ASAP7_75t_L g476 ( .A(n_93), .Y(n_476) );
INVxp67_ASAP7_75t_L g523 ( .A(n_94), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_95), .B(n_138), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_96), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g461 ( .A(n_97), .Y(n_461) );
INVx1_ASAP7_75t_L g497 ( .A(n_98), .Y(n_497) );
AND2x2_ASAP7_75t_L g513 ( .A(n_99), .B(n_143), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
OA21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_105), .B(n_111), .Y(n_103) );
NOR2xp33_ASAP7_75t_SL g742 ( .A(n_104), .B(n_112), .Y(n_742) );
INVx1_ASAP7_75t_L g763 ( .A(n_104), .Y(n_763) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g744 ( .A(n_106), .Y(n_744) );
INVx1_ASAP7_75t_SL g748 ( .A(n_106), .Y(n_748) );
INVx1_ASAP7_75t_SL g759 ( .A(n_106), .Y(n_759) );
NOR2x2_ASAP7_75t_L g738 ( .A(n_107), .B(n_726), .Y(n_738) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g725 ( .A(n_108), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x2_ASAP7_75t_L g761 ( .A(n_111), .B(n_762), .Y(n_761) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OAI222xp33_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_118), .B1(n_727), .B2(n_728), .C1(n_734), .C2(n_735), .Y(n_114) );
INVx1_ASAP7_75t_L g727 ( .A(n_115), .Y(n_727) );
INVxp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_427), .B1(n_430), .B2(n_723), .Y(n_119) );
INVx1_ASAP7_75t_L g730 ( .A(n_120), .Y(n_730) );
INVx2_ASAP7_75t_L g426 ( .A(n_121), .Y(n_426) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
XOR2x2_ASAP7_75t_L g750 ( .A(n_122), .B(n_751), .Y(n_750) );
AND3x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_345), .C(n_393), .Y(n_122) );
NOR4xp25_ASAP7_75t_L g123 ( .A(n_124), .B(n_273), .C(n_318), .D(n_332), .Y(n_123) );
OAI311xp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_189), .A3(n_216), .B1(n_226), .C1(n_241), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_153), .Y(n_125) );
OAI21xp33_ASAP7_75t_L g226 ( .A1(n_126), .A2(n_227), .B(n_229), .Y(n_226) );
AND2x2_ASAP7_75t_L g334 ( .A(n_126), .B(n_261), .Y(n_334) );
AND2x2_ASAP7_75t_L g391 ( .A(n_126), .B(n_277), .Y(n_391) );
BUFx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g284 ( .A(n_127), .B(n_182), .Y(n_284) );
AND2x2_ASAP7_75t_L g341 ( .A(n_127), .B(n_289), .Y(n_341) );
INVx1_ASAP7_75t_L g382 ( .A(n_127), .Y(n_382) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_128), .Y(n_250) );
AND2x2_ASAP7_75t_L g291 ( .A(n_128), .B(n_182), .Y(n_291) );
AND2x2_ASAP7_75t_L g295 ( .A(n_128), .B(n_183), .Y(n_295) );
INVx1_ASAP7_75t_L g307 ( .A(n_128), .Y(n_307) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_135), .B1(n_137), .B2(n_141), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx3_ASAP7_75t_L g134 ( .A(n_132), .Y(n_134) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
AND2x6_ASAP7_75t_L g443 ( .A(n_132), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
INVx1_ASAP7_75t_L g203 ( .A(n_133), .Y(n_203) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_134), .Y(n_478) );
INVx2_ASAP7_75t_L g540 ( .A(n_134), .Y(n_540) );
INVx2_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_135), .A2(n_185), .B1(n_186), .B2(n_187), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_135), .A2(n_186), .B1(n_223), .B2(n_224), .Y(n_222) );
INVx4_ASAP7_75t_L g539 ( .A(n_135), .Y(n_539) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx3_ASAP7_75t_L g141 ( .A(n_136), .Y(n_141) );
INVx1_ASAP7_75t_L g160 ( .A(n_136), .Y(n_160) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_136), .Y(n_180) );
AND2x2_ASAP7_75t_L g441 ( .A(n_136), .B(n_203), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_136), .Y(n_444) );
INVx2_ASAP7_75t_L g197 ( .A(n_138), .Y(n_197) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx3_ASAP7_75t_L g172 ( .A(n_140), .Y(n_172) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_140), .Y(n_463) );
INVx5_ASAP7_75t_L g175 ( .A(n_141), .Y(n_175) );
INVx1_ASAP7_75t_L g450 ( .A(n_142), .Y(n_450) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_143), .A2(n_155), .B(n_165), .Y(n_154) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_143), .A2(n_170), .B(n_181), .Y(n_169) );
INVx1_ASAP7_75t_L g453 ( .A(n_143), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_143), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_143), .A2(n_508), .B(n_509), .Y(n_507) );
AND2x2_ASAP7_75t_SL g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x2_ASAP7_75t_L g152 ( .A(n_144), .B(n_145), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
NAND3xp33_ASAP7_75t_L g221 ( .A(n_148), .B(n_222), .C(n_225), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_148), .A2(n_234), .B(n_237), .Y(n_233) );
BUFx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OAI21xp5_ASAP7_75t_L g155 ( .A1(n_149), .A2(n_156), .B(n_161), .Y(n_155) );
OAI21xp5_ASAP7_75t_L g170 ( .A1(n_149), .A2(n_171), .B(n_176), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_149), .A2(n_195), .B(n_200), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_149), .A2(n_209), .B(n_212), .Y(n_208) );
AND2x4_ASAP7_75t_L g440 ( .A(n_149), .B(n_441), .Y(n_440) );
INVx4_ASAP7_75t_SL g465 ( .A(n_149), .Y(n_465) );
NAND2x1p5_ASAP7_75t_L g498 ( .A(n_149), .B(n_441), .Y(n_498) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_151), .A2(n_208), .B(n_215), .Y(n_207) );
INVx4_ASAP7_75t_L g225 ( .A(n_151), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_151), .A2(n_488), .B(n_489), .Y(n_487) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_151), .Y(n_517) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g188 ( .A(n_152), .Y(n_188) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_166), .Y(n_153) );
AND2x2_ASAP7_75t_L g228 ( .A(n_154), .B(n_182), .Y(n_228) );
INVx2_ASAP7_75t_L g262 ( .A(n_154), .Y(n_262) );
AND2x2_ASAP7_75t_L g277 ( .A(n_154), .B(n_183), .Y(n_277) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_154), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_154), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g297 ( .A(n_154), .B(n_260), .Y(n_297) );
INVx1_ASAP7_75t_L g309 ( .A(n_154), .Y(n_309) );
INVx1_ASAP7_75t_L g350 ( .A(n_154), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_154), .B(n_250), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_159), .Y(n_156) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_164), .Y(n_161) );
O2A1O1Ixp5_ASAP7_75t_L g237 ( .A1(n_164), .A2(n_201), .B(n_238), .C(n_239), .Y(n_237) );
NOR2xp67_ASAP7_75t_L g166 ( .A(n_167), .B(n_182), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g227 ( .A(n_168), .B(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_168), .Y(n_255) );
AND2x2_ASAP7_75t_SL g308 ( .A(n_168), .B(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g312 ( .A(n_168), .B(n_182), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_168), .B(n_307), .Y(n_370) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g260 ( .A(n_169), .Y(n_260) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_169), .Y(n_276) );
OR2x2_ASAP7_75t_L g349 ( .A(n_169), .B(n_350), .Y(n_349) );
O2A1O1Ixp5_ASAP7_75t_SL g171 ( .A1(n_172), .A2(n_173), .B(n_174), .C(n_175), .Y(n_171) );
INVx2_ASAP7_75t_L g186 ( .A(n_175), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_175), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_175), .A2(n_235), .B(n_236), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_175), .B(n_523), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_179), .Y(n_176) );
INVx1_ASAP7_75t_L g199 ( .A(n_179), .Y(n_199) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g447 ( .A(n_180), .Y(n_447) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
BUFx2_ASAP7_75t_L g256 ( .A(n_183), .Y(n_256) );
AND2x2_ASAP7_75t_L g261 ( .A(n_183), .B(n_262), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_186), .A2(n_201), .B(n_204), .C(n_205), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_186), .A2(n_213), .B(n_214), .Y(n_212) );
INVx2_ASAP7_75t_L g193 ( .A(n_188), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_188), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_189), .B(n_244), .Y(n_407) );
INVx1_ASAP7_75t_SL g189 ( .A(n_190), .Y(n_189) );
OR2x2_ASAP7_75t_L g377 ( .A(n_190), .B(n_218), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_207), .Y(n_190) );
AND2x2_ASAP7_75t_L g253 ( .A(n_191), .B(n_244), .Y(n_253) );
INVx2_ASAP7_75t_L g265 ( .A(n_191), .Y(n_265) );
AND2x2_ASAP7_75t_L g299 ( .A(n_191), .B(n_247), .Y(n_299) );
AND2x2_ASAP7_75t_L g366 ( .A(n_191), .B(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_192), .B(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g246 ( .A(n_192), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g286 ( .A(n_192), .B(n_207), .Y(n_286) );
AND2x2_ASAP7_75t_L g303 ( .A(n_192), .B(n_304), .Y(n_303) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_206), .Y(n_192) );
OA21x2_ASAP7_75t_L g232 ( .A1(n_193), .A2(n_233), .B(n_240), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_198), .C(n_199), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_197), .A2(n_491), .B(n_492), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_197), .A2(n_501), .B(n_502), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_199), .A2(n_461), .B(n_462), .C(n_463), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_201), .A2(n_446), .B(n_448), .Y(n_445) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g229 ( .A(n_207), .B(n_230), .Y(n_229) );
INVx3_ASAP7_75t_L g247 ( .A(n_207), .Y(n_247) );
AND2x2_ASAP7_75t_L g252 ( .A(n_207), .B(n_232), .Y(n_252) );
AND2x2_ASAP7_75t_L g325 ( .A(n_207), .B(n_304), .Y(n_325) );
AND2x2_ASAP7_75t_L g390 ( .A(n_207), .B(n_380), .Y(n_390) );
OAI311xp33_ASAP7_75t_L g273 ( .A1(n_216), .A2(n_274), .A3(n_278), .B1(n_280), .C1(n_300), .Y(n_273) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g285 ( .A(n_217), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g344 ( .A(n_217), .B(n_252), .Y(n_344) );
AND2x2_ASAP7_75t_L g418 ( .A(n_217), .B(n_299), .Y(n_418) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_218), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g353 ( .A(n_218), .Y(n_353) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx3_ASAP7_75t_L g244 ( .A(n_219), .Y(n_244) );
NOR2x1_ASAP7_75t_L g316 ( .A(n_219), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g373 ( .A(n_219), .B(n_247), .Y(n_373) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
INVx1_ASAP7_75t_L g270 ( .A(n_220), .Y(n_270) );
AO21x1_ASAP7_75t_L g269 ( .A1(n_222), .A2(n_225), .B(n_270), .Y(n_269) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_225), .A2(n_458), .B(n_467), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_225), .B(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_225), .B(n_480), .Y(n_479) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_225), .A2(n_496), .B(n_503), .Y(n_495) );
INVx3_ASAP7_75t_L g525 ( .A(n_225), .Y(n_525) );
AND2x2_ASAP7_75t_L g248 ( .A(n_228), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g301 ( .A(n_228), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g381 ( .A(n_228), .B(n_382), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_229), .A2(n_261), .B1(n_281), .B2(n_285), .C(n_287), .Y(n_280) );
INVx1_ASAP7_75t_L g405 ( .A(n_230), .Y(n_405) );
OR2x2_ASAP7_75t_L g371 ( .A(n_231), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g266 ( .A(n_232), .B(n_247), .Y(n_266) );
OR2x2_ASAP7_75t_L g268 ( .A(n_232), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g293 ( .A(n_232), .Y(n_293) );
INVx2_ASAP7_75t_L g304 ( .A(n_232), .Y(n_304) );
AND2x2_ASAP7_75t_L g331 ( .A(n_232), .B(n_269), .Y(n_331) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_232), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_248), .B1(n_251), .B2(n_254), .C(n_257), .Y(n_241) );
INVx1_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
AND2x2_ASAP7_75t_L g342 ( .A(n_244), .B(n_252), .Y(n_342) );
AND2x2_ASAP7_75t_L g392 ( .A(n_244), .B(n_246), .Y(n_392) );
INVx2_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g279 ( .A(n_246), .B(n_250), .Y(n_279) );
AND2x2_ASAP7_75t_L g358 ( .A(n_246), .B(n_331), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_247), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g317 ( .A(n_247), .Y(n_317) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_248), .A2(n_328), .B(n_330), .Y(n_327) );
OR2x2_ASAP7_75t_L g271 ( .A(n_249), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g337 ( .A(n_249), .B(n_297), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_249), .B(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g314 ( .A(n_250), .B(n_283), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_250), .B(n_397), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_251), .B(n_277), .Y(n_387) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
AND2x2_ASAP7_75t_L g310 ( .A(n_252), .B(n_265), .Y(n_310) );
INVx1_ASAP7_75t_L g326 ( .A(n_253), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_263), .B1(n_267), .B2(n_271), .Y(n_257) );
INVx2_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx2_ASAP7_75t_L g289 ( .A(n_260), .Y(n_289) );
INVx1_ASAP7_75t_L g302 ( .A(n_260), .Y(n_302) );
INVx1_ASAP7_75t_L g272 ( .A(n_261), .Y(n_272) );
AND2x2_ASAP7_75t_L g343 ( .A(n_261), .B(n_289), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_261), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
OR2x2_ASAP7_75t_L g267 ( .A(n_264), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_264), .B(n_380), .Y(n_379) );
NOR2xp67_ASAP7_75t_L g411 ( .A(n_264), .B(n_412), .Y(n_411) );
INVx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g414 ( .A(n_266), .B(n_366), .Y(n_414) );
INVx1_ASAP7_75t_SL g380 ( .A(n_268), .Y(n_380) );
AND2x2_ASAP7_75t_L g320 ( .A(n_269), .B(n_304), .Y(n_320) );
INVx1_ASAP7_75t_L g367 ( .A(n_269), .Y(n_367) );
OAI222xp33_ASAP7_75t_L g408 ( .A1(n_274), .A2(n_364), .B1(n_409), .B2(n_410), .C1(n_413), .C2(n_415), .Y(n_408) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_L g329 ( .A(n_276), .Y(n_329) );
AND2x2_ASAP7_75t_L g340 ( .A(n_277), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_277), .B(n_382), .Y(n_409) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_279), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g384 ( .A(n_281), .Y(n_384) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_SL g322 ( .A(n_284), .Y(n_322) );
AND2x2_ASAP7_75t_L g401 ( .A(n_284), .B(n_362), .Y(n_401) );
AND2x2_ASAP7_75t_L g424 ( .A(n_284), .B(n_308), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_286), .B(n_320), .Y(n_319) );
OAI32xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_290), .A3(n_292), .B1(n_294), .B2(n_298), .Y(n_287) );
BUFx2_ASAP7_75t_L g362 ( .A(n_289), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_290), .B(n_308), .Y(n_389) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g328 ( .A(n_291), .B(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g396 ( .A(n_291), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g385 ( .A(n_292), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AND2x2_ASAP7_75t_L g356 ( .A(n_295), .B(n_329), .Y(n_356) );
INVx2_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
OAI221xp5_ASAP7_75t_SL g318 ( .A1(n_297), .A2(n_319), .B1(n_321), .B2(n_323), .C(n_327), .Y(n_318) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g330 ( .A(n_299), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g336 ( .A(n_299), .B(n_320), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_303), .B1(n_305), .B2(n_310), .C(n_311), .Y(n_300) );
INVx1_ASAP7_75t_L g419 ( .A(n_301), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_302), .B(n_396), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_303), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_308), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g374 ( .A(n_308), .Y(n_374) );
BUFx3_ASAP7_75t_L g397 ( .A(n_309), .Y(n_397) );
INVx1_ASAP7_75t_SL g338 ( .A(n_310), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_310), .B(n_352), .Y(n_351) );
AOI21xp33_ASAP7_75t_SL g311 ( .A1(n_312), .A2(n_313), .B(n_315), .Y(n_311) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_312), .A2(n_413), .B1(n_417), .B2(n_419), .C(n_420), .Y(n_416) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g359 ( .A(n_317), .B(n_320), .Y(n_359) );
INVx1_ASAP7_75t_L g423 ( .A(n_317), .Y(n_423) );
INVx2_ASAP7_75t_L g412 ( .A(n_320), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_320), .B(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g365 ( .A(n_325), .B(n_366), .Y(n_365) );
OAI221xp5_ASAP7_75t_SL g332 ( .A1(n_333), .A2(n_335), .B1(n_337), .B2(n_338), .C(n_339), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_342), .B1(n_343), .B2(n_344), .Y(n_339) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_341), .A2(n_403), .B1(n_404), .B2(n_406), .Y(n_402) );
OAI21xp5_ASAP7_75t_L g420 ( .A1(n_344), .A2(n_421), .B(n_424), .Y(n_420) );
NOR4xp25_ASAP7_75t_SL g345 ( .A(n_346), .B(n_354), .C(n_363), .D(n_383), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_351), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_357), .B1(n_360), .B2(n_361), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g399 ( .A(n_359), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_368), .B1(n_371), .B2(n_374), .C(n_375), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g386 ( .A(n_366), .Y(n_386) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI21xp5_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_378), .B(n_381), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI211xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B(n_387), .C(n_388), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B1(n_391), .B2(n_392), .Y(n_388) );
CKINVDCx14_ASAP7_75t_R g398 ( .A(n_392), .Y(n_398) );
NOR3xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_408), .C(n_416), .Y(n_393) );
OAI221xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_398), .B1(n_399), .B2(n_400), .C(n_402), .Y(n_394) );
INVxp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
CKINVDCx16_ASAP7_75t_R g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g731 ( .A(n_428), .Y(n_731) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g732 ( .A(n_431), .Y(n_732) );
AND3x1_ASAP7_75t_L g431 ( .A(n_432), .B(n_627), .C(n_684), .Y(n_431) );
NOR3xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_572), .C(n_608), .Y(n_432) );
OAI211xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_481), .B(n_527), .C(n_559), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_454), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g530 ( .A(n_436), .B(n_531), .Y(n_530) );
INVx5_ASAP7_75t_L g558 ( .A(n_436), .Y(n_558) );
AND2x2_ASAP7_75t_L g631 ( .A(n_436), .B(n_547), .Y(n_631) );
AND2x2_ASAP7_75t_L g669 ( .A(n_436), .B(n_575), .Y(n_669) );
AND2x2_ASAP7_75t_L g689 ( .A(n_436), .B(n_532), .Y(n_689) );
OR2x6_ASAP7_75t_L g436 ( .A(n_437), .B(n_451), .Y(n_436) );
AOI21xp5_ASAP7_75t_SL g437 ( .A1(n_438), .A2(n_442), .B(n_450), .Y(n_437) );
BUFx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx5_ASAP7_75t_L g474 ( .A(n_443), .Y(n_474) );
INVx2_ASAP7_75t_L g449 ( .A(n_447), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_449), .A2(n_476), .B(n_477), .C(n_478), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_449), .A2(n_478), .B(n_511), .C(n_512), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_454), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_469), .Y(n_454) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_455), .Y(n_570) );
AND2x2_ASAP7_75t_L g584 ( .A(n_455), .B(n_531), .Y(n_584) );
INVx1_ASAP7_75t_L g607 ( .A(n_455), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_455), .B(n_558), .Y(n_646) );
OR2x2_ASAP7_75t_L g683 ( .A(n_455), .B(n_529), .Y(n_683) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_456), .Y(n_619) );
AND2x2_ASAP7_75t_L g626 ( .A(n_456), .B(n_532), .Y(n_626) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g547 ( .A(n_457), .B(n_532), .Y(n_547) );
BUFx2_ASAP7_75t_L g575 ( .A(n_457), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_466), .Y(n_458) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_465), .A2(n_474), .B(n_520), .C(n_521), .Y(n_519) );
O2A1O1Ixp33_ASAP7_75t_SL g534 ( .A1(n_465), .A2(n_474), .B(n_535), .C(n_536), .Y(n_534) );
INVx5_ASAP7_75t_L g529 ( .A(n_469), .Y(n_529) );
BUFx2_ASAP7_75t_L g551 ( .A(n_469), .Y(n_551) );
AND2x2_ASAP7_75t_L g708 ( .A(n_469), .B(n_562), .Y(n_708) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_479), .Y(n_469) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_514), .Y(n_482) );
OAI221xp5_ASAP7_75t_L g608 ( .A1(n_483), .A2(n_609), .B1(n_616), .B2(n_617), .C(n_620), .Y(n_608) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_493), .Y(n_483) );
AND2x2_ASAP7_75t_L g515 ( .A(n_484), .B(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_484), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g543 ( .A(n_485), .B(n_494), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_485), .B(n_495), .Y(n_553) );
OR2x2_ASAP7_75t_L g564 ( .A(n_485), .B(n_516), .Y(n_564) );
AND2x2_ASAP7_75t_L g567 ( .A(n_485), .B(n_555), .Y(n_567) );
AND2x2_ASAP7_75t_L g583 ( .A(n_485), .B(n_505), .Y(n_583) );
OR2x2_ASAP7_75t_L g599 ( .A(n_485), .B(n_495), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_485), .B(n_516), .Y(n_661) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_486), .B(n_505), .Y(n_653) );
AND2x2_ASAP7_75t_L g656 ( .A(n_486), .B(n_495), .Y(n_656) );
OR2x2_ASAP7_75t_L g577 ( .A(n_493), .B(n_564), .Y(n_577) );
INVx2_ASAP7_75t_L g603 ( .A(n_493), .Y(n_603) );
OR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_505), .Y(n_493) );
AND2x2_ASAP7_75t_L g526 ( .A(n_494), .B(n_506), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_494), .B(n_516), .Y(n_582) );
OR2x2_ASAP7_75t_L g593 ( .A(n_494), .B(n_506), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_494), .B(n_555), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_494), .A2(n_686), .B1(n_688), .B2(n_690), .C(n_693), .Y(n_685) );
INVx5_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_495), .B(n_516), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B(n_499), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_505), .B(n_555), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_505), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g571 ( .A(n_505), .B(n_543), .Y(n_571) );
OR2x2_ASAP7_75t_L g615 ( .A(n_505), .B(n_516), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_505), .B(n_567), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_505), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g680 ( .A(n_505), .B(n_681), .Y(n_680) );
INVx5_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_SL g544 ( .A(n_506), .B(n_515), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_SL g548 ( .A1(n_506), .A2(n_549), .B(n_552), .C(n_556), .Y(n_548) );
OR2x2_ASAP7_75t_L g586 ( .A(n_506), .B(n_582), .Y(n_586) );
OR2x2_ASAP7_75t_L g622 ( .A(n_506), .B(n_564), .Y(n_622) );
OAI311xp33_ASAP7_75t_L g628 ( .A1(n_506), .A2(n_567), .A3(n_629), .B1(n_632), .C1(n_639), .Y(n_628) );
AND2x2_ASAP7_75t_L g679 ( .A(n_506), .B(n_516), .Y(n_679) );
AND2x2_ASAP7_75t_L g687 ( .A(n_506), .B(n_542), .Y(n_687) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_506), .Y(n_705) );
AND2x2_ASAP7_75t_L g722 ( .A(n_506), .B(n_543), .Y(n_722) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_513), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_526), .Y(n_514) );
AND2x2_ASAP7_75t_L g550 ( .A(n_515), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g706 ( .A(n_515), .Y(n_706) );
AND2x2_ASAP7_75t_L g542 ( .A(n_516), .B(n_543), .Y(n_542) );
INVx3_ASAP7_75t_L g555 ( .A(n_516), .Y(n_555) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_516), .Y(n_598) );
INVxp67_ASAP7_75t_L g637 ( .A(n_516), .Y(n_637) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_524), .Y(n_516) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_525), .A2(n_533), .B(n_541), .Y(n_532) );
AND2x2_ASAP7_75t_L g715 ( .A(n_526), .B(n_563), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_542), .B1(n_544), .B2(n_545), .C(n_548), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_529), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g568 ( .A(n_529), .B(n_558), .Y(n_568) );
AND2x2_ASAP7_75t_L g576 ( .A(n_529), .B(n_531), .Y(n_576) );
OR2x2_ASAP7_75t_L g588 ( .A(n_529), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g606 ( .A(n_529), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g630 ( .A(n_529), .B(n_631), .Y(n_630) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_529), .Y(n_650) );
AND2x2_ASAP7_75t_L g702 ( .A(n_529), .B(n_626), .Y(n_702) );
OAI31xp33_ASAP7_75t_L g710 ( .A1(n_529), .A2(n_579), .A3(n_678), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_530), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_SL g674 ( .A(n_530), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_530), .B(n_683), .Y(n_682) );
AND2x4_ASAP7_75t_L g562 ( .A(n_531), .B(n_558), .Y(n_562) );
INVx1_ASAP7_75t_L g649 ( .A(n_531), .Y(n_649) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g699 ( .A(n_532), .B(n_558), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_SL g709 ( .A(n_542), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_543), .B(n_614), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_544), .A2(n_656), .B1(n_694), .B2(n_697), .Y(n_693) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g557 ( .A(n_547), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g616 ( .A(n_547), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_547), .B(n_568), .Y(n_721) );
INVx1_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g691 ( .A(n_550), .B(n_692), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_551), .A2(n_610), .B(n_612), .Y(n_609) );
OR2x2_ASAP7_75t_L g617 ( .A(n_551), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g638 ( .A(n_551), .B(n_626), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_551), .B(n_649), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_551), .B(n_689), .Y(n_688) );
OAI221xp5_ASAP7_75t_SL g665 ( .A1(n_552), .A2(n_666), .B1(n_671), .B2(n_674), .C(n_675), .Y(n_665) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
OR2x2_ASAP7_75t_L g642 ( .A(n_553), .B(n_615), .Y(n_642) );
INVx1_ASAP7_75t_L g681 ( .A(n_553), .Y(n_681) );
INVx2_ASAP7_75t_L g657 ( .A(n_554), .Y(n_657) );
INVx1_ASAP7_75t_L g591 ( .A(n_555), .Y(n_591) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g596 ( .A(n_558), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_558), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g625 ( .A(n_558), .B(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g713 ( .A(n_558), .B(n_683), .Y(n_713) );
AOI222xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_563), .B1(n_565), .B2(n_568), .C1(n_569), .C2(n_571), .Y(n_559) );
INVxp67_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g569 ( .A(n_562), .B(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_562), .A2(n_612), .B1(n_640), .B2(n_641), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_562), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
OAI21xp33_ASAP7_75t_SL g600 ( .A1(n_571), .A2(n_601), .B(n_604), .Y(n_600) );
OAI211xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_577), .B(n_578), .C(n_600), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g578 ( .A1(n_576), .A2(n_579), .B1(n_584), .B2(n_585), .C(n_587), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_576), .B(n_664), .Y(n_663) );
INVxp67_ASAP7_75t_L g670 ( .A(n_576), .Y(n_670) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
AND2x2_ASAP7_75t_L g672 ( .A(n_581), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g589 ( .A(n_584), .Y(n_589) );
AND2x2_ASAP7_75t_L g595 ( .A(n_584), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_590), .B1(n_594), .B2(n_597), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_591), .B(n_603), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_592), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g692 ( .A(n_596), .Y(n_692) );
AND2x2_ASAP7_75t_L g711 ( .A(n_596), .B(n_626), .Y(n_711) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_603), .B(n_660), .Y(n_719) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_606), .B(n_674), .Y(n_717) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g640 ( .A(n_618), .Y(n_640) );
BUFx2_ASAP7_75t_L g664 ( .A(n_619), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_623), .B(n_625), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR3xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_643), .C(n_665), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B(n_638), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
A2O1A1Ixp33_ASAP7_75t_SL g643 ( .A1(n_644), .A2(n_647), .B(n_651), .C(n_654), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_644), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NOR2xp67_ASAP7_75t_SL g648 ( .A(n_649), .B(n_650), .Y(n_648) );
OR2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_SL g673 ( .A(n_653), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_658), .B(n_662), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
AND2x2_ASAP7_75t_L g678 ( .A(n_656), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .B1(n_680), .B2(n_682), .Y(n_675) );
INVx2_ASAP7_75t_SL g696 ( .A(n_683), .Y(n_696) );
NOR3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_700), .C(n_712), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_696), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B1(n_707), .B2(n_709), .C(n_710), .Y(n_700) );
A2O1A1Ixp33_ASAP7_75t_L g712 ( .A1(n_701), .A2(n_713), .B(n_714), .C(n_716), .Y(n_712) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVxp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_720), .B2(n_722), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g733 ( .A(n_724), .Y(n_733) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_730), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_729) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
BUFx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND2xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
AOI21xp33_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_755), .B(n_760), .Y(n_745) );
INVxp33_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g753 ( .A(n_750), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
endmodule