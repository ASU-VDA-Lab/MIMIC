module fake_jpeg_31850_n_208 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_208);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_34),
.Y(n_59)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_37),
.B(n_27),
.Y(n_82)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_13),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_49),
.B(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_14),
.B(n_1),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_32),
.B(n_30),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_78),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_55),
.B(n_63),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_16),
.B1(n_30),
.B2(n_26),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_58),
.A2(n_60),
.B1(n_81),
.B2(n_9),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_16),
.B1(n_30),
.B2(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_35),
.B(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_14),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_64),
.B(n_67),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_19),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_15),
.Y(n_76)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_15),
.B1(n_23),
.B2(n_21),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_36),
.A2(n_28),
.B1(n_25),
.B2(n_23),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_33),
.B(n_28),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_82),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_26),
.B1(n_28),
.B2(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_27),
.Y(n_84)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_34),
.B(n_27),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_34),
.B(n_1),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_88),
.A2(n_2),
.B(n_3),
.Y(n_94)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_55),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_77),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_113),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

NAND2x1_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_5),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_104),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_88),
.B1(n_75),
.B2(n_56),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_53),
.B1(n_89),
.B2(n_54),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_54),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_109),
.A2(n_112),
.B1(n_52),
.B2(n_66),
.Y(n_121)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_115),
.Y(n_128)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_119),
.Y(n_143)
);

NAND2x1_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_82),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_59),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_120),
.B(n_126),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_80),
.B(n_63),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_123),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_127),
.B1(n_130),
.B2(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_68),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_86),
.B1(n_56),
.B2(n_73),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_101),
.A2(n_104),
.B1(n_95),
.B2(n_111),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_65),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_100),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_73),
.B1(n_52),
.B2(n_66),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_65),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_136),
.B(n_91),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_72),
.B1(n_62),
.B2(n_70),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_110),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_97),
.A2(n_72),
.B1(n_69),
.B2(n_70),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_107),
.A2(n_12),
.B1(n_69),
.B2(n_114),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_133),
.A2(n_130),
.B1(n_122),
.B2(n_124),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

XOR2x1_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_122),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_141),
.A2(n_131),
.B1(n_117),
.B2(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_142),
.B(n_148),
.Y(n_160)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_105),
.C(n_102),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_156),
.C(n_151),
.Y(n_159)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_154),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_90),
.B1(n_92),
.B2(n_110),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_99),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_115),
.B1(n_106),
.B2(n_113),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_127),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_159),
.B(n_161),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_136),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_118),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_170),
.Y(n_176)
);

OA21x2_ASAP7_75t_SL g180 ( 
.A1(n_164),
.A2(n_138),
.B(n_116),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_152),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_165),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_134),
.B(n_121),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_169),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_156),
.C(n_153),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_162),
.C(n_166),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_155),
.B1(n_146),
.B2(n_140),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_175),
.B1(n_180),
.B2(n_164),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_155),
.B1(n_147),
.B2(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_118),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_179),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_166),
.A2(n_149),
.B1(n_141),
.B2(n_128),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_186),
.C(n_188),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_128),
.Y(n_184)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_174),
.B1(n_179),
.B2(n_180),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_162),
.C(n_168),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_176),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_168),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_173),
.C(n_135),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_193),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_183),
.A2(n_175),
.B1(n_169),
.B2(n_172),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_186),
.C(n_182),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_199),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_172),
.C(n_125),
.Y(n_199)
);

AOI211xp5_ASAP7_75t_SL g200 ( 
.A1(n_191),
.A2(n_120),
.B(n_12),
.C(n_69),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_135),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_201),
.A2(n_132),
.B(n_196),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_197),
.Y(n_203)
);

NOR2xp67_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_198),
.Y(n_205)
);

INVxp67_ASAP7_75t_SL g206 ( 
.A(n_204),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_202),
.C(n_205),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_98),
.Y(n_208)
);


endmodule