module fake_netlist_6_3026_n_1567 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1567);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1567;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_226;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_245;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1069;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1398;
wire n_1201;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_302;
wire n_380;
wire n_1535;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_90),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_32),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_174),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_189),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_224),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_28),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_85),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_16),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_11),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_146),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_48),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_40),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_135),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_139),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_2),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_134),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_128),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_71),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_107),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_152),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_87),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_214),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_19),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_76),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_200),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_39),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_204),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_82),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_193),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_121),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_56),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_109),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_70),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_158),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_89),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_10),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_182),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_98),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_197),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_80),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_36),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_212),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_209),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_123),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_3),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_223),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_52),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_157),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_15),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_207),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_10),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_210),
.Y(n_277)
);

BUFx2_ASAP7_75t_SL g278 ( 
.A(n_8),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_92),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_165),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_145),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_177),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_88),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_216),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_172),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_213),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_14),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_173),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_43),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_4),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_220),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_183),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_112),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_7),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_2),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_9),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_49),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_101),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_81),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_162),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_54),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_86),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_164),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_19),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_120),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_110),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_178),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_39),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_133),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_141),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_67),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_99),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_58),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_23),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_222),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_37),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_202),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_62),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_114),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_91),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_117),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_206),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_106),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_142),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_148),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_196),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_111),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_27),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_124),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_84),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_40),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_199),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_24),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_160),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_143),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_55),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_176),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_108),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_5),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_122),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_100),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_79),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_20),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_211),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_9),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_31),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_136),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_43),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_29),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_27),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_140),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_3),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_14),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_192),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_104),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_44),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_68),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_4),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_97),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_48),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_96),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_191),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_34),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_95),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_42),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_18),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_24),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_297),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_289),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_289),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_233),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_297),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_297),
.B(n_0),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_259),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_225),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_363),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_229),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_271),
.B(n_0),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_363),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_227),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_287),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_351),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_363),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_235),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_249),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_287),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_250),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_252),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_255),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_229),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_294),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_260),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_351),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_294),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_261),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_266),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_263),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_268),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_268),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_286),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_288),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_309),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_243),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_243),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_270),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_274),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_257),
.B(n_1),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_291),
.B(n_1),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_286),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_276),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_280),
.B(n_6),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_290),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_267),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_292),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_269),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_278),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_362),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_365),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_304),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_292),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_273),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_307),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_277),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_328),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_282),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_283),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g427 ( 
.A(n_240),
.B(n_6),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_346),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_358),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_228),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_360),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_367),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_232),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_307),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_239),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_243),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_R g437 ( 
.A(n_330),
.B(n_50),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_253),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_365),
.B(n_7),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_330),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_254),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_361),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_256),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_251),
.Y(n_444)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_226),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_361),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_293),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_231),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_258),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_302),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_300),
.B(n_8),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_236),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_403),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_444),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_371),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_451),
.B(n_340),
.Y(n_456)
);

OA21x2_ASAP7_75t_L g457 ( 
.A1(n_403),
.A2(n_349),
.B(n_310),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_404),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_404),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_436),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_436),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_382),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_373),
.B(n_300),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_368),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_382),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_433),
.B(n_303),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_372),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_435),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_382),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_438),
.B(n_303),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_441),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_382),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_323),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_449),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_395),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_430),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_430),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_396),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_405),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_406),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_410),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_412),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_393),
.B(n_323),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_419),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_379),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_424),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_428),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_429),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_431),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_432),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_393),
.B(n_310),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_381),
.B(n_349),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_386),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_411),
.B(n_230),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_391),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_378),
.B(n_317),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_394),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_427),
.B(n_262),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_SL g499 ( 
.A(n_437),
.B(n_234),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_417),
.B(n_230),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_416),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_407),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_375),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_380),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_408),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_384),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_383),
.B(n_264),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_418),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_385),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_387),
.B(n_388),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_389),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_392),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_397),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_413),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_415),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_421),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_439),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_423),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_425),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_376),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_426),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_390),
.Y(n_522)
);

AO22x2_ASAP7_75t_L g523 ( 
.A1(n_505),
.A2(n_234),
.B1(n_353),
.B2(n_272),
.Y(n_523)
);

NAND2x1p5_ASAP7_75t_L g524 ( 
.A(n_457),
.B(n_265),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_453),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_462),
.B(n_275),
.Y(n_526)
);

NOR3xp33_ASAP7_75t_L g527 ( 
.A(n_496),
.B(n_401),
.C(n_374),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_485),
.B(n_402),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_453),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_458),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_485),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_458),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_496),
.B(n_445),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_458),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_458),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_453),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_461),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_491),
.B(n_483),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_476),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_461),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_461),
.Y(n_541)
);

NAND2x1p5_ASAP7_75t_L g542 ( 
.A(n_457),
.B(n_279),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_479),
.Y(n_543)
);

AND2x6_ASAP7_75t_L g544 ( 
.A(n_502),
.B(n_281),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_456),
.B(n_447),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_479),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_460),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_460),
.Y(n_548)
);

NAND2x1p5_ASAP7_75t_L g549 ( 
.A(n_457),
.B(n_284),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_479),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_491),
.B(n_450),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_502),
.B(n_313),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_479),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_505),
.A2(n_366),
.B1(n_452),
.B2(n_448),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_454),
.B(n_448),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_460),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_476),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_502),
.B(n_315),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_458),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_491),
.B(n_285),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_502),
.B(n_318),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_454),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_460),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_458),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_457),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_476),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_457),
.Y(n_567)
);

AND2x2_ASAP7_75t_SL g568 ( 
.A(n_502),
.B(n_298),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_502),
.B(n_319),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_502),
.A2(n_335),
.B1(n_359),
.B2(n_299),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_493),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_458),
.Y(n_572)
);

AND3x4_ASAP7_75t_L g573 ( 
.A(n_501),
.B(n_370),
.C(n_369),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_501),
.B(n_237),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_522),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_483),
.B(n_301),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_483),
.B(n_306),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_459),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_459),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_459),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_515),
.Y(n_581)
);

NAND2x1p5_ASAP7_75t_L g582 ( 
.A(n_515),
.B(n_311),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_459),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_568),
.B(n_511),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_543),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_543),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_546),
.Y(n_587)
);

AO22x2_ASAP7_75t_L g588 ( 
.A1(n_573),
.A2(n_517),
.B1(n_522),
.B2(n_494),
.Y(n_588)
);

AO22x2_ASAP7_75t_L g589 ( 
.A1(n_573),
.A2(n_517),
.B1(n_494),
.B2(n_463),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_546),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_533),
.B(n_515),
.Y(n_591)
);

OAI221xp5_ASAP7_75t_L g592 ( 
.A1(n_545),
.A2(n_473),
.B1(n_466),
.B2(n_500),
.C(n_499),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_568),
.B(n_511),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_550),
.Y(n_594)
);

OAI221xp5_ASAP7_75t_L g595 ( 
.A1(n_570),
.A2(n_466),
.B1(n_473),
.B2(n_500),
.C(n_497),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_550),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_553),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_531),
.Y(n_598)
);

CKINVDCx14_ASAP7_75t_R g599 ( 
.A(n_528),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_553),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_571),
.Y(n_601)
);

NAND2xp33_ASAP7_75t_L g602 ( 
.A(n_581),
.B(n_515),
.Y(n_602)
);

BUFx8_ASAP7_75t_L g603 ( 
.A(n_528),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_575),
.Y(n_604)
);

AO22x2_ASAP7_75t_L g605 ( 
.A1(n_573),
.A2(n_463),
.B1(n_512),
.B2(n_506),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_538),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_538),
.Y(n_607)
);

NAND2x1p5_ASAP7_75t_L g608 ( 
.A(n_551),
.B(n_515),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_568),
.B(n_511),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_526),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_551),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_526),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_576),
.A2(n_503),
.B1(n_509),
.B2(n_504),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_562),
.B(n_510),
.Y(n_614)
);

AO22x2_ASAP7_75t_L g615 ( 
.A1(n_554),
.A2(n_463),
.B1(n_512),
.B2(n_506),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_552),
.B(n_511),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_574),
.Y(n_617)
);

NAND2x1p5_ASAP7_75t_L g618 ( 
.A(n_526),
.B(n_515),
.Y(n_618)
);

AND2x6_ASAP7_75t_SL g619 ( 
.A(n_577),
.B(n_510),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_526),
.Y(n_620)
);

AO22x2_ASAP7_75t_L g621 ( 
.A1(n_555),
.A2(n_463),
.B1(n_519),
.B2(n_498),
.Y(n_621)
);

AO22x2_ASAP7_75t_L g622 ( 
.A1(n_527),
.A2(n_463),
.B1(n_519),
.B2(n_498),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_547),
.Y(n_623)
);

AO22x2_ASAP7_75t_L g624 ( 
.A1(n_523),
.A2(n_498),
.B1(n_504),
.B2(n_503),
.Y(n_624)
);

AO22x2_ASAP7_75t_L g625 ( 
.A1(n_523),
.A2(n_498),
.B1(n_504),
.B2(n_503),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_560),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_560),
.B(n_509),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_L g628 ( 
.A(n_544),
.B(n_515),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_556),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_577),
.B(n_509),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_547),
.Y(n_631)
);

NAND2x1p5_ASAP7_75t_L g632 ( 
.A(n_539),
.B(n_516),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_556),
.Y(n_633)
);

AO22x2_ASAP7_75t_L g634 ( 
.A1(n_523),
.A2(n_498),
.B1(n_518),
.B2(n_513),
.Y(n_634)
);

AO22x2_ASAP7_75t_L g635 ( 
.A1(n_523),
.A2(n_513),
.B1(n_521),
.B2(n_518),
.Y(n_635)
);

AO22x2_ASAP7_75t_L g636 ( 
.A1(n_523),
.A2(n_513),
.B1(n_521),
.B2(n_518),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_574),
.B(n_521),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_563),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_558),
.B(n_514),
.Y(n_639)
);

AO22x2_ASAP7_75t_L g640 ( 
.A1(n_565),
.A2(n_501),
.B1(n_322),
.B2(n_324),
.Y(n_640)
);

OAI22xp33_ASAP7_75t_SL g641 ( 
.A1(n_561),
.A2(n_514),
.B1(n_520),
.B2(n_508),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_569),
.A2(n_514),
.B1(n_516),
.B2(n_544),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_565),
.B(n_514),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_565),
.B(n_516),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_567),
.B(n_520),
.Y(n_645)
);

OAI221xp5_ASAP7_75t_L g646 ( 
.A1(n_582),
.A2(n_495),
.B1(n_497),
.B2(n_475),
.C(n_482),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_563),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_567),
.B(n_516),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_544),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_525),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_525),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_582),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_536),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_539),
.B(n_495),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_544),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_536),
.Y(n_656)
);

NAND2x1p5_ASAP7_75t_L g657 ( 
.A(n_539),
.B(n_516),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_567),
.B(n_516),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_537),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_582),
.Y(n_660)
);

BUFx8_ASAP7_75t_L g661 ( 
.A(n_544),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_540),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_540),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_541),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_541),
.Y(n_665)
);

AO22x2_ASAP7_75t_L g666 ( 
.A1(n_572),
.A2(n_326),
.B1(n_336),
.B2(n_312),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_547),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_637),
.B(n_516),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_584),
.B(n_524),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_SL g670 ( 
.A(n_611),
.B(n_409),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_637),
.B(n_476),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_627),
.B(n_476),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_627),
.B(n_544),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_630),
.B(n_477),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_630),
.B(n_477),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_614),
.B(n_477),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_598),
.B(n_477),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_613),
.B(n_477),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_617),
.B(n_477),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_645),
.B(n_477),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_608),
.B(n_508),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_606),
.B(n_455),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_607),
.B(n_455),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_641),
.B(n_604),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_593),
.B(n_434),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_609),
.B(n_440),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_626),
.B(n_544),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_SL g688 ( 
.A(n_591),
.B(n_377),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_660),
.B(n_377),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_639),
.B(n_398),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_654),
.B(n_398),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_654),
.B(n_399),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_616),
.B(n_399),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_644),
.B(n_544),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_642),
.B(n_618),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_652),
.B(n_610),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_612),
.B(n_400),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_SL g698 ( 
.A(n_655),
.B(n_400),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_SL g699 ( 
.A(n_620),
.B(n_414),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_643),
.B(n_414),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_SL g701 ( 
.A(n_648),
.B(n_420),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_658),
.B(n_507),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_632),
.B(n_420),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_657),
.B(n_422),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_585),
.B(n_422),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_602),
.B(n_507),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_SL g707 ( 
.A(n_586),
.B(n_442),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_587),
.B(n_442),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_590),
.B(n_446),
.Y(n_709)
);

NAND2xp33_ASAP7_75t_SL g710 ( 
.A(n_594),
.B(n_446),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_596),
.B(n_470),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_597),
.B(n_470),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_SL g713 ( 
.A(n_600),
.B(n_238),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_601),
.B(n_470),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_SL g715 ( 
.A(n_619),
.B(n_241),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_SL g716 ( 
.A(n_629),
.B(n_241),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_633),
.B(n_242),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_638),
.B(n_507),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_647),
.B(n_242),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_592),
.B(n_507),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_650),
.B(n_507),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_651),
.B(n_244),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_653),
.B(n_244),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_656),
.B(n_245),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_659),
.B(n_246),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_SL g726 ( 
.A(n_615),
.B(n_246),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_SL g727 ( 
.A(n_615),
.B(n_247),
.Y(n_727)
);

NAND2xp33_ASAP7_75t_SL g728 ( 
.A(n_662),
.B(n_247),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_SL g729 ( 
.A(n_663),
.B(n_305),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_664),
.B(n_305),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_649),
.B(n_557),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_665),
.B(n_493),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_667),
.B(n_493),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_SL g734 ( 
.A(n_605),
.B(n_320),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_623),
.B(n_493),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_631),
.B(n_579),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_603),
.B(n_579),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_599),
.B(n_492),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_661),
.B(n_579),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_661),
.B(n_579),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_588),
.B(n_492),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_SL g742 ( 
.A(n_605),
.B(n_321),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_595),
.B(n_507),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_621),
.B(n_579),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_621),
.B(n_579),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_622),
.B(n_557),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_589),
.B(n_468),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_589),
.B(n_468),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_622),
.B(n_468),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_588),
.B(n_471),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_624),
.B(n_471),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_624),
.B(n_471),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_625),
.B(n_474),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_SL g754 ( 
.A(n_625),
.B(n_325),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_SL g755 ( 
.A(n_634),
.B(n_327),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_635),
.B(n_507),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_635),
.B(n_636),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_634),
.B(n_474),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_SL g759 ( 
.A(n_636),
.B(n_329),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_646),
.B(n_474),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_640),
.B(n_507),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_628),
.B(n_524),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_738),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_670),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_698),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_690),
.B(n_492),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_SL g767 ( 
.A(n_746),
.B(n_507),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_SL g768 ( 
.A(n_688),
.B(n_370),
.C(n_369),
.Y(n_768)
);

A2O1A1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_720),
.A2(n_354),
.B(n_341),
.C(n_344),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_694),
.A2(n_542),
.B(n_524),
.Y(n_770)
);

O2A1O1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_750),
.A2(n_364),
.B(n_488),
.C(n_482),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_743),
.A2(n_583),
.B(n_578),
.C(n_572),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_741),
.B(n_640),
.Y(n_773)
);

AND2x2_ASAP7_75t_SL g774 ( 
.A(n_746),
.B(n_462),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_731),
.B(n_542),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_701),
.A2(n_583),
.B(n_578),
.C(n_557),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_757),
.A2(n_542),
.B1(n_549),
.B2(n_666),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_SL g778 ( 
.A(n_685),
.B(n_332),
.Y(n_778)
);

BUFx12f_ASAP7_75t_L g779 ( 
.A(n_746),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_762),
.A2(n_549),
.B(n_578),
.Y(n_780)
);

OAI21x1_ASAP7_75t_L g781 ( 
.A1(n_762),
.A2(n_549),
.B(n_532),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_671),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_751),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_686),
.B(n_475),
.Y(n_784)
);

NAND2x1p5_ASAP7_75t_L g785 ( 
.A(n_739),
.B(n_566),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_752),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_702),
.A2(n_532),
.B(n_530),
.Y(n_787)
);

AOI21x1_ASAP7_75t_L g788 ( 
.A1(n_669),
.A2(n_666),
.B(n_548),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_695),
.A2(n_580),
.B(n_566),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_669),
.A2(n_580),
.B(n_566),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_696),
.B(n_486),
.Y(n_791)
);

AO31x2_ASAP7_75t_L g792 ( 
.A1(n_761),
.A2(n_472),
.A3(n_469),
.B(n_465),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_756),
.A2(n_529),
.B(n_530),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_731),
.Y(n_794)
);

AO31x2_ASAP7_75t_L g795 ( 
.A1(n_706),
.A2(n_721),
.A3(n_718),
.B(n_687),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_753),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_711),
.B(n_530),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_712),
.B(n_530),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_668),
.A2(n_580),
.B(n_534),
.Y(n_799)
);

NAND2x1p5_ASAP7_75t_L g800 ( 
.A(n_740),
.B(n_580),
.Y(n_800)
);

O2A1O1Ixp5_ASAP7_75t_SL g801 ( 
.A1(n_747),
.A2(n_465),
.B(n_469),
.C(n_472),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_680),
.A2(n_534),
.B(n_532),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_758),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_731),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_672),
.A2(n_534),
.B(n_532),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_674),
.A2(n_535),
.B(n_534),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_748),
.A2(n_745),
.B(n_744),
.Y(n_807)
);

AOI21x1_ASAP7_75t_SL g808 ( 
.A1(n_673),
.A2(n_755),
.B(n_754),
.Y(n_808)
);

AOI221x1_ASAP7_75t_L g809 ( 
.A1(n_726),
.A2(n_486),
.B1(n_487),
.B2(n_488),
.C(n_535),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_714),
.B(n_564),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_693),
.B(n_487),
.Y(n_811)
);

OAI21x1_ASAP7_75t_L g812 ( 
.A1(n_736),
.A2(n_559),
.B(n_535),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_735),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_749),
.A2(n_529),
.B(n_535),
.Y(n_814)
);

OAI21x1_ASAP7_75t_L g815 ( 
.A1(n_733),
.A2(n_564),
.B(n_559),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_700),
.B(n_334),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_676),
.B(n_559),
.Y(n_817)
);

AOI221x1_ASAP7_75t_L g818 ( 
.A1(n_727),
.A2(n_564),
.B1(n_559),
.B2(n_489),
.C(n_481),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_760),
.A2(n_564),
.B(n_529),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_678),
.A2(n_548),
.B(n_467),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_681),
.B(n_464),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_722),
.B(n_464),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_675),
.A2(n_679),
.B(n_677),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_759),
.A2(n_732),
.B(n_684),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_691),
.B(n_478),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_715),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_737),
.B(n_478),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_692),
.B(n_478),
.Y(n_828)
);

AO21x1_ASAP7_75t_L g829 ( 
.A1(n_734),
.A2(n_548),
.B(n_467),
.Y(n_829)
);

OAI21xp5_ASAP7_75t_L g830 ( 
.A1(n_717),
.A2(n_481),
.B(n_480),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_719),
.A2(n_724),
.B(n_723),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_SL g832 ( 
.A1(n_707),
.A2(n_248),
.B1(n_295),
.B2(n_296),
.Y(n_832)
);

BUFx10_ASAP7_75t_L g833 ( 
.A(n_710),
.Y(n_833)
);

A2O1A1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_742),
.A2(n_480),
.B(n_489),
.C(n_338),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_725),
.A2(n_459),
.B(n_342),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_730),
.A2(n_489),
.B(n_243),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_682),
.B(n_484),
.Y(n_837)
);

O2A1O1Ixp5_ASAP7_75t_SL g838 ( 
.A1(n_697),
.A2(n_243),
.B(n_308),
.C(n_314),
.Y(n_838)
);

OAI21x1_ASAP7_75t_SL g839 ( 
.A1(n_699),
.A2(n_130),
.B(n_159),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_703),
.A2(n_459),
.B(n_357),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_683),
.B(n_316),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_713),
.A2(n_347),
.B(n_337),
.C(n_355),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_704),
.A2(n_689),
.B(n_708),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_705),
.B(n_484),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_709),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_716),
.A2(n_348),
.B(n_331),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_L g847 ( 
.A(n_728),
.B(n_51),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_729),
.Y(n_848)
);

AO31x2_ASAP7_75t_L g849 ( 
.A1(n_720),
.A2(n_243),
.A3(n_12),
.B(n_13),
.Y(n_849)
);

CKINVDCx6p67_ASAP7_75t_R g850 ( 
.A(n_738),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_738),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_701),
.A2(n_490),
.B1(n_484),
.B2(n_243),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_750),
.A2(n_333),
.B(n_339),
.C(n_343),
.Y(n_853)
);

AO31x2_ASAP7_75t_L g854 ( 
.A1(n_720),
.A2(n_11),
.A3(n_12),
.B(n_13),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_731),
.B(n_484),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_787),
.A2(n_459),
.B(n_125),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_779),
.Y(n_857)
);

INVx6_ASAP7_75t_L g858 ( 
.A(n_833),
.Y(n_858)
);

OR2x6_ASAP7_75t_L g859 ( 
.A(n_794),
.B(n_484),
.Y(n_859)
);

AO22x1_ASAP7_75t_L g860 ( 
.A1(n_826),
.A2(n_356),
.B1(n_352),
.B2(n_350),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_804),
.Y(n_861)
);

O2A1O1Ixp5_ASAP7_75t_L g862 ( 
.A1(n_829),
.A2(n_490),
.B(n_484),
.C(n_17),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_763),
.B(n_851),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_783),
.Y(n_864)
);

INVxp67_ASAP7_75t_SL g865 ( 
.A(n_775),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_789),
.A2(n_490),
.B(n_484),
.Y(n_866)
);

OAI21x1_ASAP7_75t_L g867 ( 
.A1(n_812),
.A2(n_116),
.B(n_221),
.Y(n_867)
);

OA21x2_ASAP7_75t_L g868 ( 
.A1(n_818),
.A2(n_345),
.B(n_490),
.Y(n_868)
);

OAI22xp33_ASAP7_75t_L g869 ( 
.A1(n_764),
.A2(n_490),
.B1(n_16),
.B2(n_17),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_786),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_772),
.A2(n_490),
.B(n_115),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_850),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_796),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_827),
.Y(n_874)
);

OR2x6_ASAP7_75t_L g875 ( 
.A(n_848),
.B(n_490),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_819),
.A2(n_113),
.B(n_218),
.Y(n_876)
);

INVxp67_ASAP7_75t_SL g877 ( 
.A(n_775),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_803),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_SL g879 ( 
.A1(n_834),
.A2(n_105),
.B(n_217),
.C(n_215),
.Y(n_879)
);

OAI21x1_ASAP7_75t_L g880 ( 
.A1(n_780),
.A2(n_103),
.B(n_208),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_768),
.B(n_15),
.Y(n_881)
);

OAI21x1_ASAP7_75t_L g882 ( 
.A1(n_820),
.A2(n_102),
.B(n_205),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_813),
.Y(n_883)
);

NAND2x1p5_ASAP7_75t_L g884 ( 
.A(n_774),
.B(n_53),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_790),
.A2(n_118),
.B(n_203),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_845),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_791),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_SL g888 ( 
.A(n_764),
.B(n_21),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_791),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_773),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_890)
);

OR2x6_ASAP7_75t_L g891 ( 
.A(n_848),
.B(n_57),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_770),
.A2(n_126),
.B(n_201),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_SL g893 ( 
.A1(n_769),
.A2(n_119),
.B(n_198),
.C(n_195),
.Y(n_893)
);

OAI211xp5_ASAP7_75t_L g894 ( 
.A1(n_846),
.A2(n_22),
.B(n_25),
.C(n_26),
.Y(n_894)
);

AND2x6_ASAP7_75t_L g895 ( 
.A(n_848),
.B(n_59),
.Y(n_895)
);

AO21x2_ASAP7_75t_L g896 ( 
.A1(n_776),
.A2(n_788),
.B(n_807),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_793),
.A2(n_127),
.B(n_194),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_792),
.Y(n_898)
);

OA21x2_ASAP7_75t_L g899 ( 
.A1(n_809),
.A2(n_94),
.B(n_190),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_766),
.B(n_26),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_807),
.B(n_811),
.Y(n_901)
);

INVx4_ASAP7_75t_L g902 ( 
.A(n_827),
.Y(n_902)
);

BUFx2_ASAP7_75t_SL g903 ( 
.A(n_765),
.Y(n_903)
);

OAI21x1_ASAP7_75t_L g904 ( 
.A1(n_781),
.A2(n_129),
.B(n_188),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_844),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_833),
.Y(n_906)
);

AO31x2_ASAP7_75t_L g907 ( 
.A1(n_777),
.A2(n_30),
.A3(n_31),
.B(n_32),
.Y(n_907)
);

OAI21x1_ASAP7_75t_L g908 ( 
.A1(n_815),
.A2(n_131),
.B(n_187),
.Y(n_908)
);

INVx5_ASAP7_75t_L g909 ( 
.A(n_825),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_792),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_828),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_846),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_792),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_821),
.Y(n_914)
);

OAI22xp33_ASAP7_75t_L g915 ( 
.A1(n_767),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_784),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_843),
.B(n_138),
.Y(n_917)
);

AO21x1_ASAP7_75t_SL g918 ( 
.A1(n_824),
.A2(n_38),
.B(n_41),
.Y(n_918)
);

OAI21x1_ASAP7_75t_L g919 ( 
.A1(n_808),
.A2(n_144),
.B(n_186),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_816),
.B(n_42),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_771),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_824),
.Y(n_922)
);

INVx5_ASAP7_75t_L g923 ( 
.A(n_841),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_855),
.B(n_44),
.Y(n_924)
);

OAI21x1_ASAP7_75t_L g925 ( 
.A1(n_802),
.A2(n_147),
.B(n_185),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_797),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_798),
.Y(n_927)
);

OAI21x1_ASAP7_75t_L g928 ( 
.A1(n_814),
.A2(n_137),
.B(n_184),
.Y(n_928)
);

OAI21x1_ASAP7_75t_L g929 ( 
.A1(n_814),
.A2(n_132),
.B(n_181),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_810),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_778),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_931)
);

OAI21x1_ASAP7_75t_L g932 ( 
.A1(n_799),
.A2(n_93),
.B(n_180),
.Y(n_932)
);

OAI21x1_ASAP7_75t_L g933 ( 
.A1(n_805),
.A2(n_83),
.B(n_179),
.Y(n_933)
);

OR2x6_ASAP7_75t_L g934 ( 
.A(n_785),
.B(n_800),
.Y(n_934)
);

AOI21xp33_ASAP7_75t_SL g935 ( 
.A1(n_832),
.A2(n_45),
.B(n_46),
.Y(n_935)
);

OA21x2_ASAP7_75t_L g936 ( 
.A1(n_793),
.A2(n_149),
.B(n_175),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_831),
.B(n_219),
.Y(n_937)
);

INVxp67_ASAP7_75t_SL g938 ( 
.A(n_855),
.Y(n_938)
);

OAI21x1_ASAP7_75t_L g939 ( 
.A1(n_806),
.A2(n_78),
.B(n_170),
.Y(n_939)
);

AO21x2_ASAP7_75t_L g940 ( 
.A1(n_852),
.A2(n_77),
.B(n_169),
.Y(n_940)
);

OAI21x1_ASAP7_75t_L g941 ( 
.A1(n_801),
.A2(n_75),
.B(n_168),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_823),
.A2(n_74),
.B(n_167),
.Y(n_942)
);

OAI21x1_ASAP7_75t_L g943 ( 
.A1(n_836),
.A2(n_73),
.B(n_163),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_831),
.A2(n_47),
.B(n_49),
.C(n_60),
.Y(n_944)
);

OAI21x1_ASAP7_75t_L g945 ( 
.A1(n_817),
.A2(n_800),
.B(n_777),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_782),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_853),
.A2(n_61),
.B(n_63),
.C(n_64),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_785),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_822),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_838),
.A2(n_830),
.B(n_840),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_830),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_842),
.A2(n_65),
.B(n_66),
.C(n_69),
.Y(n_952)
);

AOI21x1_ASAP7_75t_L g953 ( 
.A1(n_835),
.A2(n_171),
.B(n_150),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_795),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_837),
.B(n_72),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_795),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_854),
.Y(n_957)
);

INVxp67_ASAP7_75t_SL g958 ( 
.A(n_767),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_849),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_854),
.Y(n_960)
);

AO21x2_ASAP7_75t_L g961 ( 
.A1(n_839),
.A2(n_151),
.B(n_153),
.Y(n_961)
);

NAND2x1p5_ASAP7_75t_L g962 ( 
.A(n_847),
.B(n_154),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_957),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_927),
.B(n_854),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_960),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_959),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_954),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_917),
.B(n_849),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_922),
.A2(n_849),
.B(n_156),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_911),
.B(n_901),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_956),
.Y(n_971)
);

OR2x6_ASAP7_75t_L g972 ( 
.A(n_934),
.B(n_155),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_858),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_898),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_896),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_880),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_910),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_896),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_913),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_864),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_948),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_873),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_878),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_883),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_858),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_877),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_863),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_868),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_877),
.Y(n_989)
);

BUFx12f_ASAP7_75t_L g990 ( 
.A(n_872),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_856),
.A2(n_161),
.B(n_876),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_868),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_865),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_938),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_909),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_901),
.B(n_926),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_874),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_889),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_904),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_930),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_945),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_949),
.B(n_914),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_936),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_936),
.Y(n_1004)
);

AO21x1_ASAP7_75t_L g1005 ( 
.A1(n_944),
.A2(n_871),
.B(n_897),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_907),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_887),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_899),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_899),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_909),
.Y(n_1010)
);

AO21x2_ASAP7_75t_L g1011 ( 
.A1(n_871),
.A2(n_950),
.B(n_866),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_909),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_862),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_903),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_907),
.Y(n_1015)
);

AOI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_920),
.A2(n_944),
.B(n_881),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_937),
.B(n_924),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_909),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_923),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_907),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_870),
.Y(n_1021)
);

OR2x2_ASAP7_75t_L g1022 ( 
.A(n_924),
.B(n_951),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_870),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_862),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_917),
.Y(n_1025)
);

INVxp67_ASAP7_75t_R g1026 ( 
.A(n_928),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_906),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_919),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_861),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_946),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_867),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_942),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_SL g1033 ( 
.A1(n_888),
.A2(n_923),
.B1(n_937),
.B2(n_894),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_918),
.B(n_949),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_908),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_929),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_948),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_948),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_934),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_882),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_934),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_892),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_943),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_892),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_958),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_906),
.Y(n_1046)
);

INVx6_ASAP7_75t_L g1047 ( 
.A(n_906),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_900),
.B(n_958),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_933),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_923),
.B(n_900),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_R g1051 ( 
.A(n_990),
.B(n_857),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_985),
.B(n_902),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_963),
.Y(n_1053)
);

NAND2xp33_ASAP7_75t_R g1054 ( 
.A(n_1034),
.B(n_891),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_985),
.B(n_902),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_985),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_987),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_996),
.B(n_923),
.Y(n_1058)
);

NAND2xp33_ASAP7_75t_R g1059 ( 
.A(n_1034),
.B(n_891),
.Y(n_1059)
);

OR2x6_ASAP7_75t_L g1060 ( 
.A(n_972),
.B(n_891),
.Y(n_1060)
);

XNOR2xp5_ASAP7_75t_L g1061 ( 
.A(n_1014),
.B(n_860),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_1046),
.B(n_857),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_1046),
.B(n_973),
.Y(n_1063)
);

OR2x6_ASAP7_75t_L g1064 ( 
.A(n_972),
.B(n_884),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_1046),
.B(n_857),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_963),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_R g1067 ( 
.A(n_990),
.B(n_888),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_R g1068 ( 
.A(n_973),
.B(n_895),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_996),
.B(n_890),
.Y(n_1069)
);

INVxp67_ASAP7_75t_L g1070 ( 
.A(n_997),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_972),
.B(n_1039),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_970),
.B(n_1048),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_1016),
.B(n_884),
.Y(n_1073)
);

INVxp67_ASAP7_75t_L g1074 ( 
.A(n_998),
.Y(n_1074)
);

BUFx10_ASAP7_75t_L g1075 ( 
.A(n_1047),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1048),
.B(n_890),
.Y(n_1076)
);

NAND2xp33_ASAP7_75t_R g1077 ( 
.A(n_1050),
.B(n_935),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_965),
.Y(n_1078)
);

NAND2xp33_ASAP7_75t_R g1079 ( 
.A(n_972),
.B(n_955),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_1027),
.B(n_859),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_R g1081 ( 
.A(n_1047),
.B(n_895),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_R g1082 ( 
.A(n_1047),
.B(n_895),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_1045),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1002),
.B(n_912),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_972),
.B(n_859),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_980),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_R g1087 ( 
.A(n_1047),
.B(n_895),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_980),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1022),
.B(n_894),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_981),
.Y(n_1090)
);

OR2x6_ASAP7_75t_L g1091 ( 
.A(n_995),
.B(n_875),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_R g1092 ( 
.A(n_1037),
.B(n_953),
.Y(n_1092)
);

NAND2xp33_ASAP7_75t_R g1093 ( 
.A(n_1017),
.B(n_875),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_1007),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_1039),
.B(n_859),
.Y(n_1095)
);

OR2x6_ASAP7_75t_L g1096 ( 
.A(n_995),
.B(n_1010),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1022),
.B(n_886),
.Y(n_1097)
);

NOR2x1_ASAP7_75t_L g1098 ( 
.A(n_993),
.B(n_905),
.Y(n_1098)
);

OR2x6_ASAP7_75t_L g1099 ( 
.A(n_1010),
.B(n_875),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_965),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_1041),
.Y(n_1101)
);

NAND2xp33_ASAP7_75t_SL g1102 ( 
.A(n_993),
.B(n_916),
.Y(n_1102)
);

CKINVDCx8_ASAP7_75t_R g1103 ( 
.A(n_981),
.Y(n_1103)
);

CKINVDCx8_ASAP7_75t_R g1104 ( 
.A(n_981),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1030),
.Y(n_1105)
);

OR2x2_ASAP7_75t_L g1106 ( 
.A(n_994),
.B(n_962),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_1037),
.B(n_940),
.Y(n_1107)
);

CKINVDCx8_ASAP7_75t_R g1108 ( 
.A(n_981),
.Y(n_1108)
);

CKINVDCx8_ASAP7_75t_R g1109 ( 
.A(n_981),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1017),
.B(n_931),
.Y(n_1110)
);

NAND2xp33_ASAP7_75t_R g1111 ( 
.A(n_968),
.B(n_897),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_1033),
.B(n_1025),
.Y(n_1112)
);

NAND2xp33_ASAP7_75t_R g1113 ( 
.A(n_968),
.B(n_885),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_R g1114 ( 
.A(n_1038),
.B(n_921),
.Y(n_1114)
);

OR2x4_ASAP7_75t_L g1115 ( 
.A(n_981),
.B(n_915),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_1038),
.B(n_962),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1102),
.A2(n_1005),
.B1(n_869),
.B2(n_1011),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1053),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1072),
.B(n_986),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1066),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1078),
.B(n_975),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1100),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1105),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1086),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1088),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1071),
.B(n_1001),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1083),
.B(n_986),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1101),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1101),
.B(n_975),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_1098),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1107),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1058),
.B(n_975),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_1094),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1106),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1071),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1076),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1110),
.B(n_978),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1096),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1069),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1096),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1089),
.B(n_978),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1095),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1060),
.B(n_978),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_1114),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1060),
.B(n_1006),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1095),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1090),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1074),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1091),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1073),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1112),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1064),
.B(n_1006),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1064),
.B(n_1015),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1057),
.B(n_1015),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1091),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1070),
.B(n_1020),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1097),
.B(n_989),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1085),
.B(n_1020),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1099),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1092),
.B(n_988),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1099),
.B(n_988),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1063),
.B(n_988),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1052),
.B(n_1001),
.Y(n_1163)
);

CKINVDCx14_ASAP7_75t_R g1164 ( 
.A(n_1067),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1103),
.B(n_992),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1115),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1104),
.B(n_992),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1108),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1128),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_1128),
.B(n_1001),
.Y(n_1170)
);

OAI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1166),
.A2(n_1079),
.B1(n_1059),
.B2(n_1054),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1136),
.B(n_989),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1118),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1118),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1118),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1136),
.B(n_964),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1132),
.B(n_1003),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1118),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1128),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1120),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1132),
.B(n_1003),
.Y(n_1181)
);

NOR2x1_ASAP7_75t_SL g1182 ( 
.A(n_1144),
.B(n_1011),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1120),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1120),
.Y(n_1184)
);

NAND2x1_ASAP7_75t_L g1185 ( 
.A(n_1144),
.B(n_994),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1128),
.B(n_1011),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_1130),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1154),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1120),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1154),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1132),
.B(n_1003),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1141),
.B(n_1004),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1138),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1124),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1122),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1139),
.B(n_964),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1124),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1154),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1156),
.Y(n_1199)
);

AOI211xp5_ASAP7_75t_L g1200 ( 
.A1(n_1130),
.A2(n_1005),
.B(n_1061),
.C(n_905),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1124),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1141),
.B(n_1004),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1141),
.B(n_1004),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1166),
.A2(n_1061),
.B1(n_1084),
.B2(n_1025),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1137),
.B(n_992),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1122),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1123),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1125),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1123),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1139),
.B(n_974),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1157),
.B(n_974),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1125),
.Y(n_1212)
);

INVx4_ASAP7_75t_L g1213 ( 
.A(n_1144),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1125),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1137),
.B(n_1008),
.Y(n_1215)
);

INVxp67_ASAP7_75t_SL g1216 ( 
.A(n_1127),
.Y(n_1216)
);

INVxp67_ASAP7_75t_SL g1217 ( 
.A(n_1127),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1121),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1134),
.B(n_1042),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1121),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1137),
.B(n_1008),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1126),
.B(n_1008),
.Y(n_1222)
);

AND2x2_ASAP7_75t_L g1223 ( 
.A(n_1126),
.B(n_1009),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1126),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1218),
.B(n_1134),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1195),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1187),
.Y(n_1227)
);

OR2x2_ASAP7_75t_L g1228 ( 
.A(n_1218),
.B(n_1156),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1173),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_1216),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1171),
.B(n_1151),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1195),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1224),
.B(n_1188),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1224),
.B(n_1146),
.Y(n_1234)
);

INVx3_ASAP7_75t_L g1235 ( 
.A(n_1224),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1174),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1216),
.B(n_1133),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1174),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1224),
.B(n_1188),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1190),
.B(n_1198),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1173),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1206),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1213),
.B(n_1164),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1175),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1206),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1190),
.B(n_1146),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1207),
.Y(n_1247)
);

NAND3xp33_ASAP7_75t_L g1248 ( 
.A(n_1200),
.B(n_1117),
.C(n_1150),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1199),
.B(n_1146),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1213),
.B(n_1164),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1218),
.B(n_1156),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_1220),
.B(n_1133),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1175),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1207),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1217),
.B(n_1150),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1220),
.B(n_1129),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1177),
.B(n_1146),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1226),
.Y(n_1258)
);

AO221x2_ASAP7_75t_L g1259 ( 
.A1(n_1248),
.A2(n_1148),
.B1(n_1151),
.B2(n_1155),
.C(n_1168),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1237),
.B(n_1217),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1255),
.B(n_1187),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1230),
.B(n_1148),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1227),
.B(n_1192),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1252),
.B(n_1192),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1231),
.A2(n_1200),
.B1(n_1077),
.B2(n_1166),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1243),
.B(n_1213),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1252),
.B(n_1192),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1257),
.B(n_1202),
.Y(n_1268)
);

NAND2xp33_ASAP7_75t_SL g1269 ( 
.A(n_1240),
.B(n_1051),
.Y(n_1269)
);

NAND2xp33_ASAP7_75t_SL g1270 ( 
.A(n_1240),
.B(n_1068),
.Y(n_1270)
);

NAND2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1249),
.B(n_1081),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1257),
.B(n_1177),
.Y(n_1272)
);

AO221x2_ASAP7_75t_L g1273 ( 
.A1(n_1232),
.A2(n_1155),
.B1(n_1168),
.B2(n_1138),
.C(n_1140),
.Y(n_1273)
);

NOR4xp25_ASAP7_75t_SL g1274 ( 
.A(n_1242),
.B(n_1093),
.C(n_1111),
.D(n_1113),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1249),
.B(n_1246),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1246),
.B(n_1202),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1245),
.B(n_1202),
.Y(n_1277)
);

INVxp67_ASAP7_75t_L g1278 ( 
.A(n_1250),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1247),
.Y(n_1279)
);

AO221x2_ASAP7_75t_L g1280 ( 
.A1(n_1254),
.A2(n_1168),
.B1(n_1140),
.B2(n_1138),
.C(n_1135),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1256),
.B(n_1177),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1235),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_R g1283 ( 
.A(n_1235),
.B(n_1056),
.Y(n_1283)
);

OAI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1256),
.A2(n_1213),
.B1(n_1185),
.B2(n_1149),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1225),
.B(n_1203),
.Y(n_1285)
);

AO221x2_ASAP7_75t_L g1286 ( 
.A1(n_1236),
.A2(n_1168),
.B1(n_1140),
.B2(n_1138),
.C(n_1135),
.Y(n_1286)
);

AO221x2_ASAP7_75t_L g1287 ( 
.A1(n_1236),
.A2(n_1140),
.B1(n_1149),
.B2(n_1159),
.C(n_969),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1234),
.B(n_1159),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1225),
.B(n_1203),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1269),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1258),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1279),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1288),
.B(n_1235),
.Y(n_1293)
);

INVx1_ASAP7_75t_SL g1294 ( 
.A(n_1283),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1277),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_1270),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_1286),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1265),
.B(n_1259),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1259),
.B(n_1234),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1261),
.B(n_1204),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1278),
.A2(n_1117),
.B1(n_1185),
.B2(n_1159),
.Y(n_1301)
);

INVx3_ASAP7_75t_L g1302 ( 
.A(n_1282),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1262),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1260),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1273),
.B(n_1233),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1263),
.A2(n_1241),
.B(n_1229),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1281),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1264),
.B(n_1228),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1273),
.B(n_1233),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1286),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1274),
.A2(n_1149),
.B1(n_1142),
.B2(n_1157),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1266),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1271),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1280),
.B(n_1239),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1267),
.B(n_1228),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1285),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1289),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1275),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_1268),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1280),
.B(n_1239),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1272),
.B(n_1182),
.Y(n_1321)
);

NAND3xp33_ASAP7_75t_L g1322 ( 
.A(n_1287),
.B(n_1145),
.C(n_1147),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1276),
.B(n_1062),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1298),
.A2(n_1287),
.B(n_1284),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1313),
.B(n_1251),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1300),
.A2(n_1182),
.B(n_1172),
.Y(n_1326)
);

NOR2xp67_ASAP7_75t_L g1327 ( 
.A(n_1297),
.B(n_1241),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1291),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1292),
.B(n_1193),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1292),
.B(n_1193),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1302),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1318),
.B(n_1251),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1290),
.B(n_1065),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1303),
.B(n_1193),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_SL g1335 ( 
.A1(n_1294),
.A2(n_1019),
.B(n_1087),
.C(n_1082),
.Y(n_1335)
);

OAI321xp33_ASAP7_75t_L g1336 ( 
.A1(n_1313),
.A2(n_1301),
.A3(n_1322),
.B1(n_1311),
.B2(n_1304),
.C(n_1310),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1304),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1319),
.B(n_1238),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1312),
.B(n_1238),
.Y(n_1339)
);

OAI32xp33_ASAP7_75t_L g1340 ( 
.A1(n_1310),
.A2(n_1196),
.A3(n_1176),
.B1(n_1186),
.B2(n_1244),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1312),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1296),
.B(n_1244),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1302),
.B(n_1293),
.Y(n_1343)
);

OAI221xp5_ASAP7_75t_L g1344 ( 
.A1(n_1299),
.A2(n_1142),
.B1(n_1196),
.B2(n_1176),
.C(n_1253),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1309),
.A2(n_1149),
.B1(n_1186),
.B2(n_1131),
.Y(n_1345)
);

AND2x4_ASAP7_75t_SL g1346 ( 
.A(n_1302),
.B(n_1075),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1307),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1305),
.A2(n_1145),
.B1(n_1116),
.B2(n_1160),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1320),
.A2(n_952),
.B(n_947),
.Y(n_1349)
);

AOI222xp33_ASAP7_75t_L g1350 ( 
.A1(n_1305),
.A2(n_1145),
.B1(n_1152),
.B2(n_1153),
.C1(n_1203),
.C2(n_1211),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1317),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1293),
.B(n_1181),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1295),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1295),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1314),
.B(n_1172),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1341),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1347),
.B(n_1316),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1328),
.Y(n_1358)
);

NOR2x1p5_ASAP7_75t_SL g1359 ( 
.A(n_1353),
.B(n_1316),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1333),
.B(n_1323),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1336),
.B(n_1348),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1354),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1331),
.B(n_1314),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1337),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1351),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1339),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1333),
.B(n_1308),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1343),
.B(n_1325),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1324),
.B(n_1308),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1342),
.B(n_1315),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1338),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1332),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1329),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1346),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1348),
.A2(n_1315),
.B1(n_1321),
.B2(n_1131),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1330),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1346),
.B(n_1321),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1344),
.B(n_1306),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1349),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1355),
.A2(n_1152),
.B1(n_1153),
.B2(n_1158),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1334),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1355),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1350),
.B(n_1306),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1352),
.Y(n_1384)
);

NOR2xp67_ASAP7_75t_L g1385 ( 
.A(n_1327),
.B(n_1241),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1345),
.B(n_1253),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1362),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1364),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1372),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1357),
.Y(n_1390)
);

INVxp33_ASAP7_75t_L g1391 ( 
.A(n_1356),
.Y(n_1391)
);

INVx4_ASAP7_75t_L g1392 ( 
.A(n_1379),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1358),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1365),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1368),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1374),
.B(n_1335),
.Y(n_1396)
);

INVx1_ASAP7_75t_SL g1397 ( 
.A(n_1382),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1366),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1371),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1384),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1363),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1360),
.B(n_1335),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1373),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1376),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1381),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1370),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1359),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1367),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1367),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1369),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1386),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1385),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1377),
.Y(n_1413)
);

INVxp33_ASAP7_75t_SL g1414 ( 
.A(n_1360),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1377),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1380),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1361),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1383),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1375),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1378),
.Y(n_1420)
);

BUFx12f_ASAP7_75t_L g1421 ( 
.A(n_1378),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1356),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1356),
.B(n_1326),
.Y(n_1423)
);

INVxp67_ASAP7_75t_L g1424 ( 
.A(n_1356),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1414),
.B(n_1340),
.Y(n_1425)
);

O2A1O1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1410),
.A2(n_952),
.B(n_947),
.C(n_879),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1422),
.Y(n_1427)
);

AOI211xp5_ASAP7_75t_L g1428 ( 
.A1(n_1417),
.A2(n_893),
.B(n_1055),
.C(n_885),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1392),
.B(n_1229),
.Y(n_1429)
);

NAND3xp33_ASAP7_75t_SL g1430 ( 
.A(n_1410),
.B(n_1109),
.C(n_1160),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1392),
.B(n_1209),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1391),
.B(n_1209),
.Y(n_1432)
);

NOR2xp67_ASAP7_75t_L g1433 ( 
.A(n_1424),
.B(n_1407),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1422),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1397),
.B(n_1179),
.Y(n_1435)
);

OAI211xp5_ASAP7_75t_L g1436 ( 
.A1(n_1418),
.A2(n_1402),
.B(n_1396),
.C(n_1420),
.Y(n_1436)
);

NOR3xp33_ASAP7_75t_L g1437 ( 
.A(n_1424),
.B(n_1147),
.C(n_1080),
.Y(n_1437)
);

NOR2x1_ASAP7_75t_L g1438 ( 
.A(n_1408),
.B(n_1000),
.Y(n_1438)
);

NOR3x1_ASAP7_75t_L g1439 ( 
.A(n_1413),
.B(n_1179),
.C(n_1210),
.Y(n_1439)
);

NAND4xp75_ASAP7_75t_L g1440 ( 
.A(n_1396),
.B(n_1160),
.C(n_1153),
.D(n_1152),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1395),
.B(n_1391),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1389),
.Y(n_1442)
);

NOR3x1_ASAP7_75t_L g1443 ( 
.A(n_1415),
.B(n_1210),
.C(n_1000),
.Y(n_1443)
);

AOI221xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1419),
.A2(n_1402),
.B1(n_1411),
.B2(n_1416),
.C(n_1423),
.Y(n_1444)
);

NAND5xp2_ASAP7_75t_L g1445 ( 
.A(n_1409),
.B(n_1030),
.C(n_1041),
.D(n_1042),
.E(n_1044),
.Y(n_1445)
);

O2A1O1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1399),
.A2(n_961),
.B(n_1012),
.C(n_1018),
.Y(n_1446)
);

NAND4xp25_ASAP7_75t_L g1447 ( 
.A(n_1406),
.B(n_1400),
.C(n_1401),
.D(n_1390),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1421),
.B(n_1219),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1387),
.Y(n_1449)
);

NAND4xp25_ASAP7_75t_L g1450 ( 
.A(n_1400),
.B(n_1158),
.C(n_1211),
.D(n_1143),
.Y(n_1450)
);

NOR3x1_ASAP7_75t_L g1451 ( 
.A(n_1405),
.B(n_1119),
.C(n_1219),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_SL g1452 ( 
.A(n_1401),
.B(n_1412),
.Y(n_1452)
);

A2O1A1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1403),
.A2(n_1212),
.B(n_1143),
.C(n_1158),
.Y(n_1453)
);

NOR3x1_ASAP7_75t_SL g1454 ( 
.A(n_1403),
.B(n_1398),
.C(n_1404),
.Y(n_1454)
);

AND5x1_ASAP7_75t_L g1455 ( 
.A(n_1393),
.B(n_866),
.C(n_1026),
.D(n_1143),
.E(n_1163),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1394),
.B(n_1212),
.Y(n_1456)
);

OAI211xp5_ASAP7_75t_SL g1457 ( 
.A1(n_1436),
.A2(n_1388),
.B(n_1029),
.C(n_950),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1425),
.A2(n_1181),
.B1(n_1191),
.B2(n_1161),
.Y(n_1458)
);

AND4x1_ASAP7_75t_L g1459 ( 
.A(n_1441),
.B(n_1165),
.C(n_1167),
.D(n_1029),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1427),
.Y(n_1460)
);

NOR4xp25_ASAP7_75t_L g1461 ( 
.A(n_1454),
.B(n_983),
.C(n_982),
.D(n_984),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1434),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1444),
.A2(n_1430),
.B1(n_1440),
.B2(n_1437),
.Y(n_1463)
);

OAI31xp33_ASAP7_75t_L g1464 ( 
.A1(n_1447),
.A2(n_1044),
.A3(n_1169),
.B(n_968),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1433),
.A2(n_1191),
.B1(n_1181),
.B2(n_1161),
.Y(n_1465)
);

O2A1O1Ixp33_ASAP7_75t_SL g1466 ( 
.A1(n_1452),
.A2(n_1169),
.B(n_1023),
.C(n_982),
.Y(n_1466)
);

NOR4xp25_ASAP7_75t_L g1467 ( 
.A(n_1442),
.B(n_983),
.C(n_984),
.D(n_1180),
.Y(n_1467)
);

INVxp67_ASAP7_75t_L g1468 ( 
.A(n_1429),
.Y(n_1468)
);

AOI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1448),
.A2(n_1184),
.B1(n_1180),
.B2(n_1119),
.C(n_1208),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1435),
.A2(n_1024),
.B1(n_1013),
.B2(n_968),
.Y(n_1470)
);

AOI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1449),
.A2(n_1184),
.B1(n_1214),
.B2(n_1208),
.C(n_1201),
.Y(n_1471)
);

NOR3xp33_ASAP7_75t_L g1472 ( 
.A(n_1431),
.B(n_939),
.C(n_925),
.Y(n_1472)
);

OAI211xp5_ASAP7_75t_L g1473 ( 
.A1(n_1432),
.A2(n_1023),
.B(n_1214),
.C(n_1201),
.Y(n_1473)
);

AOI32xp33_ASAP7_75t_L g1474 ( 
.A1(n_1438),
.A2(n_1165),
.A3(n_1167),
.B1(n_1191),
.B2(n_1161),
.Y(n_1474)
);

NAND4xp25_ASAP7_75t_SL g1475 ( 
.A(n_1446),
.B(n_1167),
.C(n_1165),
.D(n_1223),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1443),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1450),
.A2(n_1163),
.B1(n_1126),
.B2(n_940),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1453),
.A2(n_1178),
.B1(n_1183),
.B2(n_1189),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1456),
.A2(n_1126),
.B1(n_1163),
.B2(n_1222),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_SL g1480 ( 
.A(n_1428),
.B(n_1021),
.C(n_1045),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1439),
.A2(n_1194),
.B1(n_1208),
.B2(n_1201),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1445),
.A2(n_1163),
.B1(n_961),
.B2(n_1162),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1451),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1445),
.Y(n_1484)
);

AOI211xp5_ASAP7_75t_SL g1485 ( 
.A1(n_1455),
.A2(n_1032),
.B(n_1028),
.C(n_1170),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1426),
.A2(n_1163),
.B1(n_1162),
.B2(n_1013),
.Y(n_1486)
);

AOI221xp5_ASAP7_75t_L g1487 ( 
.A1(n_1425),
.A2(n_1194),
.B1(n_1197),
.B2(n_1214),
.C(n_1173),
.Y(n_1487)
);

NOR3xp33_ASAP7_75t_L g1488 ( 
.A(n_1436),
.B(n_932),
.C(n_1032),
.Y(n_1488)
);

NAND4xp25_ASAP7_75t_L g1489 ( 
.A(n_1444),
.B(n_1036),
.C(n_1028),
.D(n_1162),
.Y(n_1489)
);

AOI221xp5_ASAP7_75t_L g1490 ( 
.A1(n_1425),
.A2(n_1197),
.B1(n_1194),
.B2(n_1178),
.C(n_1183),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1461),
.A2(n_1036),
.B(n_1021),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1460),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1463),
.B(n_1197),
.Y(n_1493)
);

XNOR2xp5_ASAP7_75t_L g1494 ( 
.A(n_1483),
.B(n_1223),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1462),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1476),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1468),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1459),
.B(n_1189),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1484),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1480),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1475),
.A2(n_1223),
.B1(n_1222),
.B2(n_1189),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1489),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1457),
.A2(n_1222),
.B1(n_1178),
.B2(n_1183),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1488),
.B(n_1205),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1458),
.B(n_1170),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1467),
.B(n_1205),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1485),
.B(n_1464),
.Y(n_1507)
);

NOR2xp67_ASAP7_75t_L g1508 ( 
.A(n_1473),
.B(n_1049),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1466),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1465),
.Y(n_1510)
);

NAND4xp75_ASAP7_75t_L g1511 ( 
.A(n_1487),
.B(n_1490),
.C(n_1469),
.D(n_1471),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1481),
.B(n_1205),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1496),
.B(n_1474),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_R g1514 ( 
.A(n_1497),
.B(n_1477),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_R g1515 ( 
.A(n_1499),
.B(n_1482),
.Y(n_1515)
);

NOR3xp33_ASAP7_75t_SL g1516 ( 
.A(n_1493),
.B(n_1470),
.C(n_1478),
.Y(n_1516)
);

NAND2xp33_ASAP7_75t_SL g1517 ( 
.A(n_1509),
.B(n_1470),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1510),
.B(n_1486),
.Y(n_1518)
);

NAND2xp33_ASAP7_75t_SL g1519 ( 
.A(n_1509),
.B(n_1479),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_R g1520 ( 
.A(n_1492),
.B(n_1495),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_R g1521 ( 
.A(n_1500),
.B(n_999),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_R g1522 ( 
.A(n_1494),
.B(n_999),
.Y(n_1522)
);

NOR3xp33_ASAP7_75t_SL g1523 ( 
.A(n_1507),
.B(n_1511),
.C(n_1504),
.Y(n_1523)
);

NAND2xp33_ASAP7_75t_SL g1524 ( 
.A(n_1498),
.B(n_1221),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_R g1525 ( 
.A(n_1502),
.B(n_999),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1498),
.B(n_1472),
.Y(n_1526)
);

NOR3xp33_ASAP7_75t_SL g1527 ( 
.A(n_1491),
.B(n_1049),
.C(n_966),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_R g1528 ( 
.A(n_1506),
.B(n_999),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1503),
.B(n_1013),
.C(n_1024),
.Y(n_1529)
);

XNOR2xp5_ASAP7_75t_L g1530 ( 
.A(n_1508),
.B(n_991),
.Y(n_1530)
);

OAI211xp5_ASAP7_75t_L g1531 ( 
.A1(n_1520),
.A2(n_1512),
.B(n_1505),
.C(n_1501),
.Y(n_1531)
);

NAND2xp33_ASAP7_75t_SL g1532 ( 
.A(n_1521),
.B(n_1221),
.Y(n_1532)
);

XNOR2x1_ASAP7_75t_L g1533 ( 
.A(n_1513),
.B(n_941),
.Y(n_1533)
);

NAND2x1_ASAP7_75t_L g1534 ( 
.A(n_1516),
.B(n_1221),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1518),
.A2(n_1215),
.B1(n_1129),
.B2(n_1024),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1514),
.Y(n_1536)
);

AND4x1_ASAP7_75t_L g1537 ( 
.A(n_1523),
.B(n_1215),
.C(n_1129),
.D(n_1121),
.Y(n_1537)
);

INVxp33_ASAP7_75t_SL g1538 ( 
.A(n_1525),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1519),
.A2(n_1215),
.B1(n_1026),
.B2(n_976),
.Y(n_1539)
);

NOR3xp33_ASAP7_75t_L g1540 ( 
.A(n_1517),
.B(n_991),
.C(n_976),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1526),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1515),
.B(n_966),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1538),
.B(n_1524),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1534),
.Y(n_1544)
);

XNOR2xp5_ASAP7_75t_L g1545 ( 
.A(n_1537),
.B(n_1530),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1536),
.B(n_1527),
.Y(n_1546)
);

XOR2x2_ASAP7_75t_L g1547 ( 
.A(n_1541),
.B(n_1529),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1531),
.A2(n_1522),
.B1(n_1528),
.B2(n_1043),
.Y(n_1548)
);

XNOR2xp5_ASAP7_75t_L g1549 ( 
.A(n_1539),
.B(n_1043),
.Y(n_1549)
);

NAND2x1p5_ASAP7_75t_L g1550 ( 
.A(n_1542),
.B(n_976),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1532),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1533),
.B(n_977),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_SL g1553 ( 
.A1(n_1544),
.A2(n_1535),
.B1(n_1540),
.B2(n_976),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1551),
.Y(n_1554)
);

NOR2xp67_ASAP7_75t_L g1555 ( 
.A(n_1548),
.B(n_1035),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1547),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1545),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1554),
.A2(n_1543),
.B1(n_1552),
.B2(n_1546),
.Y(n_1558)
);

AOI31xp33_ASAP7_75t_L g1559 ( 
.A1(n_1556),
.A2(n_1550),
.A3(n_1549),
.B(n_1031),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1559),
.Y(n_1560)
);

XOR2xp5_ASAP7_75t_L g1561 ( 
.A(n_1558),
.B(n_1557),
.Y(n_1561)
);

OAI222xp33_ASAP7_75t_L g1562 ( 
.A1(n_1561),
.A2(n_1553),
.B1(n_1555),
.B2(n_1043),
.C1(n_1031),
.C2(n_1035),
.Y(n_1562)
);

AOI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1560),
.A2(n_1040),
.B1(n_979),
.B2(n_977),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1563),
.Y(n_1564)
);

OAI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1562),
.A2(n_1040),
.B(n_979),
.Y(n_1565)
);

OAI221xp5_ASAP7_75t_R g1566 ( 
.A1(n_1564),
.A2(n_1040),
.B1(n_1009),
.B2(n_971),
.C(n_967),
.Y(n_1566)
);

AOI211xp5_ASAP7_75t_L g1567 ( 
.A1(n_1566),
.A2(n_1565),
.B(n_967),
.C(n_971),
.Y(n_1567)
);


endmodule