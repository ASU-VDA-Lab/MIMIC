module fake_jpeg_27116_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx11_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_14),
.Y(n_17)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_20),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_11),
.B(n_0),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_21),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_10),
.B1(n_27),
.B2(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_33),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_14),
.C(n_20),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_18),
.Y(n_33)
);

NAND2x1_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_17),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_27),
.B1(n_17),
.B2(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_14),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_12),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_39),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_26),
.B1(n_8),
.B2(n_16),
.Y(n_43)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_35),
.B1(n_34),
.B2(n_16),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_44),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_19),
.C(n_22),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_41),
.C(n_22),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_47),
.C(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_39),
.B1(n_38),
.B2(n_15),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_38),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_52),
.B(n_3),
.Y(n_53)
);

AO21x1_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_5),
.B(n_6),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_7),
.Y(n_55)
);


endmodule