module fake_jpeg_13324_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

BUFx3_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_2),
.B(n_4),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

OR2x2_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_2),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_8),
.B(n_2),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_18),
.B(n_19),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_7),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_20),
.A2(n_22),
.B1(n_6),
.B2(n_11),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_22),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_17),
.A2(n_1),
.B1(n_9),
.B2(n_20),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_17),
.B1(n_14),
.B2(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_22),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_32),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_30),
.B1(n_25),
.B2(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_33),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_37),
.B(n_32),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_39),
.A2(n_37),
.B(n_29),
.Y(n_40)
);


endmodule