module fake_netlist_1_11241_n_854 (n_117, n_44, n_133, n_149, n_81, n_69, n_204, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_96, n_39, n_854);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_204;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_96;
input n_39;
output n_854;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_383;
wire n_288;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_809;
wire n_580;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_769;
wire n_844;
wire n_230;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_771;
wire n_735;
wire n_696;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_357;
wire n_245;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_406;
wire n_395;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_209), .Y(n_212) );
INVx1_ASAP7_75t_SL g213 ( .A(n_13), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_149), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_51), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_30), .Y(n_216) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_126), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_175), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_168), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_152), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_160), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_33), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_101), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_200), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_103), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_79), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_197), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_132), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_90), .Y(n_229) );
BUFx8_ASAP7_75t_SL g230 ( .A(n_193), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_48), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_115), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_153), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_38), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_42), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_86), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_166), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_190), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_107), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_56), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_169), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_14), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_11), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_140), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_183), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_189), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_74), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_167), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_192), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_60), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_118), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_96), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_25), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_110), .Y(n_254) );
INVxp67_ASAP7_75t_L g255 ( .A(n_6), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_176), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_13), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_180), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_62), .Y(n_259) );
INVx1_ASAP7_75t_SL g260 ( .A(n_71), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_95), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_143), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_2), .Y(n_263) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_72), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_162), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_151), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_111), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_164), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_0), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_64), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_21), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_181), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_146), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_45), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_16), .Y(n_275) );
BUFx3_ASAP7_75t_L g276 ( .A(n_26), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_39), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_100), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_102), .B(n_109), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_121), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_66), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_4), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_198), .Y(n_283) );
CKINVDCx16_ASAP7_75t_R g284 ( .A(n_9), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_23), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_194), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_105), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_117), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_196), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_182), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_55), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_43), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_123), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_83), .Y(n_294) );
INVxp33_ASAP7_75t_L g295 ( .A(n_24), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_58), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_32), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_92), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_211), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_170), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_163), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_4), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_177), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_36), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_70), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_63), .Y(n_306) );
CKINVDCx16_ASAP7_75t_R g307 ( .A(n_148), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_5), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_89), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_135), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_34), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_49), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_172), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_41), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_99), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_5), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_27), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_128), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_82), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_17), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_93), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_54), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_284), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_248), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_255), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_242), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_231), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_263), .A2(n_269), .B1(n_308), .B2(n_302), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_218), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_230), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_248), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_231), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_257), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_223), .Y(n_334) );
BUFx8_ASAP7_75t_L g335 ( .A(n_216), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_282), .B(n_1), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_255), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_231), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_307), .A2(n_3), .B1(n_6), .B2(n_7), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_316), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_236), .Y(n_341) );
INVx4_ASAP7_75t_L g342 ( .A(n_212), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_241), .B(n_3), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_247), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_231), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_295), .B(n_7), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_295), .B(n_8), .Y(n_347) );
INVx5_ASAP7_75t_L g348 ( .A(n_256), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g349 ( .A1(n_215), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_349) );
BUFx3_ASAP7_75t_L g350 ( .A(n_220), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_333), .Y(n_351) );
BUFx6f_ASAP7_75t_SL g352 ( .A(n_336), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_333), .Y(n_353) );
INVx4_ASAP7_75t_SL g354 ( .A(n_346), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_350), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_324), .B(n_271), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_348), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_336), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_348), .Y(n_359) );
NAND3xp33_ASAP7_75t_L g360 ( .A(n_324), .B(n_221), .C(n_219), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_327), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_343), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_342), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_342), .B(n_313), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_348), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_329), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_327), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_331), .B(n_275), .Y(n_368) );
OR2x6_ASAP7_75t_L g369 ( .A(n_337), .B(n_230), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_334), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_341), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_344), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_343), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_340), .B(n_313), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_326), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_327), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_328), .B(n_214), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_325), .A2(n_213), .B1(n_225), .B2(n_222), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_364), .B(n_347), .Y(n_379) );
NAND2xp33_ASAP7_75t_L g380 ( .A(n_362), .B(n_217), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_351), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_353), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_360), .A2(n_335), .B1(n_328), .B2(n_339), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_358), .B(n_335), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_366), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_362), .B(n_226), .Y(n_386) );
INVx8_ASAP7_75t_L g387 ( .A(n_352), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_370), .Y(n_388) );
A2O1A1Ixp33_ASAP7_75t_L g389 ( .A1(n_360), .A2(n_323), .B(n_235), .C(n_239), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_368), .B(n_224), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_368), .B(n_227), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_371), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_374), .B(n_229), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_372), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_356), .B(n_232), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_373), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_373), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_356), .B(n_234), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_363), .B(n_354), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_352), .A2(n_323), .B1(n_349), .B2(n_246), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_354), .B(n_326), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_357), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_355), .B(n_237), .Y(n_403) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_359), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_378), .B(n_238), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_375), .Y(n_406) );
NOR2xp67_ASAP7_75t_L g407 ( .A(n_377), .B(n_330), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_365), .Y(n_408) );
AOI21xp5_ASAP7_75t_L g409 ( .A1(n_379), .A2(n_240), .B(n_233), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_395), .B(n_228), .Y(n_410) );
AOI21xp5_ASAP7_75t_L g411 ( .A1(n_386), .A2(n_252), .B(n_244), .Y(n_411) );
NAND3xp33_ASAP7_75t_SL g412 ( .A(n_400), .B(n_264), .C(n_249), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_392), .Y(n_413) );
OAI21x1_ASAP7_75t_L g414 ( .A1(n_386), .A2(n_293), .B(n_277), .Y(n_414) );
O2A1O1Ixp5_ASAP7_75t_L g415 ( .A1(n_399), .A2(n_301), .B(n_310), .C(n_279), .Y(n_415) );
AOI21x1_ASAP7_75t_L g416 ( .A1(n_398), .A2(n_376), .B(n_261), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_394), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_396), .A2(n_267), .B(n_259), .Y(n_418) );
OAI21xp5_ASAP7_75t_L g419 ( .A1(n_385), .A2(n_270), .B(n_268), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_380), .A2(n_280), .B(n_273), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_404), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_390), .B(n_315), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_391), .B(n_369), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_397), .B(n_389), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_387), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_388), .B(n_369), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_382), .B(n_245), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_406), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_403), .A2(n_393), .B(n_381), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_405), .B(n_251), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g431 ( .A1(n_402), .A2(n_285), .B(n_281), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_401), .B(n_253), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_408), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_404), .Y(n_434) );
OAI21xp5_ASAP7_75t_L g435 ( .A1(n_401), .A2(n_290), .B(n_287), .Y(n_435) );
INVxp67_ASAP7_75t_SL g436 ( .A(n_404), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_384), .A2(n_300), .B(n_294), .Y(n_437) );
AOI21x1_ASAP7_75t_L g438 ( .A1(n_407), .A2(n_376), .B(n_303), .Y(n_438) );
OA22x2_ASAP7_75t_L g439 ( .A1(n_423), .A2(n_383), .B1(n_387), .B2(n_243), .Y(n_439) );
OAI21xp5_ASAP7_75t_L g440 ( .A1(n_429), .A2(n_312), .B(n_311), .Y(n_440) );
OAI21x1_ASAP7_75t_L g441 ( .A1(n_414), .A2(n_416), .B(n_438), .Y(n_441) );
AOI21x1_ASAP7_75t_L g442 ( .A1(n_411), .A2(n_320), .B(n_319), .Y(n_442) );
BUFx12f_ASAP7_75t_L g443 ( .A(n_425), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_424), .A2(n_387), .B(n_279), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_428), .Y(n_445) );
OAI21xp33_ASAP7_75t_L g446 ( .A1(n_422), .A2(n_296), .B(n_260), .Y(n_446) );
AND2x6_ASAP7_75t_L g447 ( .A(n_433), .B(n_250), .Y(n_447) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_421), .Y(n_448) );
OAI21x1_ASAP7_75t_L g449 ( .A1(n_421), .A2(n_434), .B(n_411), .Y(n_449) );
AO22x2_ASAP7_75t_L g450 ( .A1(n_412), .A2(n_276), .B1(n_254), .B2(n_12), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_409), .A2(n_262), .B(n_258), .Y(n_451) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_418), .A2(n_266), .B(n_265), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_413), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_410), .B(n_10), .Y(n_454) );
OA21x2_ASAP7_75t_L g455 ( .A1(n_419), .A2(n_274), .B(n_272), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_409), .B(n_278), .Y(n_456) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_434), .Y(n_457) );
OAI21x1_ASAP7_75t_L g458 ( .A1(n_415), .A2(n_291), .B(n_256), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_435), .A2(n_306), .B1(n_283), .B2(n_286), .Y(n_459) );
BUFx3_ASAP7_75t_L g460 ( .A(n_426), .Y(n_460) );
OR2x6_ASAP7_75t_L g461 ( .A(n_437), .B(n_256), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_437), .B(n_288), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_432), .Y(n_463) );
AO32x2_ASAP7_75t_L g464 ( .A1(n_420), .A2(n_345), .A3(n_332), .B1(n_338), .B2(n_15), .Y(n_464) );
NOR2x1_ASAP7_75t_SL g465 ( .A(n_417), .B(n_291), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_427), .A2(n_292), .B(n_289), .Y(n_466) );
OAI21x1_ASAP7_75t_L g467 ( .A1(n_436), .A2(n_291), .B(n_19), .Y(n_467) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_430), .A2(n_317), .B1(n_298), .B2(n_299), .C(n_304), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_431), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_425), .Y(n_470) );
INVx3_ASAP7_75t_L g471 ( .A(n_425), .Y(n_471) );
OR2x6_ASAP7_75t_L g472 ( .A(n_425), .B(n_11), .Y(n_472) );
INVx3_ASAP7_75t_L g473 ( .A(n_453), .Y(n_473) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_453), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_445), .B(n_12), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_460), .B(n_14), .Y(n_476) );
AO31x2_ASAP7_75t_L g477 ( .A1(n_465), .A2(n_345), .A3(n_338), .B(n_332), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_454), .B(n_15), .Y(n_478) );
AO32x2_ASAP7_75t_L g479 ( .A1(n_464), .A2(n_345), .A3(n_338), .B1(n_332), .B2(n_28), .Y(n_479) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_457), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_444), .A2(n_318), .B(n_305), .C(n_322), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_446), .B(n_297), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_469), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_472), .A2(n_321), .B1(n_314), .B2(n_309), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_469), .Y(n_485) );
OAI21x1_ASAP7_75t_L g486 ( .A1(n_441), .A2(n_18), .B(n_20), .Y(n_486) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_458), .A2(n_367), .B(n_361), .Y(n_487) );
OAI21x1_ASAP7_75t_L g488 ( .A1(n_449), .A2(n_22), .B(n_29), .Y(n_488) );
BUFx2_ASAP7_75t_L g489 ( .A(n_443), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_442), .Y(n_490) );
OAI21x1_ASAP7_75t_L g491 ( .A1(n_467), .A2(n_31), .B(n_35), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g492 ( .A1(n_440), .A2(n_37), .B(n_40), .C(n_44), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_470), .B(n_46), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_472), .B(n_439), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_450), .A2(n_367), .B1(n_361), .B2(n_52), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_452), .A2(n_47), .B(n_50), .C(n_53), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_471), .B(n_57), .Y(n_497) );
INVx4_ASAP7_75t_L g498 ( .A(n_447), .Y(n_498) );
INVx5_ASAP7_75t_L g499 ( .A(n_447), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_463), .B(n_59), .Y(n_500) );
INVx2_ASAP7_75t_SL g501 ( .A(n_447), .Y(n_501) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_456), .A2(n_61), .B(n_65), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_461), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_451), .A2(n_67), .B(n_68), .Y(n_504) );
BUFx2_ASAP7_75t_L g505 ( .A(n_455), .Y(n_505) );
OAI221xp5_ASAP7_75t_L g506 ( .A1(n_468), .A2(n_69), .B1(n_73), .B2(n_75), .C(n_76), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_459), .B(n_77), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_461), .Y(n_508) );
OAI21x1_ASAP7_75t_L g509 ( .A1(n_448), .A2(n_78), .B(n_80), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_455), .B(n_210), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_462), .A2(n_81), .B(n_84), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_457), .B(n_85), .Y(n_512) );
OAI21x1_ASAP7_75t_L g513 ( .A1(n_466), .A2(n_87), .B(n_88), .Y(n_513) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_441), .A2(n_91), .B(n_94), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_460), .B(n_97), .Y(n_515) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_441), .A2(n_98), .B(n_104), .Y(n_516) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_441), .A2(n_106), .B(n_108), .Y(n_517) );
BUFx2_ASAP7_75t_R g518 ( .A(n_460), .Y(n_518) );
OAI21x1_ASAP7_75t_L g519 ( .A1(n_441), .A2(n_112), .B(n_113), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_445), .B(n_114), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_445), .B(n_208), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_460), .B(n_116), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_445), .Y(n_523) );
BUFx3_ASAP7_75t_L g524 ( .A(n_443), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_440), .A2(n_119), .B(n_120), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_445), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_526), .Y(n_527) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_480), .Y(n_528) );
CKINVDCx11_ASAP7_75t_R g529 ( .A(n_524), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_490), .Y(n_530) );
INVx3_ASAP7_75t_L g531 ( .A(n_498), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_526), .Y(n_532) );
CKINVDCx6p67_ASAP7_75t_R g533 ( .A(n_489), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_523), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_520), .A2(n_122), .B(n_124), .C(n_125), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_475), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_474), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_494), .A2(n_127), .B1(n_129), .B2(n_130), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_498), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_473), .Y(n_540) );
INVx3_ASAP7_75t_L g541 ( .A(n_499), .Y(n_541) );
INVx2_ASAP7_75t_SL g542 ( .A(n_499), .Y(n_542) );
OAI21x1_ASAP7_75t_L g543 ( .A1(n_487), .A2(n_131), .B(n_133), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_473), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_476), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_476), .B(n_134), .Y(n_546) );
OAI21x1_ASAP7_75t_L g547 ( .A1(n_487), .A2(n_136), .B(n_137), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_483), .B(n_138), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_522), .B(n_207), .Y(n_549) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_483), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_485), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_520), .Y(n_552) );
OA21x2_ASAP7_75t_L g553 ( .A1(n_485), .A2(n_139), .B(n_141), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_499), .B(n_142), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_478), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_497), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_505), .B(n_144), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_525), .A2(n_145), .B(n_147), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_493), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_480), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_521), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_503), .Y(n_562) );
INVx3_ASAP7_75t_L g563 ( .A(n_501), .Y(n_563) );
BUFx3_ASAP7_75t_L g564 ( .A(n_512), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_503), .Y(n_565) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_508), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_515), .Y(n_567) );
NAND2xp33_ASAP7_75t_L g568 ( .A(n_507), .B(n_150), .Y(n_568) );
BUFx3_ASAP7_75t_L g569 ( .A(n_512), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_508), .B(n_154), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_500), .B(n_155), .Y(n_571) );
BUFx2_ASAP7_75t_L g572 ( .A(n_484), .Y(n_572) );
AND2x4_ASAP7_75t_L g573 ( .A(n_504), .B(n_156), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_518), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_477), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_479), .Y(n_576) );
CKINVDCx16_ASAP7_75t_R g577 ( .A(n_482), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_479), .Y(n_578) );
INVxp67_ASAP7_75t_R g579 ( .A(n_509), .Y(n_579) );
INVx3_ASAP7_75t_SL g580 ( .A(n_502), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_479), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_513), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_486), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_488), .Y(n_584) );
BUFx3_ASAP7_75t_L g585 ( .A(n_477), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_481), .B(n_157), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_519), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_491), .Y(n_588) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_510), .A2(n_158), .B(n_159), .Y(n_589) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_506), .A2(n_161), .B(n_165), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_502), .Y(n_591) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_477), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_514), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_517), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_514), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_516), .Y(n_596) );
OAI21x1_ASAP7_75t_L g597 ( .A1(n_511), .A2(n_171), .B(n_173), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_495), .B(n_174), .Y(n_598) );
AO21x1_ASAP7_75t_L g599 ( .A1(n_496), .A2(n_178), .B(n_179), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_492), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_526), .Y(n_601) );
OAI22xp33_ASAP7_75t_SL g602 ( .A1(n_498), .A2(n_184), .B1(n_185), .B2(n_186), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_526), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_498), .B(n_187), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_527), .Y(n_605) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_528), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_537), .B(n_188), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_532), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_534), .Y(n_609) );
BUFx2_ASAP7_75t_L g610 ( .A(n_537), .Y(n_610) );
AND2x4_ASAP7_75t_L g611 ( .A(n_540), .B(n_191), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_601), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_603), .B(n_195), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_577), .B(n_199), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_572), .A2(n_201), .B1(n_202), .B2(n_203), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_562), .B(n_206), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_551), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_555), .B(n_204), .Y(n_618) );
BUFx4f_ASAP7_75t_SL g619 ( .A(n_533), .Y(n_619) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_550), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_567), .B(n_205), .Y(n_621) );
BUFx3_ASAP7_75t_L g622 ( .A(n_528), .Y(n_622) );
BUFx4f_ASAP7_75t_SL g623 ( .A(n_539), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_530), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_546), .B(n_565), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_565), .B(n_566), .Y(n_626) );
OR2x2_ASAP7_75t_SL g627 ( .A(n_574), .B(n_549), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_566), .Y(n_628) );
INVx4_ASAP7_75t_R g629 ( .A(n_529), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_540), .B(n_544), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_545), .B(n_536), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_550), .B(n_552), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_570), .Y(n_633) );
AND2x4_ASAP7_75t_L g634 ( .A(n_531), .B(n_604), .Y(n_634) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_575), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_570), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_563), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_556), .B(n_559), .Y(n_638) );
OAI21xp33_ASAP7_75t_L g639 ( .A1(n_538), .A2(n_568), .B(n_535), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_563), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_561), .B(n_576), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_571), .B(n_560), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_586), .B(n_604), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_531), .B(n_564), .Y(n_644) );
INVxp67_ASAP7_75t_SL g645 ( .A(n_592), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_548), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_564), .B(n_569), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_569), .B(n_529), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_548), .Y(n_649) );
INVx2_ASAP7_75t_SL g650 ( .A(n_541), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_541), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_581), .B(n_578), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_542), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_568), .B(n_557), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_554), .B(n_598), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_535), .B(n_573), .Y(n_656) );
BUFx3_ASAP7_75t_L g657 ( .A(n_585), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_557), .B(n_595), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_592), .B(n_585), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_573), .B(n_589), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_589), .B(n_590), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_588), .Y(n_662) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_591), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_590), .B(n_553), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_553), .B(n_582), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_583), .B(n_587), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_543), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_584), .B(n_591), .Y(n_668) );
BUFx3_ASAP7_75t_L g669 ( .A(n_597), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_580), .B(n_596), .Y(n_670) );
OR2x2_ASAP7_75t_L g671 ( .A(n_580), .B(n_593), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g672 ( .A(n_602), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_558), .A2(n_600), .B1(n_599), .B2(n_594), .Y(n_673) );
INVx2_ASAP7_75t_SL g674 ( .A(n_547), .Y(n_674) );
NOR2x1p5_ASAP7_75t_L g675 ( .A(n_579), .B(n_558), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_537), .B(n_534), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_527), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_537), .B(n_534), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_527), .B(n_532), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_534), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_534), .Y(n_681) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_537), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_527), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_534), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_625), .B(n_610), .Y(n_685) );
BUFx2_ASAP7_75t_L g686 ( .A(n_623), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_631), .B(n_682), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_676), .Y(n_688) );
BUFx2_ASAP7_75t_L g689 ( .A(n_623), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_678), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_605), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_624), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_608), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_682), .B(n_642), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_677), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_641), .B(n_683), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_626), .B(n_609), .Y(n_697) );
BUFx2_ASAP7_75t_L g698 ( .A(n_648), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_612), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_680), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_681), .B(n_684), .Y(n_701) );
AND2x4_ASAP7_75t_L g702 ( .A(n_657), .B(n_620), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_679), .Y(n_703) );
INVx1_ASAP7_75t_SL g704 ( .A(n_620), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_630), .B(n_632), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_617), .B(n_638), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_638), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_628), .Y(n_708) );
OR2x2_ASAP7_75t_L g709 ( .A(n_641), .B(n_627), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_634), .B(n_647), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_637), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_640), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_662), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_653), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_651), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_663), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_655), .B(n_607), .Y(n_717) );
AND2x4_ASAP7_75t_L g718 ( .A(n_634), .B(n_644), .Y(n_718) );
INVxp67_ASAP7_75t_L g719 ( .A(n_635), .Y(n_719) );
AND2x4_ASAP7_75t_L g720 ( .A(n_644), .B(n_659), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_663), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_652), .Y(n_722) );
OR2x2_ASAP7_75t_L g723 ( .A(n_650), .B(n_646), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_614), .B(n_643), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_652), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_649), .B(n_636), .Y(n_726) );
AND2x4_ASAP7_75t_L g727 ( .A(n_666), .B(n_675), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_633), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_672), .B(n_621), .Y(n_729) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_645), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_613), .Y(n_731) );
INVx3_ASAP7_75t_L g732 ( .A(n_606), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_613), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_622), .Y(n_734) );
OR2x2_ASAP7_75t_L g735 ( .A(n_645), .B(n_658), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_660), .B(n_656), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_611), .B(n_622), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_611), .B(n_618), .Y(n_738) );
OR2x2_ASAP7_75t_L g739 ( .A(n_658), .B(n_654), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_621), .B(n_661), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_606), .B(n_672), .Y(n_741) );
BUFx2_ASAP7_75t_L g742 ( .A(n_619), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_616), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_706), .B(n_654), .Y(n_744) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_730), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_707), .B(n_639), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_685), .B(n_671), .Y(n_747) );
NAND2x1p5_ASAP7_75t_L g748 ( .A(n_686), .B(n_689), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_694), .B(n_670), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_687), .B(n_668), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_688), .B(n_664), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_691), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_736), .B(n_665), .Y(n_753) );
OR2x2_ASAP7_75t_L g754 ( .A(n_705), .B(n_616), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_693), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_690), .B(n_697), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_695), .Y(n_757) );
NOR2xp33_ASAP7_75t_SL g758 ( .A(n_742), .B(n_619), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_700), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_698), .B(n_669), .Y(n_760) );
OR2x2_ASAP7_75t_L g761 ( .A(n_720), .B(n_615), .Y(n_761) );
AND2x2_ASAP7_75t_L g762 ( .A(n_710), .B(n_674), .Y(n_762) );
AND2x4_ASAP7_75t_SL g763 ( .A(n_718), .B(n_629), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_701), .Y(n_764) );
AND2x4_ASAP7_75t_L g765 ( .A(n_727), .B(n_667), .Y(n_765) );
INVx2_ASAP7_75t_SL g766 ( .A(n_702), .Y(n_766) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_730), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_739), .B(n_673), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_722), .B(n_615), .Y(n_769) );
INVx3_ASAP7_75t_L g770 ( .A(n_727), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_717), .B(n_702), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_708), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_725), .B(n_713), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_699), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_713), .B(n_692), .Y(n_775) );
OAI31xp33_ASAP7_75t_L g776 ( .A1(n_729), .A2(n_709), .A3(n_738), .B(n_724), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_752), .Y(n_777) );
BUFx2_ASAP7_75t_L g778 ( .A(n_748), .Y(n_778) );
OR2x2_ASAP7_75t_L g779 ( .A(n_756), .B(n_704), .Y(n_779) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_745), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_771), .B(n_718), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_755), .Y(n_782) );
BUFx2_ASAP7_75t_L g783 ( .A(n_748), .Y(n_783) );
OR2x2_ASAP7_75t_L g784 ( .A(n_749), .B(n_704), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_757), .Y(n_785) );
OR2x2_ASAP7_75t_L g786 ( .A(n_751), .B(n_735), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_747), .B(n_741), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_772), .Y(n_788) );
INVx2_ASAP7_75t_SL g789 ( .A(n_763), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_759), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_750), .B(n_721), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_774), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_773), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_773), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_745), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_768), .B(n_703), .Y(n_796) );
INVxp67_ASAP7_75t_L g797 ( .A(n_767), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_767), .Y(n_798) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_775), .Y(n_799) );
AOI21xp33_ASAP7_75t_L g800 ( .A1(n_778), .A2(n_729), .B(n_746), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_777), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_782), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_785), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_788), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_790), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_796), .A2(n_768), .B1(n_776), .B2(n_740), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_792), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_796), .B(n_753), .Y(n_808) );
AOI31xp33_ASAP7_75t_L g809 ( .A1(n_789), .A2(n_763), .A3(n_761), .B(n_766), .Y(n_809) );
INVx3_ASAP7_75t_L g810 ( .A(n_783), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_799), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_799), .Y(n_812) );
INVxp67_ASAP7_75t_SL g813 ( .A(n_780), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_798), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_814), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_801), .B(n_797), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_802), .Y(n_817) );
BUFx2_ASAP7_75t_L g818 ( .A(n_810), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_810), .B(n_787), .Y(n_819) );
AOI211xp5_ASAP7_75t_L g820 ( .A1(n_800), .A2(n_758), .B(n_770), .C(n_766), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_803), .Y(n_821) );
AND2x2_ASAP7_75t_SL g822 ( .A(n_806), .B(n_770), .Y(n_822) );
INVx2_ASAP7_75t_L g823 ( .A(n_811), .Y(n_823) );
OAI21xp5_ASAP7_75t_L g824 ( .A1(n_820), .A2(n_809), .B(n_813), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g825 ( .A1(n_820), .A2(n_780), .B(n_797), .Y(n_825) );
AOI211xp5_ASAP7_75t_L g826 ( .A1(n_818), .A2(n_812), .B(n_769), .C(n_760), .Y(n_826) );
NOR3xp33_ASAP7_75t_L g827 ( .A(n_816), .B(n_714), .C(n_807), .Y(n_827) );
NOR4xp25_ASAP7_75t_L g828 ( .A(n_816), .B(n_821), .C(n_817), .D(n_815), .Y(n_828) );
O2A1O1Ixp33_ASAP7_75t_L g829 ( .A1(n_823), .A2(n_804), .B(n_805), .C(n_819), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_827), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_824), .A2(n_822), .B1(n_764), .B2(n_770), .Y(n_831) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_828), .Y(n_832) );
NOR3xp33_ASAP7_75t_L g833 ( .A(n_825), .B(n_733), .C(n_731), .Y(n_833) );
AND4x2_ASAP7_75t_L g834 ( .A(n_832), .B(n_826), .C(n_829), .D(n_779), .Y(n_834) );
NOR3xp33_ASAP7_75t_L g835 ( .A(n_830), .B(n_833), .C(n_831), .Y(n_835) );
NOR2x1_ASAP7_75t_L g836 ( .A(n_830), .B(n_781), .Y(n_836) );
BUFx2_ASAP7_75t_L g837 ( .A(n_836), .Y(n_837) );
NAND2x1p5_ASAP7_75t_L g838 ( .A(n_834), .B(n_784), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_838), .B(n_835), .Y(n_839) );
OAI21xp5_ASAP7_75t_L g840 ( .A1(n_837), .A2(n_808), .B(n_795), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_839), .B(n_791), .Y(n_841) );
AND2x4_ASAP7_75t_L g842 ( .A(n_840), .B(n_794), .Y(n_842) );
OAI21x1_ASAP7_75t_L g843 ( .A1(n_841), .A2(n_723), .B(n_711), .Y(n_843) );
OAI221xp5_ASAP7_75t_L g844 ( .A1(n_842), .A2(n_712), .B1(n_715), .B2(n_728), .C(n_719), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_843), .B(n_793), .Y(n_845) );
NAND3xp33_ASAP7_75t_L g846 ( .A(n_844), .B(n_743), .C(n_726), .Y(n_846) );
OAI21xp5_ASAP7_75t_SL g847 ( .A1(n_845), .A2(n_769), .B(n_737), .Y(n_847) );
OAI21xp5_ASAP7_75t_L g848 ( .A1(n_846), .A2(n_719), .B(n_754), .Y(n_848) );
AOI21xp5_ASAP7_75t_L g849 ( .A1(n_848), .A2(n_696), .B(n_744), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_847), .A2(n_734), .B1(n_765), .B2(n_716), .Y(n_850) );
OR2x6_ASAP7_75t_L g851 ( .A(n_849), .B(n_732), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_850), .B(n_732), .Y(n_852) );
OR2x4_ASAP7_75t_L g853 ( .A(n_852), .B(n_786), .Y(n_853) );
AOI21xp33_ASAP7_75t_L g854 ( .A1(n_853), .A2(n_851), .B(n_762), .Y(n_854) );
endmodule