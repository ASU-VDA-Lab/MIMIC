module fake_jpeg_14651_n_170 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_170);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_1),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_43),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_54),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_64),
.B(n_43),
.Y(n_73)
);

AO22x2_ASAP7_75t_L g114 ( 
.A1(n_73),
.A2(n_60),
.B1(n_6),
.B2(n_7),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_77),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_58),
.B1(n_64),
.B2(n_62),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_46),
.B1(n_56),
.B2(n_47),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_57),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_45),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_51),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx5_ASAP7_75t_SL g115 ( 
.A(n_91),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_100),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_104),
.B1(n_4),
.B2(n_7),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_60),
.B1(n_2),
.B2(n_3),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_114),
.B1(n_116),
.B2(n_101),
.Y(n_121)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_103),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_59),
.B1(n_52),
.B2(n_49),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_84),
.B(n_1),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_107),
.B(n_110),
.Y(n_130)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_108),
.A2(n_109),
.B1(n_4),
.B2(n_6),
.Y(n_119)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_113),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_117),
.B(n_9),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_131),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_29),
.B1(n_40),
.B2(n_39),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_8),
.Y(n_126)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_114),
.A2(n_28),
.B1(n_36),
.B2(n_35),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_114),
.C(n_104),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_136),
.Y(n_139)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_98),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_137),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_138),
.A2(n_119),
.B1(n_127),
.B2(n_120),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_133),
.B(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_142),
.A2(n_134),
.B1(n_129),
.B2(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_142),
.A2(n_136),
.B1(n_128),
.B2(n_95),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_105),
.Y(n_152)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_122),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_139),
.C(n_140),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_145),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_152),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_150),
.B(n_155),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_153),
.A2(n_151),
.B(n_148),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_156),
.B(n_157),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_106),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_111),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_8),
.C(n_9),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_10),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_10),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_12),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_13),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_14),
.B(n_15),
.Y(n_167)
);

OAI321xp33_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_16),
.A3(n_18),
.B1(n_19),
.B2(n_22),
.C(n_27),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_120),
.Y(n_169)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_169),
.B(n_30),
.CI(n_31),
.CON(n_170),
.SN(n_170)
);


endmodule