module fake_netlist_6_83_n_868 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_868);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_868;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_800;
wire n_779;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_796;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_678;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_102),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_53),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_150),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_174),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_54),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_38),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_196),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_93),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_95),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_198),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_48),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_43),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_192),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_183),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_14),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_159),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_141),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_101),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_56),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_94),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_166),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_14),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_119),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_136),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_12),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_117),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_177),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_190),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_85),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_71),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_185),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_134),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_115),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_40),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_13),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_180),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_2),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_78),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_57),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_87),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_34),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_97),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_16),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_33),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_47),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_195),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_69),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_124),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_41),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_147),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_160),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_83),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_1),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_201),
.Y(n_262)
);

BUFx2_ASAP7_75t_SL g263 ( 
.A(n_88),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_74),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_111),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_121),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_142),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_65),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_122),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_76),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_108),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_138),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_173),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_77),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_168),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_197),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_116),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_72),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_61),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_205),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_206),
.Y(n_281)
);

INVxp33_ASAP7_75t_SL g282 ( 
.A(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_221),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_228),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_221),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_229),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_221),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_221),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_261),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_221),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_221),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_242),
.Y(n_293)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_213),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_214),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_230),
.B(n_0),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_225),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_207),
.Y(n_299)
);

INVxp33_ASAP7_75t_SL g300 ( 
.A(n_263),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_227),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_211),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_208),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_233),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_234),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_211),
.Y(n_306)
);

NAND2xp33_ASAP7_75t_R g307 ( 
.A(n_209),
.B(n_0),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_240),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_245),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_215),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_248),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_266),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_277),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_253),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_210),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_264),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_274),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_212),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_216),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_237),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_217),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_271),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_252),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_218),
.B(n_1),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_219),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_256),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_220),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_329),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_290),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_301),
.Y(n_334)
);

NAND2xp33_ASAP7_75t_SL g335 ( 
.A(n_307),
.B(n_271),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_304),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_308),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_280),
.B(n_222),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_309),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_311),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_325),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_317),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_318),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_284),
.B(n_223),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_298),
.B(n_315),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_321),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_283),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_281),
.B(n_224),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_285),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_294),
.B(n_226),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_288),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_302),
.B(n_231),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_306),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_325),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_289),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_299),
.B(n_278),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_305),
.A2(n_276),
.B1(n_273),
.B2(n_272),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_287),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_291),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_292),
.Y(n_361)
);

OA21x2_ASAP7_75t_L g362 ( 
.A1(n_323),
.A2(n_326),
.B(n_293),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_300),
.B(n_297),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_293),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_295),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_312),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_286),
.Y(n_367)
);

AND2x6_ASAP7_75t_L g368 ( 
.A(n_327),
.B(n_271),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_300),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_303),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_320),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_320),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_316),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_319),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_330),
.B(n_235),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_324),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_324),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_328),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_330),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_305),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_365),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_353),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_310),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_282),
.Y(n_385)
);

INVxp33_ASAP7_75t_L g386 ( 
.A(n_359),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_282),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_343),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_354),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_343),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_351),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_373),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_341),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_345),
.B(n_313),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_236),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_373),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_238),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_373),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_341),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_341),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_345),
.B(n_239),
.Y(n_402)
);

AND2x2_ASAP7_75t_SL g403 ( 
.A(n_363),
.B(n_370),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_332),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_360),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_373),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_344),
.B(n_241),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_366),
.B(n_243),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_376),
.B(n_271),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_355),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_362),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_246),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_355),
.Y(n_413)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_376),
.Y(n_414)
);

NAND3xp33_ASAP7_75t_L g415 ( 
.A(n_367),
.B(n_366),
.C(n_359),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_334),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_381),
.B(n_247),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_376),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_333),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_368),
.B(n_249),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_336),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_337),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_355),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_335),
.A2(n_262),
.B1(n_255),
.B2(n_257),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_360),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_368),
.B(n_254),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_360),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_362),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_372),
.B(n_258),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_340),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_362),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_342),
.Y(n_433)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_368),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_346),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_377),
.B(n_259),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_368),
.B(n_260),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_347),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_335),
.A2(n_269),
.B1(n_265),
.B2(n_267),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_348),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_331),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_376),
.B(n_256),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_350),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_378),
.A2(n_270),
.B1(n_268),
.B2(n_314),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_352),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_356),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_361),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_364),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_395),
.B(n_370),
.Y(n_449)
);

NAND2x1p5_ASAP7_75t_L g450 ( 
.A(n_396),
.B(n_374),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_395),
.B(n_374),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_388),
.B(n_379),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_382),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_389),
.B(n_380),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_432),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_410),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_403),
.A2(n_358),
.B1(n_375),
.B2(n_338),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_388),
.B(n_364),
.Y(n_458)
);

A2O1A1Ixp33_ASAP7_75t_L g459 ( 
.A1(n_432),
.A2(n_357),
.B(n_349),
.C(n_256),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_410),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_404),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_384),
.Y(n_462)
);

NAND2x1_ASAP7_75t_L g463 ( 
.A(n_411),
.B(n_368),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_390),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_413),
.Y(n_465)
);

AO22x2_ASAP7_75t_L g466 ( 
.A1(n_394),
.A2(n_290),
.B1(n_3),
.B2(n_4),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_416),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_390),
.B(n_22),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_413),
.Y(n_469)
);

AO22x2_ASAP7_75t_L g470 ( 
.A1(n_415),
.A2(n_444),
.B1(n_383),
.B2(n_385),
.Y(n_470)
);

NAND2x1p5_ASAP7_75t_L g471 ( 
.A(n_396),
.B(n_23),
.Y(n_471)
);

NAND2x1p5_ASAP7_75t_L g472 ( 
.A(n_398),
.B(n_24),
.Y(n_472)
);

AO22x2_ASAP7_75t_L g473 ( 
.A1(n_391),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_411),
.B(n_429),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_421),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_403),
.A2(n_314),
.B1(n_313),
.B2(n_333),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_422),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_386),
.B(n_5),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_386),
.B(n_5),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_425),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_427),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_387),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_423),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_392),
.Y(n_484)
);

OR2x6_ASAP7_75t_SL g485 ( 
.A(n_406),
.B(n_6),
.Y(n_485)
);

OAI221xp5_ASAP7_75t_L g486 ( 
.A1(n_402),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_387),
.A2(n_397),
.B1(n_436),
.B2(n_430),
.Y(n_487)
);

AO22x2_ASAP7_75t_L g488 ( 
.A1(n_442),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_431),
.Y(n_489)
);

BUFx6f_ASAP7_75t_SL g490 ( 
.A(n_397),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_448),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_408),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_433),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_417),
.B(n_10),
.Y(n_494)
);

OAI22xp33_ASAP7_75t_SL g495 ( 
.A1(n_442),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_448),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_435),
.B(n_25),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_411),
.B(n_26),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_425),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_398),
.B(n_11),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_414),
.B(n_27),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_438),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_411),
.B(n_28),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_419),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_412),
.A2(n_113),
.B1(n_202),
.B2(n_200),
.Y(n_505)
);

BUFx8_ASAP7_75t_L g506 ( 
.A(n_441),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_446),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_414),
.Y(n_508)
);

AO22x2_ASAP7_75t_L g509 ( 
.A1(n_409),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_440),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_429),
.B(n_29),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_445),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_447),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_418),
.B(n_15),
.Y(n_514)
);

AO22x2_ASAP7_75t_L g515 ( 
.A1(n_409),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_405),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_487),
.B(n_418),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_449),
.B(n_407),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_451),
.B(n_457),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_462),
.B(n_434),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_484),
.B(n_434),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_492),
.B(n_434),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_464),
.B(n_468),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_464),
.B(n_434),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_468),
.B(n_412),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_455),
.B(n_429),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_482),
.B(n_430),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_452),
.B(n_436),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_452),
.B(n_443),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_458),
.B(n_443),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_458),
.B(n_429),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_454),
.B(n_424),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_450),
.B(n_439),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_494),
.B(n_420),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_497),
.B(n_510),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_478),
.B(n_405),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_455),
.B(n_428),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_497),
.B(n_426),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_513),
.B(n_437),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_453),
.B(n_428),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_SL g541 ( 
.A(n_508),
.B(n_400),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_461),
.B(n_400),
.Y(n_542)
);

NAND2xp33_ASAP7_75t_SL g543 ( 
.A(n_490),
.B(n_401),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_474),
.B(n_399),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_467),
.B(n_393),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_475),
.B(n_399),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_477),
.B(n_30),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_481),
.B(n_31),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_476),
.B(n_17),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_489),
.B(n_32),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_SL g551 ( 
.A(n_479),
.B(n_18),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_493),
.B(n_35),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_502),
.B(n_36),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_512),
.B(n_37),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_491),
.B(n_39),
.Y(n_555)
);

NAND2xp33_ASAP7_75t_SL g556 ( 
.A(n_514),
.B(n_19),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_507),
.B(n_516),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_SL g558 ( 
.A(n_463),
.B(n_20),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_496),
.B(n_42),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_501),
.B(n_44),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_495),
.B(n_45),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_483),
.B(n_46),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_503),
.B(n_49),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_480),
.B(n_50),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_SL g565 ( 
.A(n_463),
.B(n_20),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_SL g566 ( 
.A(n_504),
.B(n_21),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_511),
.B(n_480),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_499),
.B(n_51),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_505),
.B(n_52),
.Y(n_569)
);

NAND2xp33_ASAP7_75t_SL g570 ( 
.A(n_470),
.B(n_21),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_456),
.B(n_460),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_465),
.B(n_55),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_SL g573 ( 
.A(n_470),
.B(n_469),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_537),
.Y(n_574)
);

NAND3xp33_ASAP7_75t_L g575 ( 
.A(n_549),
.B(n_500),
.C(n_506),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_518),
.B(n_498),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_526),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_571),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_525),
.A2(n_498),
.B1(n_500),
.B2(n_466),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_536),
.B(n_527),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_528),
.B(n_459),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_R g582 ( 
.A(n_541),
.B(n_506),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_570),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_543),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_542),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_566),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_517),
.A2(n_519),
.B(n_538),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_544),
.A2(n_472),
.B(n_471),
.Y(n_588)
);

AOI211x1_ASAP7_75t_L g589 ( 
.A1(n_561),
.A2(n_486),
.B(n_473),
.C(n_515),
.Y(n_589)
);

CKINVDCx11_ASAP7_75t_R g590 ( 
.A(n_564),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_564),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_523),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_551),
.Y(n_593)
);

NOR2xp67_ASAP7_75t_SL g594 ( 
.A(n_569),
.B(n_529),
.Y(n_594)
);

OAI21x1_ASAP7_75t_L g595 ( 
.A1(n_567),
.A2(n_498),
.B(n_509),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_531),
.A2(n_534),
.B(n_539),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_564),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_532),
.B(n_466),
.C(n_485),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_530),
.B(n_58),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_535),
.B(n_488),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_540),
.B(n_488),
.Y(n_601)
);

INVxp67_ASAP7_75t_SL g602 ( 
.A(n_557),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_533),
.B(n_473),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_545),
.Y(n_604)
);

BUFx4_ASAP7_75t_SL g605 ( 
.A(n_573),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_546),
.A2(n_59),
.B(n_60),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_522),
.B(n_203),
.Y(n_607)
);

AOI21x1_ASAP7_75t_SL g608 ( 
.A1(n_558),
.A2(n_62),
.B(n_63),
.Y(n_608)
);

OAI21x1_ASAP7_75t_SL g609 ( 
.A1(n_565),
.A2(n_64),
.B(n_66),
.Y(n_609)
);

OAI21x1_ASAP7_75t_SL g610 ( 
.A1(n_556),
.A2(n_67),
.B(n_68),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_563),
.B(n_70),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_521),
.B(n_73),
.Y(n_612)
);

AOI221x1_ASAP7_75t_L g613 ( 
.A1(n_560),
.A2(n_75),
.B1(n_79),
.B2(n_80),
.C(n_81),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_524),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_520),
.B(n_82),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_547),
.A2(n_84),
.B1(n_86),
.B2(n_89),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_555),
.Y(n_617)
);

BUFx2_ASAP7_75t_SL g618 ( 
.A(n_559),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_548),
.Y(n_619)
);

AO21x2_ASAP7_75t_L g620 ( 
.A1(n_587),
.A2(n_554),
.B(n_553),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_592),
.B(n_550),
.Y(n_621)
);

NAND3xp33_ASAP7_75t_L g622 ( 
.A(n_587),
.B(n_552),
.C(n_562),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_577),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_580),
.B(n_568),
.Y(n_624)
);

NOR2xp67_ASAP7_75t_SL g625 ( 
.A(n_575),
.B(n_572),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_588),
.A2(n_90),
.B(n_91),
.Y(n_626)
);

OAI22xp33_ASAP7_75t_L g627 ( 
.A1(n_579),
.A2(n_92),
.B1(n_96),
.B2(n_98),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_581),
.A2(n_199),
.B(n_100),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_606),
.A2(n_99),
.B(n_103),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_584),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_591),
.B(n_194),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_SL g632 ( 
.A1(n_598),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_577),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_593),
.B(n_107),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_578),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_574),
.B(n_109),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_590),
.Y(n_637)
);

OAI21x1_ASAP7_75t_L g638 ( 
.A1(n_595),
.A2(n_596),
.B(n_608),
.Y(n_638)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_608),
.A2(n_110),
.B(n_112),
.Y(n_639)
);

OAI21x1_ASAP7_75t_SL g640 ( 
.A1(n_609),
.A2(n_114),
.B(n_123),
.Y(n_640)
);

OAI21x1_ASAP7_75t_L g641 ( 
.A1(n_576),
.A2(n_125),
.B(n_126),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g642 ( 
.A1(n_591),
.A2(n_127),
.B(n_128),
.Y(n_642)
);

AO31x2_ASAP7_75t_L g643 ( 
.A1(n_613),
.A2(n_129),
.A3(n_130),
.B(n_131),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_597),
.B(n_583),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_597),
.A2(n_132),
.B(n_133),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_599),
.B(n_135),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_602),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_602),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_599),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_585),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_604),
.Y(n_651)
);

AOI221xp5_ASAP7_75t_L g652 ( 
.A1(n_589),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.C(n_143),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_590),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_586),
.B(n_193),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_601),
.B(n_144),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_603),
.A2(n_145),
.B1(n_146),
.B2(n_148),
.Y(n_656)
);

AO32x2_ASAP7_75t_L g657 ( 
.A1(n_619),
.A2(n_149),
.A3(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_657)
);

INVx6_ASAP7_75t_SL g658 ( 
.A(n_582),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_584),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_582),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_617),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_635),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_623),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_633),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_651),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_650),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_644),
.B(n_600),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_647),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_649),
.Y(n_669)
);

AOI21x1_ASAP7_75t_L g670 ( 
.A1(n_638),
.A2(n_594),
.B(n_611),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_661),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_631),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_648),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_649),
.B(n_612),
.Y(n_674)
);

OA21x2_ASAP7_75t_L g675 ( 
.A1(n_639),
.A2(n_611),
.B(n_610),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_631),
.Y(n_676)
);

OAI21x1_ASAP7_75t_L g677 ( 
.A1(n_626),
.A2(n_615),
.B(n_607),
.Y(n_677)
);

AO21x2_ASAP7_75t_L g678 ( 
.A1(n_622),
.A2(n_616),
.B(n_614),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_644),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_661),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_636),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_645),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_630),
.Y(n_683)
);

BUFx4f_ASAP7_75t_L g684 ( 
.A(n_646),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_646),
.B(n_617),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_629),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_624),
.B(n_605),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_636),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_661),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_642),
.A2(n_605),
.B(n_618),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_621),
.Y(n_691)
);

AOI21x1_ASAP7_75t_L g692 ( 
.A1(n_622),
.A2(n_154),
.B(n_155),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_641),
.Y(n_693)
);

AO21x1_ASAP7_75t_SL g694 ( 
.A1(n_628),
.A2(n_156),
.B(n_157),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_655),
.Y(n_695)
);

OA21x2_ASAP7_75t_L g696 ( 
.A1(n_628),
.A2(n_158),
.B(n_161),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_654),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_697)
);

OA21x2_ASAP7_75t_L g698 ( 
.A1(n_652),
.A2(n_167),
.B(n_169),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_659),
.Y(n_699)
);

AOI21x1_ASAP7_75t_L g700 ( 
.A1(n_625),
.A2(n_170),
.B(n_171),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_620),
.Y(n_701)
);

AO21x1_ASAP7_75t_SL g702 ( 
.A1(n_656),
.A2(n_172),
.B(n_175),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_657),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_657),
.Y(n_704)
);

OAI21x1_ASAP7_75t_L g705 ( 
.A1(n_640),
.A2(n_176),
.B(n_178),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_637),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_657),
.Y(n_707)
);

NAND2xp33_ASAP7_75t_R g708 ( 
.A(n_685),
.B(n_660),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_685),
.B(n_672),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_679),
.B(n_624),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_SL g711 ( 
.A(n_704),
.B(n_637),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_R g712 ( 
.A(n_684),
.B(n_653),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_SL g713 ( 
.A(n_704),
.B(n_654),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_685),
.B(n_672),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_679),
.B(n_667),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_R g716 ( 
.A(n_684),
.B(n_634),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_666),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_667),
.B(n_632),
.Y(n_718)
);

NAND2xp33_ASAP7_75t_R g719 ( 
.A(n_695),
.B(n_658),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_668),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_690),
.B(n_627),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_691),
.B(n_632),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_666),
.B(n_643),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_681),
.B(n_652),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_672),
.B(n_643),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_688),
.B(n_627),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_671),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_R g728 ( 
.A(n_684),
.B(n_658),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_662),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_663),
.B(n_620),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_687),
.B(n_674),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_699),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_673),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_R g734 ( 
.A(n_676),
.B(n_179),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_664),
.B(n_643),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_689),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_687),
.B(n_683),
.Y(n_737)
);

XNOR2xp5_ASAP7_75t_L g738 ( 
.A(n_706),
.B(n_181),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_665),
.B(n_182),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_674),
.B(n_184),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_R g741 ( 
.A(n_698),
.B(n_186),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_706),
.B(n_680),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_731),
.B(n_703),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_715),
.B(n_704),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_709),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_710),
.B(n_729),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_713),
.A2(n_702),
.B1(n_698),
.B2(n_694),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_720),
.B(n_703),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_733),
.B(n_704),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_730),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_735),
.B(n_701),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_709),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_725),
.B(n_704),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_725),
.B(n_707),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_736),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_723),
.Y(n_756)
);

NOR2x1_ASAP7_75t_SL g757 ( 
.A(n_721),
.B(n_707),
.Y(n_757)
);

CKINVDCx6p67_ASAP7_75t_R g758 ( 
.A(n_740),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_717),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_742),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_722),
.B(n_714),
.Y(n_761)
);

AND2x2_ASAP7_75t_SL g762 ( 
.A(n_741),
.B(n_698),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_726),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_727),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_714),
.B(n_696),
.Y(n_765)
);

NOR3xp33_ASAP7_75t_L g766 ( 
.A(n_737),
.B(n_697),
.C(n_700),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_726),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_721),
.Y(n_768)
);

BUFx2_ASAP7_75t_L g769 ( 
.A(n_711),
.Y(n_769)
);

AND2x4_ASAP7_75t_SL g770 ( 
.A(n_721),
.B(n_669),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_759),
.Y(n_771)
);

BUFx8_ASAP7_75t_L g772 ( 
.A(n_769),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_753),
.B(n_696),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_752),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_748),
.Y(n_775)
);

AND2x2_ASAP7_75t_SL g776 ( 
.A(n_762),
.B(n_696),
.Y(n_776)
);

NAND2x1p5_ASAP7_75t_SL g777 ( 
.A(n_763),
.B(n_765),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_SL g778 ( 
.A1(n_762),
.A2(n_716),
.B1(n_718),
.B2(n_734),
.Y(n_778)
);

AO21x2_ASAP7_75t_L g779 ( 
.A1(n_766),
.A2(n_693),
.B(n_692),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_753),
.B(n_732),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_748),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_749),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_749),
.Y(n_783)
);

AOI211xp5_ASAP7_75t_SL g784 ( 
.A1(n_768),
.A2(n_724),
.B(n_739),
.C(n_676),
.Y(n_784)
);

OAI222xp33_ASAP7_75t_L g785 ( 
.A1(n_769),
.A2(n_738),
.B1(n_700),
.B2(n_692),
.C1(n_676),
.C2(n_670),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_767),
.B(n_678),
.Y(n_786)
);

INVx5_ASAP7_75t_SL g787 ( 
.A(n_758),
.Y(n_787)
);

NAND2xp67_ASAP7_75t_L g788 ( 
.A(n_780),
.B(n_770),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_771),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_771),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_775),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_780),
.B(n_743),
.Y(n_792)
);

AND2x4_ASAP7_75t_SL g793 ( 
.A(n_773),
.B(n_758),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_775),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_783),
.B(n_743),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_774),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_782),
.B(n_767),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_781),
.Y(n_798)
);

NOR2x1_ASAP7_75t_L g799 ( 
.A(n_796),
.B(n_785),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_797),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_793),
.Y(n_801)
);

NAND2xp33_ASAP7_75t_SL g802 ( 
.A(n_792),
.B(n_708),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_793),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_801),
.B(n_795),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_800),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_803),
.B(n_787),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_799),
.A2(n_778),
.B1(n_776),
.B2(n_787),
.Y(n_807)
);

AOI21xp33_ASAP7_75t_SL g808 ( 
.A1(n_807),
.A2(n_760),
.B(n_719),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_805),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_806),
.B(n_798),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_809),
.B(n_804),
.Y(n_811)
);

NOR2x1_ASAP7_75t_SL g812 ( 
.A(n_810),
.B(n_807),
.Y(n_812)
);

NAND2x1_ASAP7_75t_L g813 ( 
.A(n_810),
.B(n_791),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_811),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_813),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_812),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_811),
.Y(n_817)
);

NAND3xp33_ASAP7_75t_L g818 ( 
.A(n_816),
.B(n_808),
.C(n_802),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_814),
.B(n_787),
.Y(n_819)
);

NAND3xp33_ASAP7_75t_SL g820 ( 
.A(n_817),
.B(n_712),
.C(n_728),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_815),
.Y(n_821)
);

OAI21xp33_ASAP7_75t_L g822 ( 
.A1(n_816),
.A2(n_768),
.B(n_776),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_816),
.B(n_787),
.Y(n_823)
);

NAND4xp25_ASAP7_75t_L g824 ( 
.A(n_816),
.B(n_784),
.C(n_764),
.D(n_747),
.Y(n_824)
);

NOR3xp33_ASAP7_75t_SL g825 ( 
.A(n_818),
.B(n_746),
.C(n_772),
.Y(n_825)
);

CKINVDCx6p67_ASAP7_75t_R g826 ( 
.A(n_823),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_SL g827 ( 
.A1(n_821),
.A2(n_680),
.B1(n_772),
.B2(n_755),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_819),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_820),
.A2(n_822),
.B(n_824),
.Y(n_829)
);

AOI31xp33_ASAP7_75t_L g830 ( 
.A1(n_818),
.A2(n_772),
.A3(n_794),
.B(n_798),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_818),
.A2(n_779),
.B1(n_770),
.B2(n_774),
.Y(n_831)
);

AOI221xp5_ASAP7_75t_L g832 ( 
.A1(n_818),
.A2(n_777),
.B1(n_790),
.B2(n_789),
.C(n_779),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_828),
.B(n_794),
.Y(n_833)
);

NOR2x1_ASAP7_75t_L g834 ( 
.A(n_830),
.B(n_779),
.Y(n_834)
);

BUFx12f_ASAP7_75t_L g835 ( 
.A(n_826),
.Y(n_835)
);

INVxp67_ASAP7_75t_SL g836 ( 
.A(n_827),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_829),
.B(n_705),
.C(n_786),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_831),
.Y(n_838)
);

NAND2x1p5_ASAP7_75t_L g839 ( 
.A(n_825),
.B(n_705),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_832),
.B(n_761),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_828),
.B(n_761),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_835),
.B(n_745),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_836),
.B(n_782),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_L g844 ( 
.A(n_838),
.B(n_750),
.C(n_763),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_834),
.B(n_745),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_841),
.B(n_833),
.Y(n_846)
);

NAND2xp33_ASAP7_75t_SL g847 ( 
.A(n_840),
.B(n_669),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_R g848 ( 
.A(n_839),
.B(n_187),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_R g849 ( 
.A(n_837),
.B(n_188),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_843),
.Y(n_850)
);

OA22x2_ASAP7_75t_L g851 ( 
.A1(n_842),
.A2(n_745),
.B1(n_781),
.B2(n_750),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_846),
.Y(n_852)
);

AOI222xp33_ASAP7_75t_L g853 ( 
.A1(n_847),
.A2(n_757),
.B1(n_773),
.B2(n_690),
.C1(n_694),
.C2(n_702),
.Y(n_853)
);

AOI211xp5_ASAP7_75t_L g854 ( 
.A1(n_845),
.A2(n_669),
.B(n_765),
.C(n_788),
.Y(n_854)
);

NAND4xp25_ASAP7_75t_L g855 ( 
.A(n_844),
.B(n_848),
.C(n_849),
.D(n_752),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_850),
.Y(n_856)
);

NAND3x1_ASAP7_75t_L g857 ( 
.A(n_852),
.B(n_670),
.C(n_744),
.Y(n_857)
);

AO21x2_ASAP7_75t_L g858 ( 
.A1(n_855),
.A2(n_777),
.B(n_757),
.Y(n_858)
);

XNOR2x1_ASAP7_75t_L g859 ( 
.A(n_851),
.B(n_189),
.Y(n_859)
);

XOR2xp5_ASAP7_75t_L g860 ( 
.A(n_859),
.B(n_854),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_856),
.B(n_858),
.Y(n_861)
);

NOR2x1_ASAP7_75t_L g862 ( 
.A(n_857),
.B(n_853),
.Y(n_862)
);

AOI31xp33_ASAP7_75t_L g863 ( 
.A1(n_861),
.A2(n_860),
.A3(n_862),
.B(n_783),
.Y(n_863)
);

OAI322xp33_ASAP7_75t_L g864 ( 
.A1(n_863),
.A2(n_693),
.A3(n_751),
.B1(n_669),
.B2(n_756),
.C1(n_682),
.C2(n_686),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_864),
.A2(n_678),
.B1(n_669),
.B2(n_756),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_865),
.Y(n_866)
);

OAI221xp5_ASAP7_75t_R g867 ( 
.A1(n_866),
.A2(n_191),
.B1(n_678),
.B2(n_677),
.C(n_675),
.Y(n_867)
);

AOI211xp5_ASAP7_75t_L g868 ( 
.A1(n_867),
.A2(n_677),
.B(n_751),
.C(n_754),
.Y(n_868)
);


endmodule