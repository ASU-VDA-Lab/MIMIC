module fake_jpeg_22841_n_257 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_11),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

AOI21xp33_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_0),
.B(n_1),
.Y(n_30)
);

NAND2xp33_ASAP7_75t_SL g50 ( 
.A(n_30),
.B(n_1),
.Y(n_50)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_32),
.Y(n_42)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_26),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_53),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_19),
.B1(n_28),
.B2(n_16),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_56),
.B1(n_24),
.B2(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_19),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_54),
.C(n_37),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_51),
.B(n_20),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_30),
.B(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_34),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_16),
.B1(n_17),
.B2(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_59),
.Y(n_63)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_65),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_79),
.B1(n_31),
.B2(n_39),
.Y(n_101)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_74),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_24),
.B1(n_29),
.B2(n_23),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_24),
.B1(n_23),
.B2(n_15),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_71),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_76),
.C(n_52),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_49),
.B1(n_50),
.B2(n_46),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_75),
.B(n_27),
.C(n_18),
.Y(n_91)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_47),
.A2(n_38),
.B(n_34),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_80),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

AO22x2_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_22),
.B1(n_27),
.B2(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_43),
.A2(n_15),
.B1(n_25),
.B2(n_14),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_81),
.A2(n_56),
.B1(n_43),
.B2(n_45),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_88),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_84),
.B(n_101),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_90),
.C(n_95),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_76),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_44),
.B1(n_58),
.B2(n_40),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_99),
.B1(n_79),
.B2(n_61),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_42),
.C(n_55),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_31),
.B(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_40),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_96),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_42),
.C(n_53),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_59),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_42),
.C(n_41),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_42),
.C(n_63),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_73),
.A2(n_79),
.B1(n_62),
.B2(n_74),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_61),
.Y(n_117)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_66),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_79),
.B(n_60),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_112),
.B(n_119),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_107),
.B(n_109),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_74),
.B1(n_65),
.B2(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_70),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_90),
.Y(n_136)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_122),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_123),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_70),
.B(n_14),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_100),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_120),
.Y(n_130)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_97),
.C(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_2),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_2),
.Y(n_147)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_128),
.Y(n_167)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_82),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_143),
.B(n_145),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_110),
.A2(n_93),
.B1(n_94),
.B2(n_92),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_124),
.B1(n_106),
.B2(n_120),
.Y(n_156)
);

AO22x1_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_89),
.B1(n_93),
.B2(n_84),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_104),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_147),
.B(n_110),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_152),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_132),
.A2(n_121),
.B1(n_116),
.B2(n_115),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_150),
.A2(n_156),
.B1(n_157),
.B2(n_163),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_136),
.B(n_116),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_121),
.B1(n_114),
.B2(n_107),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_105),
.B(n_119),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_161),
.A2(n_165),
.B(n_147),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_134),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_145),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_113),
.B1(n_109),
.B2(n_126),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_129),
.B(n_126),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_140),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_63),
.B(n_86),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_103),
.B1(n_86),
.B2(n_25),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_170),
.B1(n_77),
.B2(n_103),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_169),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_103),
.B1(n_77),
.B2(n_14),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_172),
.Y(n_190)
);

OAI21x1_ASAP7_75t_SL g172 ( 
.A1(n_161),
.A2(n_143),
.B(n_165),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_167),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_173),
.B(n_174),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

A2O1A1O1Ixp25_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_139),
.B(n_146),
.C(n_141),
.D(n_130),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_179),
.Y(n_196)
);

AO22x1_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_140),
.B1(n_137),
.B2(n_133),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_189),
.B(n_147),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_154),
.A2(n_133),
.B1(n_135),
.B2(n_128),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_183),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_155),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_182),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_195),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_157),
.B1(n_150),
.B2(n_158),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_198),
.B1(n_199),
.B2(n_184),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_152),
.B1(n_149),
.B2(n_160),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_160),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_186),
.C(n_189),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_148),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_188),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_203),
.A2(n_127),
.B(n_27),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_207),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_186),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_211),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_201),
.A2(n_180),
.B1(n_178),
.B2(n_176),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_213),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_178),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_217),
.B(n_203),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_22),
.C(n_27),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_215),
.C(n_195),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_22),
.C(n_18),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_18),
.B1(n_22),
.B2(n_4),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_202),
.Y(n_225)
);

XNOR2x1_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_8),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_220),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_191),
.C(n_196),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_223),
.C(n_215),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_196),
.C(n_194),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_207),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_217),
.A2(n_193),
.B(n_204),
.C(n_9),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_227),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_8),
.B(n_13),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_10),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_232),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_235),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_21),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_222),
.A2(n_7),
.B(n_13),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_237),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_21),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_219),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_238),
.A2(n_221),
.B1(n_6),
.B2(n_11),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_233),
.A2(n_223),
.B1(n_221),
.B2(n_224),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_244),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_242),
.A2(n_231),
.B1(n_3),
.B2(n_4),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_248),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_11),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_12),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_247),
.B(n_240),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_245),
.Y(n_253)
);

AOI322xp5_ASAP7_75t_L g255 ( 
.A1(n_253),
.A2(n_254),
.A3(n_252),
.B1(n_12),
.B2(n_4),
.C1(n_5),
.C2(n_3),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_241),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_255),
.B(n_2),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g257 ( 
.A(n_256),
.Y(n_257)
);


endmodule