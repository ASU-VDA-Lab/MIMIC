module fake_jpeg_10818_n_420 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_420);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_420;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx11_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_50),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_54),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_16),
.B(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_67),
.Y(n_109)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_56),
.Y(n_96)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_13),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_59),
.B(n_84),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_60),
.B(n_73),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_16),
.B(n_12),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_17),
.B(n_9),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_69),
.B(n_79),
.Y(n_127)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_76),
.Y(n_108)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_17),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_74),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_23),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_75),
.B(n_77),
.Y(n_138)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_23),
.B(n_9),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_45),
.B1(n_18),
.B2(n_37),
.Y(n_111)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_27),
.B(n_8),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_86),
.B(n_92),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_31),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_31),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_33),
.B1(n_46),
.B2(n_44),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_97),
.A2(n_122),
.B1(n_129),
.B2(n_83),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_49),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_98),
.B(n_121),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_53),
.B(n_33),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_101),
.B(n_83),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_48),
.A2(n_25),
.B1(n_39),
.B2(n_43),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_104),
.A2(n_114),
.B1(n_145),
.B2(n_80),
.Y(n_151)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_111),
.A2(n_131),
.B1(n_18),
.B2(n_26),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_63),
.A2(n_87),
.B1(n_91),
.B2(n_71),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_66),
.A2(n_44),
.B1(n_25),
.B2(n_39),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_72),
.A2(n_39),
.B1(n_25),
.B2(n_24),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_56),
.A2(n_43),
.B1(n_30),
.B2(n_32),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_85),
.B(n_32),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_85),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_81),
.A2(n_26),
.B1(n_30),
.B2(n_37),
.Y(n_145)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_54),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_151),
.A2(n_165),
.B1(n_143),
.B2(n_124),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_109),
.B(n_45),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_152),
.B(n_162),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_153),
.A2(n_78),
.B(n_52),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_157),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_108),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_155),
.B(n_163),
.C(n_100),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_125),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_142),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_158),
.B(n_169),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_89),
.B1(n_88),
.B2(n_74),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_159),
.A2(n_185),
.B1(n_100),
.B2(n_96),
.Y(n_197)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_50),
.C(n_49),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_164),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_122),
.A2(n_129),
.B1(n_97),
.B2(n_145),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_134),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_170),
.Y(n_196)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_116),
.B(n_90),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_107),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_173),
.A2(n_184),
.B1(n_132),
.B2(n_143),
.Y(n_202)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_90),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_175),
.B(n_180),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_102),
.B(n_0),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_176),
.B(n_187),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_112),
.B(n_0),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_178),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_113),
.B(n_1),
.Y(n_178)
);

BUFx8_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_181),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_182),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_126),
.B(n_140),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_186),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_106),
.A2(n_93),
.B1(n_4),
.B2(n_5),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_115),
.B(n_3),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_110),
.B(n_52),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_128),
.B(n_141),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_120),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_96),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_190),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_199),
.B1(n_184),
.B2(n_200),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g198 ( 
.A(n_156),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_153),
.A2(n_105),
.B1(n_124),
.B2(n_123),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_154),
.A2(n_132),
.B(n_139),
.C(n_99),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_200),
.A2(n_179),
.B(n_170),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_165),
.A2(n_139),
.B1(n_136),
.B2(n_135),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_202),
.A2(n_203),
.B1(n_212),
.B2(n_166),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_215),
.C(n_219),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_151),
.A2(n_123),
.B1(n_136),
.B2(n_130),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_155),
.B(n_117),
.C(n_103),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_216),
.B(n_218),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_181),
.C(n_183),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_181),
.A2(n_3),
.B(n_4),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_4),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_225),
.A2(n_201),
.B1(n_212),
.B2(n_219),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_226),
.B(n_233),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_177),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_234),
.Y(n_265)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_229),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_230),
.A2(n_241),
.B(n_220),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_221),
.B(n_178),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_208),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_191),
.B(n_186),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_235),
.B(n_238),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_208),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_237),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_171),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_196),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_239),
.A2(n_243),
.B1(n_224),
.B2(n_222),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_196),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_240),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_223),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_242),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_203),
.A2(n_172),
.B1(n_182),
.B2(n_150),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_209),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_251),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_191),
.B(n_149),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_246),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_160),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_216),
.B(n_205),
.Y(n_267)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_222),
.Y(n_250)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_179),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_192),
.Y(n_252)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_248),
.B(n_210),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_227),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_256),
.A2(n_270),
.B1(n_271),
.B2(n_243),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_232),
.B(n_245),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_260),
.A2(n_269),
.B(n_238),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_215),
.C(n_214),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_266),
.B(n_207),
.C(n_193),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_267),
.B(n_234),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_232),
.A2(n_218),
.B(n_224),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_225),
.A2(n_199),
.B1(n_213),
.B2(n_205),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_237),
.A2(n_197),
.B1(n_150),
.B2(n_213),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_274),
.Y(n_283)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_228),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_279),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_259),
.A2(n_273),
.B1(n_239),
.B2(n_276),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_281),
.A2(n_284),
.B(n_293),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_277),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_285),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_275),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_244),
.Y(n_286)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_286),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_277),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_291),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_260),
.A2(n_236),
.B(n_240),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_288),
.A2(n_295),
.B(n_272),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_297),
.C(n_303),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_265),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_296),
.B1(n_274),
.B2(n_269),
.Y(n_308)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_257),
.Y(n_294)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_294),
.Y(n_316)
);

AO32x1_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_242),
.A3(n_251),
.B1(n_230),
.B2(n_247),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_271),
.A2(n_246),
.B1(n_233),
.B2(n_235),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_224),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_298),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_261),
.B(n_250),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_253),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_252),
.Y(n_300)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_300),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_252),
.Y(n_301)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_301),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_264),
.Y(n_302)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_302),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_254),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_304),
.B(n_324),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_300),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_318),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_266),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_312),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_308),
.A2(n_320),
.B1(n_298),
.B2(n_268),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_262),
.C(n_278),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_309),
.C(n_312),
.Y(n_332)
);

AO22x1_ASAP7_75t_L g341 ( 
.A1(n_311),
.A2(n_295),
.B1(n_289),
.B2(n_294),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_279),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_288),
.A2(n_275),
.B(n_263),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_313),
.A2(n_295),
.B(n_285),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_283),
.A2(n_258),
.B1(n_257),
.B2(n_262),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_296),
.A2(n_258),
.B1(n_268),
.B2(n_229),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_286),
.B(n_193),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_323),
.B(n_253),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_293),
.A2(n_281),
.B(n_283),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_284),
.Y(n_331)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_280),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_327),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_301),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_333),
.Y(n_360)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_331),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_335),
.C(n_337),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_299),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_287),
.C(n_282),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_336),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_291),
.C(n_285),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_314),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_338),
.B(n_344),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_340),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_341),
.A2(n_315),
.B(n_313),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_325),
.B(n_231),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_342),
.B(n_343),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_292),
.C(n_289),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_280),
.C(n_206),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_345),
.B(n_326),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_346),
.A2(n_321),
.B1(n_318),
.B2(n_316),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_319),
.B(n_207),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_347),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_352),
.A2(n_341),
.B(n_345),
.Y(n_369)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_353),
.Y(n_368)
);

INVx13_ASAP7_75t_L g354 ( 
.A(n_344),
.Y(n_354)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_343),
.A2(n_321),
.B1(n_306),
.B2(n_315),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_355),
.A2(n_357),
.B1(n_323),
.B2(n_327),
.Y(n_372)
);

NOR3xp33_ASAP7_75t_SL g357 ( 
.A(n_334),
.B(n_306),
.C(n_311),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_329),
.Y(n_358)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_358),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_333),
.B(n_319),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_359),
.B(n_361),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_337),
.A2(n_335),
.B1(n_328),
.B2(n_324),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_362),
.A2(n_339),
.B1(n_317),
.B2(n_316),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_349),
.Y(n_365)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_365),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_350),
.B(n_332),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_367),
.B(n_375),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_369),
.A2(n_361),
.B(n_360),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_349),
.B(n_339),
.C(n_330),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_374),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_372),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_373),
.A2(n_368),
.B1(n_378),
.B2(n_370),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_268),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_348),
.B(n_253),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_351),
.Y(n_376)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_376),
.Y(n_385)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_358),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_377),
.B(n_355),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_359),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_390),
.Y(n_395)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_381),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_378),
.B(n_360),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_317),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_369),
.A2(n_363),
.B(n_362),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_386),
.A2(n_388),
.B(n_368),
.Y(n_394)
);

AOI221xp5_ASAP7_75t_L g387 ( 
.A1(n_373),
.A2(n_356),
.B1(n_363),
.B2(n_353),
.C(n_357),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_387),
.B(n_206),
.Y(n_398)
);

NOR2x1_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_371),
.Y(n_391)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_391),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_385),
.B(n_366),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_393),
.B(n_398),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_400),
.Y(n_402)
);

AND2x2_ASAP7_75t_SL g401 ( 
.A(n_396),
.B(n_390),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_384),
.A2(n_354),
.B1(n_194),
.B2(n_204),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_397),
.A2(n_399),
.B(n_388),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_204),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_379),
.B(n_167),
.Y(n_400)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_401),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_381),
.Y(n_403)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_403),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_386),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_404),
.B(n_407),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_406),
.A2(n_392),
.B1(n_393),
.B2(n_380),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_411),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_173),
.C(n_167),
.Y(n_411)
);

AOI21x1_ASAP7_75t_SL g413 ( 
.A1(n_410),
.A2(n_405),
.B(n_401),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_413),
.A2(n_415),
.B(n_5),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_409),
.A2(n_161),
.B(n_180),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_414),
.A2(n_412),
.B1(n_168),
.B2(n_7),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_416),
.A2(n_417),
.B1(n_5),
.B2(n_6),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_418),
.B(n_6),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_419),
.B(n_6),
.Y(n_420)
);


endmodule