module real_jpeg_28838_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_286, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_286;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_281;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_105;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_202;
wire n_244;
wire n_179;
wire n_167;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_283;
wire n_81;
wire n_85;
wire n_181;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g73 ( 
.A(n_0),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_1),
.Y(n_100)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_1),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_4),
.A2(n_18),
.B1(n_19),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_4),
.A2(n_23),
.B1(n_26),
.B2(n_33),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_4),
.A2(n_33),
.B1(n_71),
.B2(n_72),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_4),
.A2(n_33),
.B1(n_50),
.B2(n_52),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_6),
.A2(n_18),
.B1(n_19),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_6),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_6),
.A2(n_23),
.B1(n_26),
.B2(n_60),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_6),
.A2(n_60),
.B1(n_71),
.B2(n_72),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_6),
.A2(n_50),
.B1(n_52),
.B2(n_60),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_7),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_7),
.A2(n_17),
.B1(n_23),
.B2(n_26),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_7),
.A2(n_17),
.B1(n_50),
.B2(n_52),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_7),
.A2(n_17),
.B1(n_71),
.B2(n_72),
.Y(n_209)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_8),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_10),
.A2(n_23),
.B1(n_26),
.B2(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_11),
.A2(n_18),
.B1(n_19),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_11),
.A2(n_23),
.B1(n_26),
.B2(n_44),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_23),
.B(n_25),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_11),
.A2(n_44),
.B1(n_71),
.B2(n_72),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_11),
.A2(n_44),
.B1(n_50),
.B2(n_52),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_11),
.B(n_22),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_11),
.A2(n_50),
.B(n_149),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g171 ( 
.A1(n_11),
.A2(n_68),
.B(n_72),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_11),
.B(n_49),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_36),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_34),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_29),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_20),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_16),
.A2(n_22),
.B1(n_27),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_18),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_19),
.B1(n_24),
.B2(n_25),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_18),
.A2(n_24),
.B(n_44),
.C(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_21),
.B(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_22),
.A2(n_27),
.B1(n_43),
.B2(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx5_ASAP7_75t_SL g26 ( 
.A(n_23),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_23),
.A2(n_44),
.B(n_51),
.C(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_30),
.B(n_38),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_41),
.B(n_42),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_75),
.B(n_284),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_39),
.B(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_39),
.B(n_282),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_45),
.CI(n_56),
.CON(n_39),
.SN(n_39)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_41),
.A2(n_42),
.B(n_59),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_43),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_44),
.A2(n_50),
.B(n_69),
.C(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_44),
.B(n_102),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_44),
.B(n_70),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_49),
.B1(n_53),
.B2(n_62),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_48),
.B(n_87),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_49),
.A2(n_62),
.B(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_50),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_52),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_88),
.Y(n_107)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_55),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.C(n_63),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_84),
.B1(n_90),
.B2(n_91),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_57),
.B(n_91),
.C(n_92),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_57),
.A2(n_90),
.B1(n_106),
.B2(n_130),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_57),
.B(n_130),
.C(n_225),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_57),
.A2(n_90),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_61),
.A2(n_63),
.B1(n_263),
.B2(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_61),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_63),
.A2(n_260),
.B1(n_261),
.B2(n_263),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_63),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_74),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_70),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_111),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_66),
.A2(n_70),
.B1(n_111),
.B2(n_118),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_66),
.A2(n_70),
.B1(n_74),
.B2(n_230),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_70),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_71),
.B(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_99),
.Y(n_98)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_281),
.B(n_283),
.Y(n_75)
);

OAI321xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_255),
.A3(n_274),
.B1(n_279),
.B2(n_280),
.C(n_286),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_238),
.B(n_254),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_219),
.B(n_237),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_141),
.B(n_202),
.C(n_218),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_127),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_81),
.B(n_127),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_103),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_82),
.B(n_104),
.C(n_114),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_92),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_84),
.B(n_136),
.C(n_139),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_84),
.A2(n_91),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_84),
.A2(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_84),
.B(n_244),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_89),
.B(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_96),
.A2(n_134),
.B1(n_173),
.B2(n_176),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_96),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_96),
.B(n_186),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_96),
.B(n_163),
.C(n_175),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_124),
.B(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_98),
.B(n_99),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_98),
.A2(n_102),
.B1(n_123),
.B2(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_113),
.B2(n_114),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.C(n_112),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_108),
.B1(n_109),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_106),
.A2(n_115),
.B1(n_116),
.B2(n_130),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_107),
.Y(n_262)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_112),
.A2(n_131),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_112),
.A2(n_131),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_112),
.A2(n_131),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_112),
.B(n_261),
.C(n_263),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_112),
.B(n_268),
.C(n_273),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_121),
.B2(n_122),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_115),
.A2(n_116),
.B1(n_170),
.B2(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_115),
.B(n_122),
.Y(n_212)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_130),
.C(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_116),
.B(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_119),
.B(n_120),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_120),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_133),
.C(n_135),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_128),
.B(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_129),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_131),
.B(n_212),
.C(n_214),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_133),
.B(n_135),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_139),
.B1(n_140),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_136),
.B(n_183),
.Y(n_182)
);

INVx5_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_201),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_196),
.B(n_200),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_166),
.B(n_195),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_154),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_145),
.B(n_154),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_150),
.B1(n_151),
.B2(n_153),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_147),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_153),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_152),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_160),
.B2(n_161),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_163),
.C(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_157),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_158),
.B(n_179),
.Y(n_188)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_162),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_163),
.A2(n_165),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_163),
.A2(n_165),
.B1(n_208),
.B2(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_163),
.B(n_208),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_190),
.B(n_194),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_177),
.B(n_189),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_172),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_170),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_174),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_181),
.B(n_188),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_185),
.B(n_187),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_192),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_198),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_203),
.B(n_204),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_216),
.B2(n_217),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_211),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_211),
.C(n_217),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_208),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_216),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_221),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_236),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_227),
.B2(n_228),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_228),
.C(n_236),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_232),
.B1(n_233),
.B2(n_235),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_229),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_233),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_233),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_L g265 ( 
.A1(n_233),
.A2(n_247),
.B(n_249),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_239),
.B(n_240),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_252),
.B2(n_253),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_246),
.C(n_253),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_257),
.C(n_264),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_257),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_252),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_266),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_266),
.Y(n_280)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_264),
.A2(n_265),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_273),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_276),
.Y(n_279)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);


endmodule