module real_jpeg_16939_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_620;
wire n_578;
wire n_332;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_469;
wire n_98;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_594;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_572;
wire n_155;
wire n_586;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_0),
.A2(n_21),
.B(n_632),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_0),
.B(n_633),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_1),
.A2(n_59),
.B1(n_63),
.B2(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_1),
.A2(n_63),
.B1(n_146),
.B2(n_152),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_1),
.A2(n_63),
.B1(n_289),
.B2(n_293),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_2),
.B(n_162),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_2),
.A2(n_211),
.B(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_2),
.Y(n_378)
);

OAI32xp33_ASAP7_75t_L g453 ( 
.A1(n_2),
.A2(n_454),
.A3(n_457),
.B1(n_460),
.B2(n_465),
.Y(n_453)
);

OAI32xp33_ASAP7_75t_L g489 ( 
.A1(n_2),
.A2(n_454),
.A3(n_457),
.B1(n_460),
.B2(n_465),
.Y(n_489)
);

OAI32xp33_ASAP7_75t_L g491 ( 
.A1(n_2),
.A2(n_454),
.A3(n_457),
.B1(n_460),
.B2(n_465),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_SL g501 ( 
.A1(n_2),
.A2(n_378),
.B1(n_502),
.B2(n_505),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_2),
.B(n_55),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_2),
.A2(n_217),
.B1(n_480),
.B2(n_590),
.Y(n_589)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_3),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_3),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_3),
.A2(n_88),
.B1(n_187),
.B2(n_312),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_3),
.A2(n_187),
.B1(n_446),
.B2(n_449),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_3),
.A2(n_187),
.B1(n_373),
.B2(n_525),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_4),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_4),
.Y(n_232)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_4),
.Y(n_308)
);

BUFx5_ASAP7_75t_L g395 ( 
.A(n_4),
.Y(n_395)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_5),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_5),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_6),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_6),
.A2(n_102),
.B1(n_107),
.B2(n_110),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_6),
.A2(n_102),
.B1(n_280),
.B2(n_282),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_6),
.A2(n_102),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_7),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_7),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_7),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_8),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_8),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_8),
.A2(n_196),
.B1(n_343),
.B2(n_346),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_8),
.A2(n_115),
.B1(n_196),
.B2(n_401),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_8),
.A2(n_196),
.B1(n_469),
.B2(n_474),
.Y(n_468)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_9),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_10),
.A2(n_246),
.B1(n_248),
.B2(n_250),
.Y(n_245)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_10),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_10),
.A2(n_250),
.B1(n_361),
.B2(n_366),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_10),
.A2(n_250),
.B1(n_517),
.B2(n_521),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_SL g590 ( 
.A1(n_10),
.A2(n_250),
.B1(n_584),
.B2(n_591),
.Y(n_590)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_11),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_11),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_11),
.Y(n_222)
);

BUFx4f_ASAP7_75t_L g473 ( 
.A(n_11),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_12),
.A2(n_115),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_12),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_12),
.A2(n_107),
.B1(n_252),
.B2(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_12),
.A2(n_252),
.B1(n_494),
.B2(n_497),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_SL g571 ( 
.A1(n_12),
.A2(n_252),
.B1(n_572),
.B2(n_576),
.Y(n_571)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_13),
.A2(n_87),
.B1(n_91),
.B2(n_92),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_13),
.A2(n_91),
.B1(n_110),
.B2(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_13),
.A2(n_91),
.B1(n_234),
.B2(n_239),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_13),
.A2(n_91),
.B1(n_260),
.B2(n_263),
.Y(n_259)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_15),
.A2(n_115),
.B1(n_117),
.B2(n_119),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_15),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_15),
.A2(n_119),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_15),
.A2(n_119),
.B1(n_270),
.B2(n_274),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_15),
.A2(n_119),
.B1(n_404),
.B2(n_407),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_16),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_16),
.Y(n_262)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_16),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_16),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_16),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_17),
.A2(n_162),
.B1(n_164),
.B2(n_167),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_17),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_17),
.A2(n_167),
.B1(n_270),
.B2(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_17),
.A2(n_64),
.B1(n_167),
.B2(n_316),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_17),
.A2(n_167),
.B1(n_373),
.B2(n_374),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_19),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_19),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_177),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_176),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_155),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_25),
.B(n_155),
.Y(n_176)
);

BUFx24_ASAP7_75t_SL g634 ( 
.A(n_25),
.Y(n_634)
);

FAx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_68),
.CI(n_103),
.CON(n_25),
.SN(n_25)
);

OAI21xp33_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_55),
.B(n_57),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g111 ( 
.A(n_27),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_27),
.A2(n_55),
.B1(n_185),
.B2(n_192),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_27),
.A2(n_55),
.B1(n_420),
.B2(n_421),
.Y(n_419)
);

OA21x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_37),
.B(n_43),
.Y(n_27)
);

INVxp33_ASAP7_75t_L g465 ( 
.A(n_28),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_35),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_36),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_36),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_41),
.Y(n_174)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B1(n_49),
.B2(n_52),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_47),
.Y(n_388)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_48),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g275 ( 
.A(n_48),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_48),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_48),
.Y(n_448)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_51),
.Y(n_139)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_51),
.Y(n_151)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_56),
.A2(n_58),
.B1(n_106),
.B2(n_111),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_56),
.A2(n_106),
.B1(n_111),
.B2(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_56),
.A2(n_111),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_56),
.A2(n_111),
.B1(n_328),
.B2(n_334),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_L g359 ( 
.A1(n_56),
.A2(n_111),
.B1(n_328),
.B2(n_360),
.Y(n_359)
);

OAI22x1_ASAP7_75t_L g402 ( 
.A1(n_56),
.A2(n_111),
.B1(n_315),
.B2(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_56),
.A2(n_111),
.B1(n_360),
.B2(n_501),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_67),
.Y(n_333)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_67),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_85),
.B1(n_97),
.B2(n_98),
.Y(n_68)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_69),
.A2(n_97),
.B1(n_114),
.B2(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_69),
.A2(n_97),
.B1(n_245),
.B2(n_251),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_69),
.A2(n_97),
.B1(n_251),
.B2(n_311),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_69),
.A2(n_97),
.B1(n_245),
.B2(n_336),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_69),
.A2(n_97),
.B1(n_311),
.B2(n_400),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_69),
.A2(n_97),
.B1(n_161),
.B2(n_400),
.Y(n_429)
);

AO21x2_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_76),
.B(n_80),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_76),
.A2(n_201),
.B1(n_210),
.B2(n_212),
.Y(n_200)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AO22x2_ASAP7_75t_L g80 ( 
.A1(n_78),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_80),
.A2(n_86),
.B1(n_113),
.B2(n_120),
.Y(n_112)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_81),
.Y(n_198)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_82),
.Y(n_409)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_90),
.Y(n_247)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2x1_ASAP7_75t_R g377 ( 
.A(n_97),
.B(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_112),
.C(n_121),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_104),
.A2(n_105),
.B1(n_121),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_109),
.Y(n_318)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_109),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_115),
.Y(n_253)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_121),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_121),
.B(n_170),
.C(n_175),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_121),
.B(n_170),
.Y(n_619)
);

OA21x2_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_136),
.B(n_145),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_122),
.B(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_122),
.A2(n_136),
.B1(n_269),
.B2(n_298),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_122),
.A2(n_136),
.B1(n_145),
.B2(n_423),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_122),
.A2(n_136),
.B1(n_445),
.B2(n_493),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_122),
.A2(n_136),
.B1(n_493),
.B2(n_516),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_122),
.A2(n_136),
.B1(n_516),
.B2(n_561),
.Y(n_560)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_123),
.A2(n_341),
.B1(n_342),
.B2(n_350),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_123),
.A2(n_259),
.B1(n_341),
.B2(n_387),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_123),
.A2(n_341),
.B1(n_342),
.B2(n_444),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_123),
.B(n_378),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_128),
.B1(n_132),
.B2(n_134),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_126),
.Y(n_549)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_129),
.Y(n_228)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_130),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_130),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_131),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_133),
.Y(n_292)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_136),
.B(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_136),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_144),
.Y(n_522)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_151),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_151),
.Y(n_496)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_151),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_154),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.C(n_168),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_157),
.A2(n_160),
.B1(n_175),
.B2(n_628),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_157),
.Y(n_628)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_160),
.A2(n_175),
.B1(n_619),
.B2(n_620),
.Y(n_618)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_164),
.Y(n_339)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_165),
.Y(n_401)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_166),
.Y(n_312)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_169),
.B(n_627),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_171),
.Y(n_421)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_609),
.B(n_629),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_434),
.B(n_604),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_379),
.C(n_414),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_319),
.B(n_351),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_182),
.B(n_319),
.C(n_606),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_254),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_183),
.B(n_255),
.C(n_294),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_199),
.C(n_243),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_184),
.A2(n_243),
.B1(n_244),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_184),
.Y(n_322)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_185),
.Y(n_334)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_192),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_195),
.Y(n_365)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_195),
.Y(n_510)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_199),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_216),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_200),
.B(n_216),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_206),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_223),
.B1(n_229),
.B2(n_233),
.Y(n_216)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_217),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_217),
.A2(n_233),
.B1(n_279),
.B2(n_304),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_217),
.A2(n_288),
.B(n_393),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_217),
.A2(n_524),
.B1(n_528),
.B2(n_532),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_217),
.A2(n_571),
.B1(n_590),
.B2(n_594),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

INVx5_ASAP7_75t_L g480 ( 
.A(n_218),
.Y(n_480)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_220),
.Y(n_376)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_221),
.Y(n_293)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_222),
.Y(n_281)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_222),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g223 ( 
.A(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_224),
.A2(n_277),
.B1(n_372),
.B2(n_376),
.Y(n_371)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_228),
.Y(n_375)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_239),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_294),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_276),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_268),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_257),
.A2(n_268),
.B(n_276),
.Y(n_410)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_261),
.Y(n_498)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_262),
.Y(n_450)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_266),
.Y(n_349)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_267),
.Y(n_273)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_267),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_267),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_270),
.B(n_378),
.Y(n_550)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_284),
.B2(n_287),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_277),
.A2(n_372),
.B1(n_468),
.B2(n_478),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_277),
.A2(n_478),
.B1(n_570),
.B2(n_578),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_281),
.Y(n_547)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_290),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_292),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_309),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_295),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_303),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_296),
.A2(n_297),
.B1(n_303),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_298),
.Y(n_350)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_303),
.Y(n_325)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_307),
.Y(n_531)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_307),
.Y(n_596)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_313),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_310),
.B(n_382),
.C(n_383),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_313),
.Y(n_383)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_323),
.C(n_326),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_320),
.B(n_353),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_326),
.Y(n_353)
);

MAJx2_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_335),
.C(n_340),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_340),
.Y(n_356)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_333),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_335),
.B(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_354),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_352),
.B(n_354),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_357),
.C(n_358),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_355),
.B(n_437),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_357),
.B(n_358),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_370),
.C(n_377),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_359),
.B(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_370),
.A2(n_371),
.B1(n_377),
.B2(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_377),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_378),
.B(n_461),
.Y(n_460)
);

OAI21xp33_ASAP7_75t_SL g561 ( 
.A1(n_378),
.A2(n_550),
.B(n_562),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_378),
.B(n_586),
.Y(n_585)
);

A2O1A1O1Ixp25_ASAP7_75t_L g604 ( 
.A1(n_379),
.A2(n_414),
.B(n_605),
.C(n_607),
.D(n_608),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_413),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_380),
.B(n_413),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_381),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_397),
.B1(n_411),
.B2(n_412),
.Y(n_384)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_385),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_385),
.B(n_412),
.C(n_433),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_386),
.A2(n_391),
.B1(n_392),
.B2(n_396),
.Y(n_385)
);

INVxp33_ASAP7_75t_SL g396 ( 
.A(n_386),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_386),
.B(n_392),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_387),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_391),
.A2(n_392),
.B1(n_428),
.B2(n_429),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_391),
.A2(n_429),
.B(n_431),
.Y(n_616)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx12f_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_410),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_402),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_399),
.B(n_402),
.C(n_410),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_403),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_415),
.B(n_432),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_415),
.B(n_432),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_416),
.B(n_613),
.C(n_614),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_425),
.Y(n_417)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_418),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_419),
.A2(n_422),
.B(n_424),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_419),
.B(n_422),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_424),
.B(n_618),
.Y(n_617)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_424),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_425),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_426),
.A2(n_427),
.B1(n_430),
.B2(n_431),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_430),
.Y(n_431)
);

AOI21x1_ASAP7_75t_L g434 ( 
.A1(n_435),
.A2(n_481),
.B(n_603),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_436),
.B(n_438),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_436),
.B(n_438),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_443),
.C(n_451),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_439),
.A2(n_440),
.B1(n_484),
.B2(n_485),
.Y(n_483)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_443),
.A2(n_451),
.B1(n_452),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_443),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_466),
.Y(n_452)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_466),
.A2(n_467),
.B1(n_489),
.B2(n_490),
.Y(n_488)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_468),
.Y(n_532)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_473),
.Y(n_577)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_477),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_482),
.A2(n_511),
.B(n_602),
.Y(n_481)
);

NOR2xp67_ASAP7_75t_SL g482 ( 
.A(n_483),
.B(n_487),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_483),
.B(n_487),
.Y(n_602)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_492),
.C(n_499),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_488),
.B(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_492),
.A2(n_499),
.B1(n_500),
.B2(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_492),
.Y(n_537)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

AOI21x1_ASAP7_75t_SL g511 ( 
.A1(n_512),
.A2(n_538),
.B(n_601),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_SL g512 ( 
.A(n_513),
.B(n_535),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_513),
.B(n_535),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_523),
.C(n_533),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_514),
.A2(n_515),
.B1(n_533),
.B2(n_534),
.Y(n_566)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_523),
.B(n_566),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_524),
.Y(n_578)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx4_ASAP7_75t_SL g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_531),
.Y(n_588)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_539),
.A2(n_567),
.B(n_600),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_565),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_540),
.B(n_565),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_559),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_541),
.A2(n_559),
.B1(n_560),
.B2(n_580),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

OAI32xp33_ASAP7_75t_L g541 ( 
.A1(n_542),
.A2(n_545),
.A3(n_548),
.B1(n_550),
.B2(n_551),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_552),
.B(n_556),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx8_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_568),
.A2(n_581),
.B(n_599),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_569),
.B(n_579),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_569),
.B(n_579),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_572),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_574),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_582),
.A2(n_592),
.B(n_598),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_583),
.B(n_589),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_584),
.B(n_585),
.Y(n_583)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_593),
.B(n_597),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_593),
.B(n_597),
.Y(n_598)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_611),
.B(n_621),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_612),
.B(n_615),
.Y(n_611)
);

NAND2x1p5_ASAP7_75t_L g630 ( 
.A(n_612),
.B(n_615),
.Y(n_630)
);

XOR2x2_ASAP7_75t_SL g615 ( 
.A(n_616),
.B(n_617),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_616),
.B(n_624),
.C(n_625),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_618),
.Y(n_624)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_619),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

OAI21x1_ASAP7_75t_SL g629 ( 
.A1(n_622),
.A2(n_630),
.B(n_631),
.Y(n_629)
);

NOR2xp67_ASAP7_75t_L g622 ( 
.A(n_623),
.B(n_626),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_623),
.B(n_626),
.Y(n_631)
);


endmodule