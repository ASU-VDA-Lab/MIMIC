module fake_ariane_100_n_120 (n_8, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_50, n_38, n_2, n_47, n_18, n_32, n_28, n_37, n_9, n_51, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_52, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_53, n_21, n_23, n_35, n_10, n_25, n_120);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_51;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_52;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_53;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_120;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_119;
wire n_90;
wire n_110;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_106;
wire n_111;
wire n_115;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_100;
wire n_62;
wire n_76;
wire n_103;
wire n_79;
wire n_84;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_82;
wire n_57;
wire n_70;
wire n_117;
wire n_85;
wire n_94;
wire n_101;
wire n_58;
wire n_65;
wire n_112;
wire n_73;
wire n_77;
wire n_118;
wire n_93;
wire n_61;
wire n_108;
wire n_102;
wire n_81;
wire n_87;
wire n_55;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_116;
wire n_104;
wire n_78;
wire n_63;
wire n_59;
wire n_99;
wire n_54;

INVx2_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_25),
.B(n_6),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_8),
.B(n_4),
.Y(n_59)
);

AND2x4_ASAP7_75t_L g60 ( 
.A(n_0),
.B(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_12),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_29),
.B1(n_52),
.B2(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_14),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

OAI21x1_ASAP7_75t_L g70 ( 
.A1(n_27),
.A2(n_34),
.B(n_36),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_30),
.B(n_18),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_7),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_32),
.B(n_2),
.Y(n_84)
);

BUFx4f_ASAP7_75t_SL g85 ( 
.A(n_64),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_65),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_55),
.B(n_0),
.Y(n_87)
);

OR2x6_ASAP7_75t_SL g88 ( 
.A(n_54),
.B(n_5),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_17),
.B(n_20),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_21),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_23),
.Y(n_95)
);

OAI21x1_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_61),
.B(n_76),
.Y(n_96)
);

AOI222xp33_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_62),
.B1(n_60),
.B2(n_81),
.C1(n_80),
.C2(n_79),
.Y(n_97)
);

OAI21x1_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_77),
.B(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

OAI21x1_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_69),
.B(n_74),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_91),
.B(n_92),
.C(n_73),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_59),
.B1(n_57),
.B2(n_78),
.Y(n_102)
);

NAND2x1p5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_94),
.Y(n_103)
);

OAI21x1_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_78),
.B(n_72),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_85),
.B1(n_72),
.B2(n_93),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_93),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_111),
.A2(n_106),
.B1(n_108),
.B2(n_102),
.Y(n_113)
);

OAI211xp5_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_107),
.B(n_101),
.C(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_109),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_114),
.A2(n_110),
.B1(n_93),
.B2(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_24),
.Y(n_117)
);

NAND4xp75_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_116),
.C(n_33),
.D(n_35),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_31),
.B1(n_38),
.B2(n_41),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_119),
.A2(n_45),
.B1(n_49),
.B2(n_51),
.Y(n_120)
);


endmodule