module fake_netlist_6_1177_n_1728 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1728);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1728;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_33),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_32),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_18),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_119),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_138),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_120),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_151),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_56),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_55),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_45),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_85),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_73),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_29),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_18),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_98),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_55),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_26),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_70),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_32),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_51),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_4),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_115),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_125),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_41),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_40),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_105),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_91),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_21),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_83),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_23),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_30),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_124),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_22),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_54),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_82),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_46),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_66),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_87),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_110),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_34),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_92),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_45),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_94),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_84),
.Y(n_204)
);

INVxp67_ASAP7_75t_SL g205 ( 
.A(n_78),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_20),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_142),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_7),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_52),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_16),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_102),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_53),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_81),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_23),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_50),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_63),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_17),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_33),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_26),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_58),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_71),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_51),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_30),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_16),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_21),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_44),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_19),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_93),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_34),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_53),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_146),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_107),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_5),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_20),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_46),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_145),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_61),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_13),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_132),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_67),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_13),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_126),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_79),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_15),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_108),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_49),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_89),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_80),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_74),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_64),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_114),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_149),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_38),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_22),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_72),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_9),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_17),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_99),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_109),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_130),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_39),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_10),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_88),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_148),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_144),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_101),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_4),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_97),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_19),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_6),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_7),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_122),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_35),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_60),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_54),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_77),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_96),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_143),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_27),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_44),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_103),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_100),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_1),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_40),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_36),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_141),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_14),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_86),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_48),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_59),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_75),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_48),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_62),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_24),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_139),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_10),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_106),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_3),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_43),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_36),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_49),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_29),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_8),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_150),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_24),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_57),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_140),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_156),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_202),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_R g310 ( 
.A(n_284),
.B(n_147),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_246),
.B(n_0),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_156),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_218),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_157),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_158),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_170),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_218),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_218),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_204),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_0),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_218),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_174),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_300),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_159),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_218),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_202),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_160),
.Y(n_327)
);

INVxp33_ASAP7_75t_SL g328 ( 
.A(n_306),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_232),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_202),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_174),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_161),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_206),
.B(n_1),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_155),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_194),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_268),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_288),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_281),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_165),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_169),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_155),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_171),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_181),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_182),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_194),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_167),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_188),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_195),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_197),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_304),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_224),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_199),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_167),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_292),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_288),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_224),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_248),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_203),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_235),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_207),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_216),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_220),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_221),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_235),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_253),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_228),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_168),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_231),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_237),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_166),
.B(n_2),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_253),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_168),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_240),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_250),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_175),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_175),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_178),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_292),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_178),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_251),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_179),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_252),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_179),
.Y(n_383)
);

NOR2x1_ASAP7_75t_L g384 ( 
.A(n_313),
.B(n_245),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_313),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_314),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_317),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_309),
.B(n_307),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_309),
.B(n_255),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_326),
.B(n_245),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_317),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_318),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_318),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_316),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_308),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_321),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_316),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_321),
.B(n_259),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_325),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_308),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_337),
.B(n_323),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_316),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_325),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_330),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_330),
.B(n_260),
.Y(n_407)
);

BUFx8_ASAP7_75t_L g408 ( 
.A(n_378),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_315),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_345),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_334),
.B(n_261),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_375),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_334),
.B(n_261),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_341),
.B(n_153),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_375),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_376),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_331),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_354),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_320),
.B(n_189),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_345),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_377),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_351),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_378),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_328),
.B(n_185),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_379),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_351),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_341),
.B(n_263),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_346),
.B(n_265),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_379),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_381),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_346),
.B(n_302),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_353),
.B(n_153),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_370),
.B(n_242),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_381),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_353),
.B(n_173),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_356),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_383),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_383),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_367),
.B(n_266),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_324),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_355),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_367),
.B(n_272),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_356),
.Y(n_446)
);

AND2x6_ASAP7_75t_L g447 ( 
.A(n_333),
.B(n_173),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_312),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_359),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_372),
.B(n_198),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_312),
.Y(n_451)
);

BUFx8_ASAP7_75t_L g452 ( 
.A(n_337),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_385),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_327),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_395),
.B(n_322),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_332),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_385),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_412),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_393),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_390),
.Y(n_460)
);

INVx4_ASAP7_75t_SL g461 ( 
.A(n_447),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_393),
.Y(n_462)
);

OAI22xp33_ASAP7_75t_L g463 ( 
.A1(n_421),
.A2(n_322),
.B1(n_333),
.B2(n_162),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_447),
.A2(n_238),
.B1(n_206),
.B2(n_241),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_394),
.Y(n_465)
);

BUFx8_ASAP7_75t_SL g466 ( 
.A(n_444),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_388),
.B(n_339),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_310),
.Y(n_468)
);

OR2x6_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_166),
.Y(n_469)
);

INVx5_ASAP7_75t_L g470 ( 
.A(n_447),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_393),
.Y(n_471)
);

OR2x6_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_172),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_387),
.Y(n_473)
);

CKINVDCx12_ASAP7_75t_R g474 ( 
.A(n_412),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_390),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_388),
.B(n_340),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_447),
.A2(n_435),
.B1(n_438),
.B2(n_415),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_415),
.B(n_372),
.Y(n_478)
);

BUFx16f_ASAP7_75t_R g479 ( 
.A(n_452),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_396),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_452),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_387),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_389),
.B(n_342),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_396),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_391),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_452),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_415),
.B(n_359),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_390),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_396),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_389),
.B(n_343),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_392),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_392),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_421),
.A2(n_275),
.B1(n_190),
.B2(n_283),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_394),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_386),
.B(n_357),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_399),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_427),
.B(n_344),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_427),
.B(n_347),
.Y(n_499)
);

AND3x1_ASAP7_75t_L g500 ( 
.A(n_395),
.B(n_241),
.C(n_238),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_400),
.B(n_348),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_400),
.B(n_349),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_394),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_403),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_403),
.Y(n_505)
);

HB1xp67_ASAP7_75t_SL g506 ( 
.A(n_452),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_415),
.B(n_364),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_394),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_413),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_408),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_410),
.B(n_352),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_399),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_415),
.B(n_364),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_410),
.B(n_358),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_430),
.B(n_360),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_390),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_398),
.B(n_362),
.Y(n_517)
);

OR2x6_ASAP7_75t_L g518 ( 
.A(n_443),
.B(n_172),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_413),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_435),
.B(n_365),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_399),
.Y(n_521)
);

BUFx8_ASAP7_75t_SL g522 ( 
.A(n_444),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_412),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_398),
.B(n_363),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_452),
.Y(n_525)
);

NAND2xp33_ASAP7_75t_SL g526 ( 
.A(n_448),
.B(n_361),
.Y(n_526)
);

INVx4_ASAP7_75t_L g527 ( 
.A(n_394),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_390),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_410),
.B(n_366),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_435),
.B(n_368),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_416),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_435),
.B(n_369),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_435),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_394),
.Y(n_534)
);

AND2x2_ASAP7_75t_SL g535 ( 
.A(n_438),
.B(n_198),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_438),
.B(n_373),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_416),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_438),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_410),
.B(n_374),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_438),
.B(n_380),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_410),
.B(n_382),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_430),
.B(n_213),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_417),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_417),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_431),
.B(n_213),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_420),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_394),
.Y(n_547)
);

OR2x6_ASAP7_75t_L g548 ( 
.A(n_450),
.B(n_407),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_450),
.B(n_365),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_397),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_420),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_423),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_450),
.B(n_243),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_423),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_431),
.B(n_319),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_425),
.Y(n_556)
);

AND3x2_ASAP7_75t_L g557 ( 
.A(n_448),
.B(n_177),
.C(n_176),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_397),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_397),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_442),
.B(n_329),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_397),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_450),
.B(n_274),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_425),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_447),
.A2(n_302),
.B1(n_303),
.B2(n_180),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_397),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_450),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_428),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_397),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_397),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_447),
.A2(n_180),
.B1(n_303),
.B2(n_301),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_426),
.B(n_371),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_447),
.A2(n_183),
.B1(n_301),
.B2(n_191),
.Y(n_572)
);

INVx6_ASAP7_75t_L g573 ( 
.A(n_402),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_414),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_402),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_414),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_447),
.A2(n_183),
.B1(n_191),
.B2(n_296),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_402),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_442),
.B(n_278),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_445),
.B(n_290),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_408),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_414),
.A2(n_193),
.B1(n_209),
.B2(n_296),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_402),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_426),
.A2(n_200),
.B1(n_212),
.B2(n_210),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_445),
.B(n_213),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_402),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_401),
.A2(n_208),
.B1(n_233),
.B2(n_230),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_402),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_402),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_428),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_407),
.B(n_336),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_434),
.B(n_291),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_432),
.Y(n_593)
);

BUFx6f_ASAP7_75t_SL g594 ( 
.A(n_432),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_433),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_434),
.B(n_384),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_433),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_437),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_437),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_405),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_434),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_L g602 ( 
.A(n_451),
.B(n_187),
.C(n_305),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_535),
.B(n_515),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g604 ( 
.A(n_510),
.B(n_408),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_454),
.B(n_451),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_535),
.B(n_405),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_535),
.A2(n_217),
.B1(n_254),
.B2(n_234),
.Y(n_607)
);

AND3x4_ASAP7_75t_L g608 ( 
.A(n_601),
.B(n_311),
.C(n_338),
.Y(n_608)
);

AND2x2_ASAP7_75t_SL g609 ( 
.A(n_477),
.B(n_176),
.Y(n_609)
);

INVxp33_ASAP7_75t_L g610 ( 
.A(n_455),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_456),
.A2(n_350),
.B1(n_205),
.B2(n_295),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_458),
.B(n_418),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_458),
.B(n_405),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_533),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_533),
.Y(n_615)
);

BUFx8_ASAP7_75t_L g616 ( 
.A(n_510),
.Y(n_616)
);

A2O1A1Ixp33_ASAP7_75t_L g617 ( 
.A1(n_523),
.A2(n_576),
.B(n_574),
.C(n_538),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_523),
.B(n_408),
.Y(n_618)
);

O2A1O1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_574),
.A2(n_440),
.B(n_441),
.C(n_222),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_576),
.B(n_601),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_538),
.B(n_405),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_478),
.B(n_418),
.Y(n_622)
);

INVx6_ASAP7_75t_L g623 ( 
.A(n_488),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_488),
.B(n_440),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_459),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_459),
.Y(n_626)
);

O2A1O1Ixp33_ASAP7_75t_L g627 ( 
.A1(n_596),
.A2(n_441),
.B(n_222),
.C(n_270),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_566),
.B(n_405),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_460),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_474),
.A2(n_384),
.B1(n_408),
.B2(n_201),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_530),
.B(n_419),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_478),
.B(n_405),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_460),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_470),
.B(n_405),
.Y(n_634)
);

NOR3xp33_ASAP7_75t_L g635 ( 
.A(n_463),
.B(n_526),
.C(n_555),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_455),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_467),
.B(n_406),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_475),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_548),
.A2(n_258),
.B1(n_186),
.B2(n_177),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_475),
.Y(n_640)
);

NAND3xp33_ASAP7_75t_L g641 ( 
.A(n_494),
.B(n_592),
.C(n_602),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_501),
.B(n_419),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_481),
.B(n_213),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_489),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_571),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_489),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_476),
.B(n_483),
.Y(n_647)
);

NOR3xp33_ASAP7_75t_L g648 ( 
.A(n_560),
.B(n_196),
.C(n_184),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_491),
.B(n_406),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_516),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_474),
.A2(n_201),
.B1(n_186),
.B2(n_192),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_517),
.B(n_524),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_507),
.B(n_406),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_532),
.B(n_154),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_536),
.B(n_236),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_516),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_507),
.B(n_406),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_SL g658 ( 
.A1(n_494),
.A2(n_311),
.B1(n_164),
.B2(n_215),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_462),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_508),
.A2(n_449),
.B(n_409),
.Y(n_660)
);

NOR3xp33_ASAP7_75t_L g661 ( 
.A(n_591),
.B(n_163),
.C(n_256),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_462),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_540),
.B(n_219),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_470),
.B(n_406),
.Y(n_664)
);

OAI221xp5_ASAP7_75t_L g665 ( 
.A1(n_582),
.A2(n_193),
.B1(n_209),
.B2(n_214),
.C(n_217),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_528),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_513),
.B(n_406),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_513),
.B(n_520),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_471),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_L g670 ( 
.A(n_579),
.B(n_170),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_520),
.B(n_549),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_549),
.B(n_406),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_528),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_SL g674 ( 
.A1(n_539),
.A2(n_249),
.B1(n_236),
.B2(n_211),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_470),
.B(n_170),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_498),
.B(n_223),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_580),
.B(n_404),
.Y(n_677)
);

AND2x6_ASAP7_75t_L g678 ( 
.A(n_550),
.B(n_192),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_553),
.B(n_404),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_571),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_501),
.B(n_236),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_480),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_502),
.B(n_446),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_509),
.B(n_519),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_480),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_570),
.A2(n_271),
.B1(n_270),
.B2(n_279),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_509),
.B(n_404),
.Y(n_687)
);

NOR3xp33_ASAP7_75t_L g688 ( 
.A(n_499),
.B(n_225),
.C(n_226),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_484),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_502),
.B(n_227),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_519),
.Y(n_691)
);

OR2x6_ASAP7_75t_L g692 ( 
.A(n_469),
.B(n_472),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_531),
.B(n_404),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_531),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_548),
.A2(n_277),
.B1(n_247),
.B2(n_211),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_500),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_537),
.B(n_404),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_484),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_548),
.A2(n_562),
.B(n_468),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_542),
.B(n_545),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_572),
.A2(n_267),
.B1(n_214),
.B2(n_234),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_537),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_543),
.B(n_422),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_577),
.A2(n_279),
.B1(n_294),
.B2(n_271),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_548),
.A2(n_258),
.B1(n_264),
.B2(n_276),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_470),
.B(n_170),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_543),
.B(n_544),
.Y(n_707)
);

NOR2xp67_ASAP7_75t_L g708 ( 
.A(n_481),
.B(n_446),
.Y(n_708)
);

O2A1O1Ixp33_ASAP7_75t_L g709 ( 
.A1(n_585),
.A2(n_294),
.B(n_254),
.C(n_267),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_544),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_587),
.B(n_229),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_470),
.B(n_170),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_R g713 ( 
.A(n_581),
.B(n_244),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_548),
.A2(n_286),
.B1(n_282),
.B2(n_277),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_496),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_546),
.B(n_422),
.Y(n_716)
);

INVx5_ASAP7_75t_L g717 ( 
.A(n_534),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_511),
.B(n_236),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_490),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_514),
.B(n_257),
.Y(n_720)
);

AO22x2_ASAP7_75t_L g721 ( 
.A1(n_479),
.A2(n_239),
.B1(n_247),
.B2(n_264),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_529),
.B(n_262),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_546),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_541),
.B(n_269),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_551),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_551),
.B(n_552),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_552),
.B(n_422),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_550),
.A2(n_449),
.B(n_439),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_490),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_470),
.B(n_170),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_497),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_554),
.B(n_422),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_SL g733 ( 
.A(n_594),
.B(n_273),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_461),
.B(n_170),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_469),
.A2(n_297),
.B1(n_239),
.B2(n_276),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_584),
.B(n_371),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_469),
.A2(n_297),
.B1(n_282),
.B2(n_286),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_554),
.B(n_429),
.Y(n_738)
);

NAND3xp33_ASAP7_75t_L g739 ( 
.A(n_584),
.B(n_299),
.C(n_280),
.Y(n_739)
);

AND2x6_ASAP7_75t_SL g740 ( 
.A(n_469),
.B(n_285),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_556),
.B(n_249),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_557),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_556),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_563),
.B(n_422),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_497),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_469),
.A2(n_170),
.B1(n_249),
.B2(n_429),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_558),
.A2(n_429),
.B(n_439),
.Y(n_747)
);

OAI22xp33_ASAP7_75t_L g748 ( 
.A1(n_472),
.A2(n_287),
.B1(n_289),
.B2(n_298),
.Y(n_748)
);

BUFx2_ASAP7_75t_L g749 ( 
.A(n_466),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_563),
.B(n_429),
.Y(n_750)
);

AO22x1_ASAP7_75t_L g751 ( 
.A1(n_567),
.A2(n_249),
.B1(n_429),
.B2(n_439),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_522),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_567),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_590),
.B(n_424),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_564),
.A2(n_170),
.B1(n_411),
.B2(n_409),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_590),
.B(n_424),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_593),
.B(n_595),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_464),
.A2(n_449),
.B1(n_411),
.B2(n_409),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_593),
.B(n_424),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_472),
.Y(n_760)
);

BUFx8_ASAP7_75t_L g761 ( 
.A(n_594),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_595),
.B(n_424),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_461),
.B(n_424),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_597),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_597),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_598),
.B(n_424),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_461),
.B(n_424),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_512),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_598),
.B(n_411),
.Y(n_769)
);

INVx8_ASAP7_75t_L g770 ( 
.A(n_594),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_599),
.Y(n_771)
);

OR2x6_ASAP7_75t_L g772 ( 
.A(n_472),
.B(n_2),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_599),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_652),
.B(n_453),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_606),
.A2(n_559),
.B(n_527),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_603),
.B(n_607),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_605),
.B(n_726),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_694),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_632),
.A2(n_559),
.B(n_527),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_636),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_607),
.A2(n_472),
.B1(n_518),
.B2(n_506),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_699),
.A2(n_559),
.B(n_527),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_683),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_764),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_605),
.B(n_518),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_647),
.B(n_461),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_610),
.B(n_518),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_749),
.Y(n_788)
);

OAI321xp33_ASAP7_75t_L g789 ( 
.A1(n_773),
.A2(n_518),
.A3(n_482),
.B1(n_457),
.B2(n_453),
.C(n_485),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_637),
.A2(n_588),
.B(n_534),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_764),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_726),
.B(n_457),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_609),
.A2(n_773),
.B(n_711),
.C(n_757),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_757),
.B(n_473),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_680),
.Y(n_795)
);

AOI21xp33_ASAP7_75t_L g796 ( 
.A1(n_711),
.A2(n_518),
.B(n_581),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_694),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_609),
.B(n_473),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_646),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_702),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_702),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_SL g802 ( 
.A1(n_692),
.A2(n_588),
.B(n_600),
.Y(n_802)
);

AOI21x1_ASAP7_75t_L g803 ( 
.A1(n_634),
.A2(n_558),
.B(n_589),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_649),
.A2(n_588),
.B(n_547),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_623),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_623),
.Y(n_806)
);

AOI21x1_ASAP7_75t_L g807 ( 
.A1(n_664),
.A2(n_565),
.B(n_569),
.Y(n_807)
);

OAI21xp33_ASAP7_75t_L g808 ( 
.A1(n_612),
.A2(n_485),
.B(n_482),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_654),
.B(n_663),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_646),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_617),
.A2(n_575),
.B(n_569),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_679),
.A2(n_534),
.B(n_547),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_641),
.B(n_575),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_623),
.A2(n_492),
.B1(n_493),
.B2(n_504),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_654),
.B(n_486),
.Y(n_815)
);

AOI21xp33_ASAP7_75t_L g816 ( 
.A1(n_676),
.A2(n_505),
.B(n_486),
.Y(n_816)
);

AOI221xp5_ASAP7_75t_SL g817 ( 
.A1(n_665),
.A2(n_504),
.B1(n_505),
.B2(n_492),
.C(n_493),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_663),
.B(n_583),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_752),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_680),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_668),
.A2(n_583),
.B(n_586),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_624),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_624),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_760),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_622),
.B(n_487),
.Y(n_825)
);

BUFx12f_ASAP7_75t_L g826 ( 
.A(n_761),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_612),
.B(n_525),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_700),
.A2(n_573),
.B1(n_586),
.B2(n_578),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_691),
.B(n_465),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_710),
.B(n_465),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_614),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_653),
.A2(n_547),
.B(n_534),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_671),
.A2(n_465),
.B(n_586),
.Y(n_833)
);

O2A1O1Ixp5_ASAP7_75t_L g834 ( 
.A1(n_769),
.A2(n_512),
.B(n_521),
.C(n_503),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_631),
.B(n_521),
.C(n_578),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_747),
.A2(n_495),
.B(n_578),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_645),
.B(n_495),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_615),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_723),
.B(n_495),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_657),
.A2(n_561),
.B(n_547),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_667),
.A2(n_561),
.B(n_547),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_629),
.Y(n_842)
);

OAI21xp33_ASAP7_75t_L g843 ( 
.A1(n_676),
.A2(n_503),
.B(n_568),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_672),
.A2(n_561),
.B(n_534),
.Y(n_844)
);

NOR2x1_ASAP7_75t_L g845 ( 
.A(n_708),
.B(n_568),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_621),
.A2(n_561),
.B(n_600),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_677),
.A2(n_568),
.B(n_503),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_725),
.B(n_561),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_770),
.Y(n_849)
);

O2A1O1Ixp33_ASAP7_75t_SL g850 ( 
.A1(n_639),
.A2(n_8),
.B(n_9),
.C(n_11),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_717),
.A2(n_600),
.B(n_573),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_743),
.B(n_573),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_717),
.A2(n_573),
.B(n_68),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_620),
.B(n_65),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_717),
.A2(n_136),
.B(n_128),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_633),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_631),
.B(n_11),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_717),
.A2(n_127),
.B(n_123),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_635),
.A2(n_121),
.B1(n_117),
.B2(n_116),
.Y(n_859)
);

NOR2xp67_ASAP7_75t_L g860 ( 
.A(n_700),
.B(n_113),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_628),
.A2(n_112),
.B(n_111),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_720),
.A2(n_12),
.B(n_14),
.C(n_15),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_753),
.B(n_12),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_765),
.B(n_25),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_720),
.A2(n_25),
.B(n_27),
.C(n_28),
.Y(n_865)
);

BUFx4f_ASAP7_75t_L g866 ( 
.A(n_770),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_692),
.Y(n_867)
);

A2O1A1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_722),
.A2(n_28),
.B(n_31),
.C(n_35),
.Y(n_868)
);

OAI321xp33_ASAP7_75t_L g869 ( 
.A1(n_748),
.A2(n_31),
.A3(n_37),
.B1(n_38),
.B2(n_39),
.C(n_41),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_692),
.A2(n_104),
.B1(n_95),
.B2(n_90),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_722),
.A2(n_37),
.B(n_42),
.C(n_43),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_771),
.B(n_42),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_684),
.B(n_707),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_736),
.B(n_47),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_638),
.B(n_47),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_640),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_644),
.B(n_69),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_650),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_613),
.A2(n_76),
.B(n_52),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_656),
.B(n_50),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_666),
.A2(n_56),
.B1(n_57),
.B2(n_673),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_690),
.B(n_724),
.Y(n_882)
);

BUFx8_ASAP7_75t_L g883 ( 
.A(n_642),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_664),
.A2(n_693),
.B(n_716),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_696),
.B(n_690),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_715),
.B(n_611),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_687),
.A2(n_744),
.B(n_738),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_724),
.A2(n_714),
.B(n_619),
.C(n_709),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_648),
.B(n_661),
.Y(n_889)
);

INVx4_ASAP7_75t_L g890 ( 
.A(n_770),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_748),
.B(n_697),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_761),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_742),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_772),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_625),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_703),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_727),
.A2(n_750),
.B(n_732),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_626),
.B(n_689),
.Y(n_898)
);

OAI21xp33_ASAP7_75t_L g899 ( 
.A1(n_674),
.A2(n_739),
.B(n_643),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_754),
.A2(n_762),
.B(n_766),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_659),
.B(n_662),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_686),
.A2(n_701),
.B(n_704),
.C(n_627),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_669),
.B(n_719),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_713),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_682),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_756),
.A2(n_767),
.B(n_763),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_681),
.B(n_713),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_735),
.A2(n_737),
.B1(n_686),
.B2(n_701),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_685),
.B(n_698),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_729),
.B(n_745),
.Y(n_910)
);

AOI21xp33_ASAP7_75t_L g911 ( 
.A1(n_695),
.A2(n_705),
.B(n_718),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_731),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_618),
.B(n_655),
.Y(n_913)
);

AND2x2_ASAP7_75t_SL g914 ( 
.A(n_604),
.B(n_704),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_768),
.Y(n_915)
);

OAI21xp33_ASAP7_75t_L g916 ( 
.A1(n_651),
.A2(n_688),
.B(n_741),
.Y(n_916)
);

AO22x1_ASAP7_75t_L g917 ( 
.A1(n_608),
.A2(n_616),
.B1(n_678),
.B2(n_772),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_763),
.A2(n_767),
.B(n_670),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_734),
.A2(n_660),
.B(n_759),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_675),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_746),
.A2(n_630),
.B(n_733),
.C(n_728),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_675),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_678),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_678),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_751),
.B(n_758),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_678),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_678),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_758),
.A2(n_755),
.B(n_734),
.C(n_712),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_772),
.A2(n_755),
.B1(n_608),
.B2(n_706),
.Y(n_929)
);

AOI21xp33_ASAP7_75t_L g930 ( 
.A1(n_658),
.A2(n_616),
.B(n_721),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_706),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_712),
.B(n_730),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_730),
.B(n_740),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_721),
.B(n_652),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_721),
.A2(n_603),
.B1(n_607),
.B2(n_652),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_606),
.A2(n_535),
.B(n_632),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_603),
.B(n_652),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_699),
.A2(n_617),
.B(n_632),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_603),
.B(n_652),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_606),
.A2(n_535),
.B(n_632),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_603),
.B(n_652),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_622),
.B(n_605),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_652),
.B(n_603),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_652),
.B(n_603),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_764),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_652),
.B(n_603),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_605),
.B(n_652),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_603),
.B(n_652),
.Y(n_948)
);

CKINVDCx6p67_ASAP7_75t_R g949 ( 
.A(n_749),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_652),
.B(n_603),
.Y(n_950)
);

NOR2xp67_ASAP7_75t_L g951 ( 
.A(n_641),
.B(n_410),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_605),
.B(n_652),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_603),
.B(n_652),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_622),
.B(n_605),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_699),
.A2(n_617),
.B(n_632),
.Y(n_955)
);

NAND2x1p5_ASAP7_75t_L g956 ( 
.A(n_646),
.B(n_533),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_652),
.B(n_603),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_605),
.A2(n_458),
.B(n_574),
.C(n_523),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_603),
.A2(n_652),
.B1(n_647),
.B2(n_635),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_947),
.B(n_952),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_912),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_831),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_947),
.B(n_952),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_882),
.A2(n_809),
.B1(n_785),
.B2(n_885),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_780),
.Y(n_965)
);

BUFx4f_ASAP7_75t_SL g966 ( 
.A(n_826),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_777),
.B(n_943),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_895),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_793),
.A2(n_957),
.B1(n_950),
.B2(n_946),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_944),
.B(n_942),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_954),
.B(n_797),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_SL g972 ( 
.A1(n_793),
.A2(n_877),
.B(n_888),
.C(n_786),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_885),
.B(n_886),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_959),
.A2(n_785),
.B1(n_774),
.B2(n_873),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_780),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_936),
.A2(n_940),
.B(n_939),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_799),
.Y(n_977)
);

AO21x2_ASAP7_75t_L g978 ( 
.A1(n_938),
.A2(n_955),
.B(n_847),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_928),
.A2(n_941),
.B(n_937),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_SL g980 ( 
.A1(n_913),
.A2(n_787),
.B(n_796),
.C(n_958),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_783),
.B(n_827),
.Y(n_981)
);

AO32x1_ASAP7_75t_L g982 ( 
.A1(n_935),
.A2(n_857),
.A3(n_814),
.B1(n_828),
.B2(n_781),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_788),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_941),
.B(n_948),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_949),
.Y(n_985)
);

CKINVDCx11_ASAP7_75t_R g986 ( 
.A(n_892),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_915),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_795),
.B(n_820),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_867),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_784),
.Y(n_990)
);

NOR2xp67_ASAP7_75t_L g991 ( 
.A(n_849),
.B(n_890),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_797),
.B(n_822),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_904),
.B(n_795),
.Y(n_993)
);

BUFx8_ASAP7_75t_L g994 ( 
.A(n_819),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_820),
.B(n_815),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_825),
.B(n_874),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_948),
.B(n_953),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_953),
.B(n_934),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_797),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_778),
.B(n_800),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_776),
.A2(n_798),
.B1(n_794),
.B2(n_792),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_SL g1002 ( 
.A(n_849),
.B(n_890),
.Y(n_1002)
);

INVx6_ASAP7_75t_L g1003 ( 
.A(n_867),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_801),
.B(n_896),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_867),
.B(n_823),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_916),
.A2(n_899),
.B(n_913),
.C(n_911),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_905),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_776),
.A2(n_914),
.B1(n_925),
.B2(n_797),
.Y(n_1008)
);

AO21x1_ASAP7_75t_L g1009 ( 
.A1(n_891),
.A2(n_813),
.B(n_877),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_791),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_799),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_945),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_838),
.Y(n_1013)
);

AOI21xp33_ASAP7_75t_L g1014 ( 
.A1(n_914),
.A2(n_908),
.B(n_929),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_837),
.B(n_808),
.Y(n_1015)
);

INVxp67_ASAP7_75t_SL g1016 ( 
.A(n_956),
.Y(n_1016)
);

O2A1O1Ixp5_ASAP7_75t_L g1017 ( 
.A1(n_891),
.A2(n_813),
.B(n_818),
.C(n_816),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_860),
.A2(n_810),
.B1(n_823),
.B2(n_951),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_898),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_805),
.B(n_806),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_810),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_842),
.B(n_856),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_901),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_867),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_822),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_775),
.A2(n_790),
.B(n_804),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_787),
.B(n_889),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_822),
.B(n_854),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_903),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_862),
.A2(n_865),
.B(n_871),
.C(n_868),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_909),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_862),
.A2(n_865),
.B(n_871),
.C(n_868),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_822),
.B(n_907),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_842),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_824),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_856),
.B(n_854),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_876),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_R g1038 ( 
.A(n_866),
.B(n_893),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_824),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_894),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_956),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_894),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_902),
.B(n_863),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_SL g1044 ( 
.A1(n_933),
.A2(n_859),
.B1(n_881),
.B2(n_870),
.Y(n_1044)
);

NOR3xp33_ASAP7_75t_L g1045 ( 
.A(n_917),
.B(n_869),
.C(n_930),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_883),
.Y(n_1046)
);

OAI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_789),
.A2(n_872),
.B1(n_864),
.B2(n_880),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_866),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_779),
.A2(n_782),
.B(n_846),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_824),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_902),
.B(n_876),
.Y(n_1051)
);

INVxp67_ASAP7_75t_L g1052 ( 
.A(n_875),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_876),
.B(n_878),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_876),
.A2(n_878),
.B1(n_786),
.B2(n_931),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_878),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_900),
.A2(n_844),
.B(n_832),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_928),
.A2(n_897),
.B(n_884),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_840),
.A2(n_841),
.B(n_833),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_817),
.B(n_887),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_910),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_920),
.B(n_922),
.Y(n_1061)
);

INVx3_ASAP7_75t_SL g1062 ( 
.A(n_926),
.Y(n_1062)
);

AND2x6_ASAP7_75t_L g1063 ( 
.A(n_923),
.B(n_924),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_812),
.A2(n_821),
.B(n_932),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_921),
.A2(n_918),
.B(n_906),
.C(n_843),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_848),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_802),
.A2(n_836),
.B(n_919),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_835),
.B(n_839),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_845),
.B(n_852),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_926),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_829),
.B(n_830),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_SL g1072 ( 
.A(n_879),
.B(n_858),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_811),
.A2(n_927),
.B1(n_851),
.B2(n_807),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_850),
.B(n_861),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_803),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_853),
.B(n_855),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_834),
.B(n_850),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_834),
.B(n_947),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_947),
.B(n_952),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_912),
.Y(n_1080)
);

O2A1O1Ixp33_ASAP7_75t_SL g1081 ( 
.A1(n_793),
.A2(n_809),
.B(n_882),
.C(n_877),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_942),
.B(n_954),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_947),
.B(n_952),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_780),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_831),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_947),
.B(n_952),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_SL g1087 ( 
.A(n_882),
.B(n_809),
.C(n_947),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_949),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_L g1089 ( 
.A(n_882),
.B(n_605),
.C(n_947),
.Y(n_1089)
);

NOR2x1p5_ASAP7_75t_L g1090 ( 
.A(n_882),
.B(n_581),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_947),
.B(n_952),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_912),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_947),
.B(n_952),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_947),
.B(n_952),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_947),
.A2(n_952),
.B1(n_882),
.B2(n_809),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_867),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_943),
.A2(n_535),
.B(n_944),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_942),
.B(n_954),
.Y(n_1098)
);

CKINVDCx16_ASAP7_75t_R g1099 ( 
.A(n_788),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_947),
.B(n_952),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_942),
.B(n_954),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_947),
.B(n_952),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_799),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_L g1104 ( 
.A1(n_813),
.A2(n_699),
.B(n_818),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1086),
.B(n_1094),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_962),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1049),
.A2(n_1026),
.B(n_1056),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_960),
.B(n_963),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1067),
.A2(n_1097),
.B(n_1065),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_960),
.B(n_963),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1089),
.A2(n_1006),
.B(n_1102),
.C(n_1100),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1100),
.A2(n_1102),
.B(n_1095),
.C(n_1014),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1079),
.A2(n_1091),
.B1(n_1093),
.B2(n_1083),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1085),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1057),
.A2(n_974),
.B(n_976),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_967),
.A2(n_964),
.B1(n_970),
.B2(n_1089),
.Y(n_1116)
);

OA21x2_ASAP7_75t_L g1117 ( 
.A1(n_1017),
.A2(n_979),
.B(n_1059),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1061),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_965),
.Y(n_1119)
);

NAND2xp33_ASAP7_75t_SL g1120 ( 
.A(n_1038),
.B(n_1048),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_969),
.B(n_1082),
.Y(n_1121)
);

AO22x1_ASAP7_75t_L g1122 ( 
.A1(n_973),
.A2(n_1045),
.B1(n_994),
.B2(n_993),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1007),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_1025),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1017),
.A2(n_997),
.B(n_1043),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_989),
.Y(n_1126)
);

INVx3_ASAP7_75t_SL g1127 ( 
.A(n_985),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_989),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_975),
.Y(n_1129)
);

AOI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1072),
.A2(n_1077),
.B(n_1104),
.Y(n_1130)
);

INVx8_ASAP7_75t_L g1131 ( 
.A(n_1025),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1087),
.A2(n_973),
.B(n_1081),
.C(n_980),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1028),
.B(n_1005),
.Y(n_1133)
);

AOI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1073),
.A2(n_1078),
.B(n_1064),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1098),
.B(n_1101),
.Y(n_1135)
);

AO32x2_ASAP7_75t_L g1136 ( 
.A1(n_1008),
.A2(n_1001),
.A3(n_1044),
.B1(n_1032),
.B2(n_1030),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1088),
.Y(n_1137)
);

AOI221x1_ASAP7_75t_L g1138 ( 
.A1(n_1045),
.A2(n_1087),
.B1(n_1027),
.B2(n_1058),
.C(n_1074),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1051),
.A2(n_995),
.B1(n_1036),
.B2(n_1027),
.Y(n_1139)
);

NAND3x1_ASAP7_75t_L g1140 ( 
.A(n_981),
.B(n_988),
.C(n_1033),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_998),
.B(n_997),
.Y(n_1141)
);

AOI21xp33_ASAP7_75t_L g1142 ( 
.A1(n_1047),
.A2(n_978),
.B(n_998),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1004),
.Y(n_1143)
);

AOI21x1_ASAP7_75t_L g1144 ( 
.A1(n_984),
.A2(n_1018),
.B(n_1069),
.Y(n_1144)
);

AO32x2_ASAP7_75t_L g1145 ( 
.A1(n_982),
.A2(n_972),
.A3(n_1009),
.B1(n_978),
.B2(n_1070),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1012),
.Y(n_1146)
);

AO21x1_ASAP7_75t_L g1147 ( 
.A1(n_1047),
.A2(n_1068),
.B(n_1054),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1071),
.A2(n_1076),
.B(n_1068),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1013),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_989),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_968),
.Y(n_1151)
);

NOR2xp67_ASAP7_75t_SL g1152 ( 
.A(n_1099),
.B(n_983),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_994),
.Y(n_1153)
);

AOI21xp33_ASAP7_75t_L g1154 ( 
.A1(n_996),
.A2(n_995),
.B(n_1052),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1076),
.A2(n_1016),
.B(n_982),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_987),
.Y(n_1156)
);

OA21x2_ASAP7_75t_L g1157 ( 
.A1(n_1075),
.A2(n_1015),
.B(n_1052),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1016),
.A2(n_982),
.B(n_1053),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1033),
.B(n_1084),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1041),
.A2(n_1022),
.B(n_971),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1003),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_977),
.A2(n_1103),
.B(n_1021),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1019),
.A2(n_1029),
.B(n_1023),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1031),
.A2(n_1066),
.B(n_1060),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1000),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_SL g1166 ( 
.A1(n_1037),
.A2(n_1055),
.B(n_1070),
.Y(n_1166)
);

BUFx4f_ASAP7_75t_SL g1167 ( 
.A(n_1040),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_977),
.A2(n_1103),
.B(n_1011),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1028),
.A2(n_1066),
.B1(n_1010),
.B2(n_990),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_992),
.A2(n_1002),
.B(n_1000),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_999),
.A2(n_1005),
.B(n_1020),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_961),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1034),
.A2(n_1003),
.B1(n_1024),
.B2(n_1096),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_999),
.A2(n_1021),
.B(n_1011),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_991),
.A2(n_1025),
.B(n_1050),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1080),
.B(n_1092),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1090),
.A2(n_1063),
.B(n_1062),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1025),
.A2(n_1039),
.B(n_1050),
.Y(n_1178)
);

NOR2x1_ASAP7_75t_R g1179 ( 
.A(n_986),
.B(n_1046),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1024),
.B(n_1096),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1063),
.A2(n_1039),
.B(n_1050),
.Y(n_1181)
);

OA21x2_ASAP7_75t_L g1182 ( 
.A1(n_1042),
.A2(n_1063),
.B(n_1039),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1063),
.A2(n_1003),
.B(n_1035),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1024),
.A2(n_1096),
.B(n_966),
.C(n_1035),
.Y(n_1184)
);

AND2x6_ASAP7_75t_L g1185 ( 
.A(n_1024),
.B(n_1096),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1035),
.A2(n_1009),
.A3(n_1065),
.B(n_1073),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_966),
.A2(n_947),
.B(n_952),
.C(n_1086),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1086),
.A2(n_947),
.B(n_952),
.C(n_1094),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1049),
.A2(n_782),
.B(n_1026),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_983),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1067),
.A2(n_1097),
.B(n_944),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1067),
.A2(n_1097),
.B(n_944),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_965),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1049),
.A2(n_782),
.B(n_1026),
.Y(n_1194)
);

O2A1O1Ixp5_ASAP7_75t_L g1195 ( 
.A1(n_1086),
.A2(n_809),
.B(n_882),
.C(n_947),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1097),
.A2(n_1014),
.B(n_1017),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_962),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1086),
.A2(n_1094),
.B1(n_947),
.B2(n_952),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_985),
.Y(n_1199)
);

AO21x2_ASAP7_75t_L g1200 ( 
.A1(n_1057),
.A2(n_976),
.B(n_1067),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1009),
.A2(n_1065),
.A3(n_1073),
.B(n_976),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1067),
.A2(n_1097),
.B(n_944),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1035),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_983),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1097),
.A2(n_1014),
.B(n_1017),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1097),
.A2(n_1014),
.B(n_1017),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1086),
.B(n_1094),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1067),
.A2(n_1097),
.B(n_944),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_962),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1067),
.A2(n_1097),
.B(n_944),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1067),
.A2(n_1097),
.B(n_944),
.Y(n_1211)
);

AOI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1072),
.A2(n_1077),
.B(n_1104),
.Y(n_1212)
);

OA21x2_ASAP7_75t_L g1213 ( 
.A1(n_1057),
.A2(n_1017),
.B(n_979),
.Y(n_1213)
);

NOR2xp67_ASAP7_75t_L g1214 ( 
.A(n_1052),
.B(n_715),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_962),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_SL g1216 ( 
.A1(n_1006),
.A2(n_793),
.B(n_882),
.C(n_809),
.Y(n_1216)
);

AO31x2_ASAP7_75t_L g1217 ( 
.A1(n_1009),
.A2(n_1065),
.A3(n_1073),
.B(n_976),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1097),
.A2(n_1014),
.B(n_1017),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1067),
.A2(n_1097),
.B(n_944),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_973),
.B(n_947),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1067),
.A2(n_1097),
.B(n_944),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_983),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1086),
.B(n_1094),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1097),
.A2(n_1014),
.B(n_1017),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_SL g1225 ( 
.A(n_1086),
.B(n_793),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1067),
.A2(n_1097),
.B(n_944),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1049),
.A2(n_782),
.B(n_1026),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1049),
.A2(n_782),
.B(n_1026),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_973),
.B(n_947),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1067),
.A2(n_1097),
.B(n_944),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_SL g1231 ( 
.A1(n_974),
.A2(n_793),
.B(n_1006),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1067),
.A2(n_1097),
.B(n_944),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1097),
.A2(n_1014),
.B(n_1017),
.Y(n_1233)
);

AO21x2_ASAP7_75t_L g1234 ( 
.A1(n_1057),
.A2(n_976),
.B(n_1067),
.Y(n_1234)
);

CKINVDCx16_ASAP7_75t_R g1235 ( 
.A(n_1099),
.Y(n_1235)
);

O2A1O1Ixp5_ASAP7_75t_SL g1236 ( 
.A1(n_1014),
.A2(n_1077),
.B(n_882),
.C(n_813),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1049),
.A2(n_782),
.B(n_1026),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1097),
.A2(n_1014),
.B(n_1017),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1028),
.B(n_1005),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_989),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1067),
.A2(n_1097),
.B(n_944),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_965),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1180),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1190),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1220),
.B(n_1229),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1225),
.A2(n_1198),
.B1(n_1116),
.B2(n_1147),
.Y(n_1246)
);

INVx4_ASAP7_75t_L g1247 ( 
.A(n_1131),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1204),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_1235),
.Y(n_1249)
);

BUFx12f_ASAP7_75t_L g1250 ( 
.A(n_1137),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1225),
.A2(n_1105),
.B1(n_1207),
.B2(n_1223),
.Y(n_1251)
);

INVx6_ASAP7_75t_L g1252 ( 
.A(n_1131),
.Y(n_1252)
);

INVx6_ASAP7_75t_L g1253 ( 
.A(n_1131),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1106),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1105),
.A2(n_1207),
.B1(n_1223),
.B2(n_1108),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1222),
.Y(n_1256)
);

BUFx8_ASAP7_75t_L g1257 ( 
.A(n_1193),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1108),
.A2(n_1110),
.B1(n_1116),
.B2(n_1113),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1135),
.B(n_1159),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_SL g1260 ( 
.A1(n_1110),
.A2(n_1113),
.B1(n_1136),
.B2(n_1141),
.Y(n_1260)
);

CKINVDCx6p67_ASAP7_75t_R g1261 ( 
.A(n_1127),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1141),
.A2(n_1121),
.B1(n_1165),
.B2(n_1135),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_SL g1263 ( 
.A1(n_1136),
.A2(n_1139),
.B1(n_1238),
.B2(n_1206),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_SL g1264 ( 
.A1(n_1136),
.A2(n_1139),
.B1(n_1238),
.B2(n_1206),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1142),
.A2(n_1121),
.B1(n_1154),
.B2(n_1125),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1167),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1142),
.A2(n_1154),
.B1(n_1125),
.B2(n_1233),
.Y(n_1267)
);

CKINVDCx6p67_ASAP7_75t_R g1268 ( 
.A(n_1153),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1196),
.A2(n_1233),
.B1(n_1224),
.B2(n_1205),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1242),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1214),
.A2(n_1148),
.B1(n_1115),
.B2(n_1205),
.Y(n_1271)
);

OAI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1143),
.A2(n_1164),
.B1(n_1169),
.B2(n_1129),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1114),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1218),
.A2(n_1213),
.B1(n_1163),
.B2(n_1164),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1197),
.Y(n_1275)
);

INVx6_ASAP7_75t_L g1276 ( 
.A(n_1124),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1151),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1187),
.A2(n_1188),
.B1(n_1122),
.B2(n_1140),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1199),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1133),
.B(n_1239),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1152),
.A2(n_1112),
.B1(n_1239),
.B2(n_1133),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1180),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1119),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1200),
.A2(n_1234),
.B1(n_1169),
.B2(n_1129),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1111),
.B(n_1118),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1109),
.A2(n_1234),
.B1(n_1200),
.B2(n_1149),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1209),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1215),
.Y(n_1288)
);

BUFx4f_ASAP7_75t_L g1289 ( 
.A(n_1185),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1119),
.Y(n_1290)
);

OAI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1138),
.A2(n_1123),
.B1(n_1146),
.B2(n_1156),
.Y(n_1291)
);

CKINVDCx14_ASAP7_75t_R g1292 ( 
.A(n_1120),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1176),
.Y(n_1293)
);

CKINVDCx6p67_ASAP7_75t_R g1294 ( 
.A(n_1161),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1172),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1157),
.Y(n_1296)
);

BUFx4f_ASAP7_75t_SL g1297 ( 
.A(n_1126),
.Y(n_1297)
);

CKINVDCx11_ASAP7_75t_R g1298 ( 
.A(n_1179),
.Y(n_1298)
);

NAND2x1p5_ASAP7_75t_L g1299 ( 
.A(n_1181),
.B(n_1177),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1128),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1231),
.A2(n_1170),
.B1(n_1132),
.B2(n_1171),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1155),
.A2(n_1216),
.B1(n_1117),
.B2(n_1221),
.Y(n_1302)
);

BUFx5_ASAP7_75t_L g1303 ( 
.A(n_1185),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1191),
.A2(n_1241),
.B1(n_1192),
.B2(n_1232),
.Y(n_1304)
);

CKINVDCx11_ASAP7_75t_R g1305 ( 
.A(n_1128),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1203),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1128),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1117),
.A2(n_1219),
.B1(n_1202),
.B2(n_1226),
.Y(n_1308)
);

BUFx4_ASAP7_75t_SL g1309 ( 
.A(n_1184),
.Y(n_1309)
);

OAI21xp33_ASAP7_75t_L g1310 ( 
.A1(n_1236),
.A2(n_1211),
.B(n_1230),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1203),
.Y(n_1311)
);

CKINVDCx11_ASAP7_75t_R g1312 ( 
.A(n_1150),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1208),
.A2(n_1210),
.B1(n_1158),
.B2(n_1160),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1195),
.A2(n_1182),
.B1(n_1185),
.B2(n_1173),
.Y(n_1314)
);

OAI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1182),
.A2(n_1144),
.B1(n_1173),
.B2(n_1124),
.Y(n_1315)
);

INVx5_ASAP7_75t_L g1316 ( 
.A(n_1150),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1174),
.A2(n_1166),
.B1(n_1183),
.B2(n_1240),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1183),
.A2(n_1168),
.B1(n_1162),
.B2(n_1107),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1186),
.B(n_1178),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1175),
.A2(n_1134),
.B1(n_1130),
.B2(n_1212),
.Y(n_1320)
);

BUFx12f_ASAP7_75t_L g1321 ( 
.A(n_1186),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1189),
.A2(n_1194),
.B1(n_1227),
.B2(n_1228),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1145),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1237),
.A2(n_1145),
.B1(n_1201),
.B2(n_1217),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1201),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1217),
.A2(n_1225),
.B1(n_1094),
.B2(n_1086),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1217),
.Y(n_1327)
);

INVx5_ASAP7_75t_L g1328 ( 
.A(n_1185),
.Y(n_1328)
);

BUFx8_ASAP7_75t_L g1329 ( 
.A(n_1193),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1220),
.B(n_1086),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1198),
.A2(n_1094),
.B1(n_1086),
.B2(n_963),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_SL g1332 ( 
.A1(n_1225),
.A2(n_1094),
.B1(n_1086),
.B2(n_952),
.Y(n_1332)
);

BUFx4f_ASAP7_75t_SL g1333 ( 
.A(n_1190),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1220),
.A2(n_1094),
.B1(n_1086),
.B2(n_1089),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1198),
.A2(n_1094),
.B1(n_1086),
.B2(n_963),
.Y(n_1335)
);

INVx6_ASAP7_75t_L g1336 ( 
.A(n_1131),
.Y(n_1336)
);

OAI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1198),
.A2(n_1095),
.B1(n_1083),
.B2(n_1091),
.Y(n_1337)
);

INVx8_ASAP7_75t_L g1338 ( 
.A(n_1131),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1220),
.A2(n_1094),
.B1(n_1086),
.B2(n_1089),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1193),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1225),
.A2(n_1094),
.B1(n_1086),
.B2(n_952),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1235),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1119),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1198),
.A2(n_1094),
.B1(n_1086),
.B2(n_963),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1135),
.B(n_1082),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1220),
.A2(n_1094),
.B1(n_1086),
.B2(n_1089),
.Y(n_1346)
);

BUFx10_ASAP7_75t_L g1347 ( 
.A(n_1137),
.Y(n_1347)
);

INVxp67_ASAP7_75t_SL g1348 ( 
.A(n_1148),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1258),
.B(n_1260),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1296),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1276),
.Y(n_1351)
);

OA21x2_ASAP7_75t_L g1352 ( 
.A1(n_1310),
.A2(n_1304),
.B(n_1324),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1290),
.Y(n_1353)
);

BUFx4f_ASAP7_75t_SL g1354 ( 
.A(n_1250),
.Y(n_1354)
);

CKINVDCx14_ASAP7_75t_R g1355 ( 
.A(n_1298),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1299),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1325),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1323),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1326),
.B(n_1263),
.Y(n_1359)
);

NOR2x1_ASAP7_75t_SL g1360 ( 
.A(n_1301),
.B(n_1328),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1331),
.A2(n_1335),
.B1(n_1344),
.B2(n_1278),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1319),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1321),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1327),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1254),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1326),
.B(n_1263),
.Y(n_1366)
);

AO21x2_ASAP7_75t_L g1367 ( 
.A1(n_1322),
.A2(n_1315),
.B(n_1320),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1273),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1348),
.Y(n_1369)
);

AOI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1285),
.A2(n_1275),
.B(n_1288),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1315),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1287),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1276),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1291),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1267),
.B(n_1269),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1330),
.B(n_1245),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1293),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1262),
.A2(n_1291),
.B(n_1337),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1264),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1313),
.A2(n_1304),
.B(n_1318),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1264),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1318),
.B(n_1271),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1267),
.B(n_1269),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1286),
.A2(n_1274),
.B(n_1317),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1286),
.Y(n_1385)
);

INVx2_ASAP7_75t_SL g1386 ( 
.A(n_1316),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1260),
.B(n_1265),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1316),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1274),
.A2(n_1317),
.B(n_1284),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1258),
.B(n_1255),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1265),
.A2(n_1246),
.B(n_1311),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1343),
.Y(n_1392)
);

BUFx2_ASAP7_75t_R g1393 ( 
.A(n_1283),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1332),
.B(n_1341),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1306),
.A2(n_1281),
.B(n_1295),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1262),
.Y(n_1396)
);

INVx4_ASAP7_75t_L g1397 ( 
.A(n_1328),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1340),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1272),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1277),
.A2(n_1308),
.B(n_1282),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1345),
.B(n_1259),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1255),
.B(n_1337),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1303),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1251),
.B(n_1346),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1303),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1302),
.Y(n_1406)
);

INVx2_ASAP7_75t_SL g1407 ( 
.A(n_1316),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1302),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1289),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1270),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1314),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1251),
.B(n_1332),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1314),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1308),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1341),
.B(n_1243),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1334),
.B(n_1346),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1334),
.B(n_1339),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1280),
.B(n_1247),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1289),
.A2(n_1339),
.B(n_1280),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1309),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1361),
.A2(n_1292),
.B(n_1342),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1376),
.B(n_1266),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1401),
.B(n_1402),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1394),
.A2(n_1416),
.B1(n_1412),
.B2(n_1417),
.Y(n_1424)
);

AOI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1417),
.A2(n_1359),
.B1(n_1366),
.B2(n_1387),
.C(n_1374),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1412),
.A2(n_1249),
.B1(n_1307),
.B2(n_1261),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1384),
.A2(n_1309),
.B(n_1297),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1364),
.B(n_1300),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1364),
.B(n_1312),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1359),
.B(n_1305),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_SL g1431 ( 
.A(n_1393),
.B(n_1333),
.Y(n_1431)
);

OR2x6_ASAP7_75t_L g1432 ( 
.A(n_1369),
.B(n_1338),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1350),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1366),
.B(n_1294),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1411),
.B(n_1279),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1419),
.B(n_1347),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1413),
.B(n_1347),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1402),
.B(n_1329),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1410),
.B(n_1244),
.Y(n_1439)
);

A2O1A1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1416),
.A2(n_1338),
.B(n_1248),
.C(n_1256),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1375),
.A2(n_1383),
.B(n_1349),
.C(n_1404),
.Y(n_1441)
);

AO22x2_ASAP7_75t_L g1442 ( 
.A1(n_1375),
.A2(n_1257),
.B1(n_1329),
.B2(n_1297),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1362),
.B(n_1268),
.Y(n_1443)
);

NOR2x1_ASAP7_75t_SL g1444 ( 
.A(n_1370),
.B(n_1333),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1413),
.B(n_1357),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1350),
.Y(n_1446)
);

AOI221xp5_ASAP7_75t_L g1447 ( 
.A1(n_1387),
.A2(n_1257),
.B1(n_1253),
.B2(n_1252),
.C(n_1336),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1392),
.B(n_1253),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1356),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1365),
.Y(n_1450)
);

AO21x1_ASAP7_75t_L g1451 ( 
.A1(n_1349),
.A2(n_1336),
.B(n_1383),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1420),
.A2(n_1336),
.B1(n_1404),
.B2(n_1390),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1403),
.B(n_1405),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1379),
.B(n_1381),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1379),
.B(n_1381),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1415),
.B(n_1362),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1356),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1380),
.A2(n_1400),
.B(n_1384),
.Y(n_1458)
);

AO21x1_ASAP7_75t_L g1459 ( 
.A1(n_1374),
.A2(n_1390),
.B(n_1399),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1368),
.B(n_1385),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1385),
.B(n_1371),
.Y(n_1461)
);

AO32x2_ASAP7_75t_L g1462 ( 
.A1(n_1397),
.A2(n_1386),
.A3(n_1388),
.B1(n_1407),
.B2(n_1358),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1403),
.B(n_1405),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1371),
.B(n_1414),
.Y(n_1464)
);

INVxp67_ASAP7_75t_L g1465 ( 
.A(n_1353),
.Y(n_1465)
);

A2O1A1Ixp33_ASAP7_75t_L g1466 ( 
.A1(n_1419),
.A2(n_1389),
.B(n_1396),
.C(n_1382),
.Y(n_1466)
);

O2A1O1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1420),
.A2(n_1378),
.B(n_1396),
.C(n_1398),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1393),
.B(n_1398),
.Y(n_1468)
);

A2O1A1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1389),
.A2(n_1382),
.B(n_1408),
.C(n_1406),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1414),
.B(n_1372),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1450),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_L g1472 ( 
.A(n_1422),
.B(n_1438),
.Y(n_1472)
);

NOR2xp67_ASAP7_75t_L g1473 ( 
.A(n_1449),
.B(n_1457),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1433),
.Y(n_1474)
);

NOR2x1p5_ASAP7_75t_L g1475 ( 
.A(n_1443),
.B(n_1409),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1456),
.B(n_1461),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1433),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1436),
.A2(n_1378),
.B1(n_1382),
.B2(n_1363),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1453),
.B(n_1463),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1470),
.B(n_1378),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1453),
.B(n_1367),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1470),
.B(n_1378),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1463),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1446),
.Y(n_1484)
);

OR2x6_ASAP7_75t_SL g1485 ( 
.A(n_1464),
.B(n_1363),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1464),
.B(n_1367),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1446),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1425),
.A2(n_1382),
.B1(n_1363),
.B2(n_1408),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1460),
.B(n_1406),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1463),
.B(n_1352),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1437),
.A2(n_1409),
.B1(n_1418),
.B2(n_1391),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1437),
.A2(n_1409),
.B1(n_1418),
.B2(n_1391),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1458),
.B(n_1352),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1462),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1459),
.B(n_1377),
.Y(n_1495)
);

AOI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1424),
.A2(n_1409),
.B1(n_1418),
.B2(n_1395),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1474),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1474),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1477),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1494),
.B(n_1469),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1490),
.B(n_1462),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1473),
.B(n_1481),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1471),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1471),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1472),
.B(n_1451),
.Y(n_1505)
);

AND2x4_ASAP7_75t_SL g1506 ( 
.A(n_1496),
.B(n_1432),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1485),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1488),
.A2(n_1451),
.B1(n_1452),
.B2(n_1459),
.Y(n_1508)
);

OAI322xp33_ASAP7_75t_L g1509 ( 
.A1(n_1486),
.A2(n_1467),
.A3(n_1423),
.B1(n_1465),
.B2(n_1426),
.C1(n_1454),
.C2(n_1455),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1489),
.B(n_1439),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1484),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1493),
.A2(n_1495),
.B(n_1482),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1476),
.B(n_1445),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1484),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1487),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1487),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1478),
.A2(n_1442),
.B1(n_1441),
.B2(n_1435),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1485),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_1485),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1496),
.A2(n_1466),
.B1(n_1426),
.B2(n_1442),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1483),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1495),
.A2(n_1360),
.B(n_1444),
.Y(n_1522)
);

AOI221xp5_ASAP7_75t_L g1523 ( 
.A1(n_1480),
.A2(n_1421),
.B1(n_1442),
.B2(n_1455),
.C(n_1454),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1501),
.B(n_1479),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1511),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1511),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1503),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1497),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1501),
.B(n_1479),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1503),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1512),
.B(n_1476),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1520),
.A2(n_1442),
.B1(n_1434),
.B2(n_1447),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1501),
.B(n_1479),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1503),
.Y(n_1534)
);

NAND2xp33_ASAP7_75t_SL g1535 ( 
.A(n_1505),
.B(n_1475),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1504),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1502),
.B(n_1521),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1502),
.B(n_1473),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1504),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1514),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1512),
.B(n_1480),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1512),
.B(n_1476),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1507),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1514),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1497),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1498),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1502),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1515),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1498),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1499),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1516),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1500),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1543),
.B(n_1507),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1527),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1545),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1545),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1535),
.B(n_1355),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1535),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1527),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1532),
.A2(n_1520),
.B1(n_1517),
.B2(n_1508),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1527),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1546),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1546),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1527),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1530),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1530),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1530),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1530),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1552),
.B(n_1500),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1525),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1532),
.A2(n_1517),
.B1(n_1523),
.B2(n_1434),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1534),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1525),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1534),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1526),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1526),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_SL g1577 ( 
.A(n_1543),
.B(n_1509),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1552),
.B(n_1500),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1541),
.B(n_1512),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1540),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1543),
.B(n_1507),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1540),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1544),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1541),
.B(n_1512),
.Y(n_1584)
);

NOR4xp25_ASAP7_75t_L g1585 ( 
.A(n_1531),
.B(n_1509),
.C(n_1523),
.D(n_1519),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1524),
.B(n_1510),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1544),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1534),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_SL g1589 ( 
.A(n_1538),
.B(n_1431),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1534),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1548),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1536),
.Y(n_1592)
);

NOR2xp67_ASAP7_75t_L g1593 ( 
.A(n_1547),
.B(n_1538),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1524),
.B(n_1513),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1569),
.Y(n_1595)
);

INVxp33_ASAP7_75t_L g1596 ( 
.A(n_1557),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1558),
.B(n_1589),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1553),
.B(n_1581),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1570),
.Y(n_1599)
);

AND2x4_ASAP7_75t_SL g1600 ( 
.A(n_1553),
.B(n_1547),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1569),
.B(n_1531),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1570),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1581),
.B(n_1593),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1577),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1573),
.Y(n_1605)
);

NOR3xp33_ASAP7_75t_L g1606 ( 
.A(n_1560),
.B(n_1468),
.C(n_1448),
.Y(n_1606)
);

AOI22x1_ASAP7_75t_L g1607 ( 
.A1(n_1585),
.A2(n_1519),
.B1(n_1518),
.B2(n_1430),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1560),
.B(n_1518),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1566),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1555),
.Y(n_1610)
);

NAND2x1p5_ASAP7_75t_L g1611 ( 
.A(n_1571),
.B(n_1427),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1593),
.B(n_1538),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1571),
.A2(n_1430),
.B1(n_1427),
.B2(n_1435),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1578),
.B(n_1538),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1573),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1578),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1586),
.B(n_1524),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1594),
.B(n_1531),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1555),
.B(n_1538),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1575),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1556),
.B(n_1538),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1556),
.B(n_1547),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1562),
.B(n_1529),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1562),
.B(n_1547),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1563),
.B(n_1542),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1563),
.B(n_1547),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1579),
.B(n_1542),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1579),
.B(n_1542),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1575),
.B(n_1529),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1598),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1599),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1598),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1606),
.B(n_1529),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1603),
.Y(n_1634)
);

OAI32xp33_ASAP7_75t_L g1635 ( 
.A1(n_1611),
.A2(n_1584),
.A3(n_1591),
.B1(n_1576),
.B2(n_1580),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1600),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1599),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1604),
.B(n_1533),
.Y(n_1638)
);

AOI211xp5_ASAP7_75t_L g1639 ( 
.A1(n_1608),
.A2(n_1584),
.B(n_1522),
.C(n_1440),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1602),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1597),
.A2(n_1506),
.B1(n_1475),
.B2(n_1537),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1602),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1607),
.A2(n_1522),
.B(n_1576),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1605),
.Y(n_1644)
);

NAND2x1_ASAP7_75t_L g1645 ( 
.A(n_1603),
.B(n_1537),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1605),
.Y(n_1646)
);

NOR3xp33_ASAP7_75t_SL g1647 ( 
.A(n_1607),
.B(n_1354),
.C(n_1580),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1616),
.B(n_1533),
.Y(n_1648)
);

AOI321xp33_ASAP7_75t_L g1649 ( 
.A1(n_1613),
.A2(n_1491),
.A3(n_1492),
.B1(n_1493),
.B2(n_1429),
.C(n_1587),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1600),
.Y(n_1650)
);

AOI31xp33_ASAP7_75t_L g1651 ( 
.A1(n_1596),
.A2(n_1429),
.A3(n_1443),
.B(n_1428),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1613),
.A2(n_1583),
.B(n_1582),
.Y(n_1652)
);

NOR2xp67_ASAP7_75t_SL g1653 ( 
.A(n_1595),
.B(n_1409),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1610),
.B(n_1614),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1654),
.Y(n_1655)
);

OAI21xp33_ASAP7_75t_L g1656 ( 
.A1(n_1647),
.A2(n_1611),
.B(n_1614),
.Y(n_1656)
);

AOI211xp5_ASAP7_75t_SL g1657 ( 
.A1(n_1643),
.A2(n_1652),
.B(n_1639),
.C(n_1651),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1654),
.Y(n_1658)
);

AOI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1635),
.A2(n_1611),
.B1(n_1610),
.B2(n_1621),
.C(n_1619),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1632),
.A2(n_1633),
.B1(n_1630),
.B2(n_1638),
.Y(n_1660)
);

OAI21xp5_ASAP7_75t_SL g1661 ( 
.A1(n_1641),
.A2(n_1621),
.B(n_1619),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1630),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1654),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1631),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1650),
.A2(n_1620),
.B1(n_1615),
.B2(n_1617),
.Y(n_1665)
);

OAI21xp33_ASAP7_75t_L g1666 ( 
.A1(n_1647),
.A2(n_1623),
.B(n_1629),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1634),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1634),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1648),
.B(n_1618),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1637),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1636),
.A2(n_1612),
.B1(n_1506),
.B2(n_1622),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1645),
.Y(n_1672)
);

OAI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1649),
.A2(n_1601),
.B1(n_1612),
.B2(n_1618),
.C(n_1615),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1663),
.B(n_1650),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1655),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1657),
.A2(n_1642),
.B(n_1640),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1668),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1655),
.Y(n_1678)
);

NAND2xp33_ASAP7_75t_L g1679 ( 
.A(n_1655),
.B(n_1644),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1658),
.Y(n_1680)
);

OAI31xp33_ASAP7_75t_L g1681 ( 
.A1(n_1656),
.A2(n_1646),
.A3(n_1601),
.B(n_1622),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1658),
.B(n_1624),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1660),
.B(n_1625),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1660),
.B(n_1624),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1678),
.B(n_1662),
.Y(n_1685)
);

NAND4xp25_ASAP7_75t_L g1686 ( 
.A(n_1674),
.B(n_1665),
.C(n_1659),
.D(n_1671),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1674),
.B(n_1667),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1683),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1677),
.B(n_1666),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_1675),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1680),
.Y(n_1691)
);

NOR3x1_ASAP7_75t_L g1692 ( 
.A(n_1684),
.B(n_1661),
.C(n_1664),
.Y(n_1692)
);

NAND3xp33_ASAP7_75t_L g1693 ( 
.A(n_1676),
.B(n_1665),
.C(n_1667),
.Y(n_1693)
);

OAI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1681),
.A2(n_1673),
.B1(n_1669),
.B2(n_1672),
.C(n_1670),
.Y(n_1694)
);

AOI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1693),
.A2(n_1679),
.B1(n_1682),
.B2(n_1672),
.C(n_1653),
.Y(n_1695)
);

AOI211xp5_ASAP7_75t_SL g1696 ( 
.A1(n_1688),
.A2(n_1679),
.B(n_1620),
.C(n_1626),
.Y(n_1696)
);

AOI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1694),
.A2(n_1653),
.B1(n_1626),
.B2(n_1625),
.C(n_1609),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1687),
.Y(n_1698)
);

AOI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1686),
.A2(n_1609),
.B1(n_1628),
.B2(n_1627),
.C(n_1567),
.Y(n_1699)
);

NOR4xp25_ASAP7_75t_L g1700 ( 
.A(n_1685),
.B(n_1628),
.C(n_1627),
.D(n_1567),
.Y(n_1700)
);

AOI222xp33_ASAP7_75t_L g1701 ( 
.A1(n_1689),
.A2(n_1587),
.B1(n_1582),
.B2(n_1591),
.C1(n_1583),
.C2(n_1567),
.Y(n_1701)
);

AOI32xp33_ASAP7_75t_L g1702 ( 
.A1(n_1696),
.A2(n_1695),
.A3(n_1698),
.B1(n_1690),
.B2(n_1697),
.Y(n_1702)
);

OAI211xp5_ASAP7_75t_L g1703 ( 
.A1(n_1700),
.A2(n_1691),
.B(n_1692),
.C(n_1574),
.Y(n_1703)
);

O2A1O1Ixp33_ASAP7_75t_L g1704 ( 
.A1(n_1699),
.A2(n_1701),
.B(n_1554),
.C(n_1592),
.Y(n_1704)
);

AOI222xp33_ASAP7_75t_L g1705 ( 
.A1(n_1697),
.A2(n_1566),
.B1(n_1568),
.B2(n_1590),
.C1(n_1572),
.C2(n_1574),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1697),
.A2(n_1537),
.B1(n_1592),
.B2(n_1554),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1698),
.B(n_1537),
.Y(n_1707)
);

NOR2x1_ASAP7_75t_L g1708 ( 
.A(n_1703),
.B(n_1566),
.Y(n_1708)
);

XNOR2x1_ASAP7_75t_L g1709 ( 
.A(n_1707),
.B(n_1428),
.Y(n_1709)
);

NAND4xp75_ASAP7_75t_L g1710 ( 
.A(n_1706),
.B(n_1590),
.C(n_1568),
.D(n_1572),
.Y(n_1710)
);

NOR2x1_ASAP7_75t_L g1711 ( 
.A(n_1704),
.B(n_1568),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1705),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1712),
.A2(n_1702),
.B(n_1574),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1709),
.B(n_1559),
.Y(n_1714)
);

NOR3xp33_ASAP7_75t_L g1715 ( 
.A(n_1708),
.B(n_1590),
.C(n_1572),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1714),
.A2(n_1710),
.B1(n_1711),
.B2(n_1564),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_SL g1717 ( 
.A1(n_1716),
.A2(n_1713),
.B1(n_1715),
.B2(n_1561),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1717),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1717),
.A2(n_1588),
.B1(n_1559),
.B2(n_1565),
.C(n_1561),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1718),
.A2(n_1588),
.B1(n_1565),
.B2(n_1564),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1719),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1537),
.B1(n_1536),
.B2(n_1539),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1720),
.B(n_1536),
.Y(n_1723)
);

INVxp33_ASAP7_75t_L g1724 ( 
.A(n_1723),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1724),
.A2(n_1722),
.B(n_1537),
.Y(n_1725)
);

INVxp67_ASAP7_75t_SL g1726 ( 
.A(n_1725),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1726),
.A2(n_1528),
.B1(n_1549),
.B2(n_1550),
.C(n_1551),
.Y(n_1727)
);

AOI211xp5_ASAP7_75t_L g1728 ( 
.A1(n_1727),
.A2(n_1409),
.B(n_1351),
.C(n_1373),
.Y(n_1728)
);


endmodule