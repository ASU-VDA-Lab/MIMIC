module fake_jpeg_7788_n_256 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_SL g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_1),
.B(n_2),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_3),
.Y(n_61)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_21),
.B1(n_31),
.B2(n_30),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_54),
.B1(n_59),
.B2(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_51),
.B(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_21),
.B1(n_31),
.B2(n_30),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_20),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_61),
.B(n_64),
.C(n_23),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_21),
.B1(n_31),
.B2(n_20),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_56),
.A2(n_69),
.B1(n_6),
.B2(n_8),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_20),
.B1(n_30),
.B2(n_26),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_34),
.B1(n_32),
.B2(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_3),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_19),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_35),
.A2(n_29),
.B1(n_23),
.B2(n_28),
.Y(n_69)
);

OAI32xp33_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_24),
.A3(n_28),
.B1(n_18),
.B2(n_29),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_49),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_24),
.B1(n_28),
.B2(n_18),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_23),
.B1(n_29),
.B2(n_18),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_100),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_87),
.Y(n_121)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

BUFx2_ASAP7_75t_SL g116 ( 
.A(n_84),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_25),
.B1(n_17),
.B2(n_7),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_98),
.B1(n_58),
.B2(n_46),
.Y(n_118)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_88),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_25),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_17),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_3),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_6),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_50),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_54),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_101),
.A2(n_102),
.B1(n_59),
.B2(n_64),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_50),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_108),
.B1(n_124),
.B2(n_95),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_100),
.A2(n_67),
.B1(n_64),
.B2(n_49),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g111 ( 
.A(n_87),
.B(n_64),
.CI(n_49),
.CON(n_111),
.SN(n_111)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_75),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_9),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_67),
.B(n_58),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_83),
.B(n_88),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_86),
.B1(n_82),
.B2(n_97),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_80),
.A2(n_49),
.B1(n_46),
.B2(n_65),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_65),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_85),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_118),
.A2(n_89),
.B1(n_74),
.B2(n_73),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_129),
.A2(n_130),
.B1(n_135),
.B2(n_136),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_79),
.C(n_81),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_134),
.C(n_138),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_132),
.A2(n_133),
.B(n_137),
.Y(n_178)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_70),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_101),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_98),
.B1(n_85),
.B2(n_83),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_85),
.B1(n_94),
.B2(n_75),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_72),
.C(n_77),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_141),
.B(n_129),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_144),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_125),
.A2(n_72),
.B1(n_84),
.B2(n_12),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_127),
.B(n_113),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_99),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_90),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_149),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_146),
.B(n_111),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_11),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_150),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_148),
.A2(n_150),
.B1(n_154),
.B2(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_103),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_113),
.B(n_14),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_151),
.B(n_105),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_16),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_153),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_16),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_122),
.A2(n_126),
.B1(n_112),
.B2(n_127),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_16),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_155),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_156),
.A2(n_166),
.B(n_175),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_122),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_126),
.B1(n_107),
.B2(n_117),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_164),
.A2(n_176),
.B1(n_143),
.B2(n_131),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_151),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_111),
.C(n_104),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_173),
.C(n_154),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_104),
.Y(n_168)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_142),
.B(n_141),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_133),
.B(n_148),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_132),
.B(n_105),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_177),
.A2(n_110),
.B1(n_114),
.B2(n_14),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_161),
.Y(n_211)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_186),
.Y(n_212)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_168),
.B(n_170),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_191),
.B1(n_193),
.B2(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

AOI22x1_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_149),
.B1(n_114),
.B2(n_146),
.Y(n_191)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_178),
.A3(n_175),
.B1(n_169),
.B2(n_176),
.C1(n_146),
.C2(n_171),
.Y(n_192)
);

OAI322xp33_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_159),
.A3(n_177),
.B1(n_173),
.B2(n_167),
.C1(n_160),
.C2(n_157),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_174),
.A2(n_140),
.B1(n_139),
.B2(n_110),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_198),
.B1(n_199),
.B2(n_166),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_196),
.Y(n_210)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_178),
.B(n_170),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_206),
.B(n_208),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_180),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_195),
.A2(n_191),
.B1(n_156),
.B2(n_187),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_204),
.B1(n_186),
.B2(n_190),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_191),
.A2(n_194),
.B1(n_184),
.B2(n_185),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_161),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_209),
.C(n_211),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_188),
.B(n_163),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_173),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_214),
.C(n_182),
.Y(n_222)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_209),
.A2(n_184),
.B1(n_199),
.B2(n_197),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_217),
.A2(n_225),
.B1(n_226),
.B2(n_207),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_220),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_189),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_219),
.B(n_223),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_208),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_224),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_181),
.B1(n_182),
.B2(n_193),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_200),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_219),
.B(n_223),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_220),
.A2(n_210),
.B1(n_206),
.B2(n_213),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_228),
.B(n_232),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_157),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_179),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_222),
.C(n_218),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_234),
.A2(n_221),
.B(n_211),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_240),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_229),
.A2(n_215),
.B(n_226),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_241),
.C(n_234),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_SL g239 ( 
.A(n_231),
.B(n_215),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_235),
.Y(n_245)
);

AOI31xp33_ASAP7_75t_SL g242 ( 
.A1(n_227),
.A2(n_162),
.A3(n_221),
.B(n_15),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_242),
.B(n_15),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_235),
.B(n_227),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_245),
.A2(n_247),
.B(n_230),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_228),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_248),
.A2(n_249),
.B(n_251),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_243),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_250),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_252),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_254),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_253),
.Y(n_256)
);


endmodule