module fake_jpeg_13336_n_582 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_582);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_582;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_11),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx5_ASAP7_75t_SL g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_15),
.B(n_13),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_60),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_63),
.B(n_66),
.Y(n_133)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_37),
.B(n_0),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_31),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_67),
.B(n_73),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_70),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_31),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_74),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_76),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_15),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_77),
.B(n_81),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_78),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_37),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_82),
.B(n_88),
.Y(n_162)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_31),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_89),
.Y(n_154)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_90),
.Y(n_168)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_91),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_94),
.B(n_97),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_96),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_24),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_24),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g153 ( 
.A(n_100),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_28),
.B(n_0),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_101),
.B(n_102),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_28),
.B(n_1),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_23),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_103),
.B(n_108),
.Y(n_160)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_23),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_18),
.B(n_1),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_2),
.Y(n_130)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_34),
.Y(n_111)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_29),
.Y(n_113)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_23),
.Y(n_115)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_35),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_116),
.B(n_53),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_20),
.Y(n_117)
);

BUFx4f_ASAP7_75t_SL g180 ( 
.A(n_117),
.Y(n_180)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_35),
.Y(n_120)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_126),
.B(n_155),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_81),
.A2(n_22),
.B(n_117),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_127),
.A2(n_169),
.B(n_60),
.C(n_69),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_130),
.B(n_141),
.Y(n_204)
);

BUFx8_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_134),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_30),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_64),
.A2(n_56),
.B1(n_47),
.B2(n_38),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_146),
.B(n_62),
.Y(n_225)
);

BUFx16f_ASAP7_75t_L g147 ( 
.A(n_60),
.Y(n_147)
);

INVx6_ASAP7_75t_SL g216 ( 
.A(n_147),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_74),
.B(n_20),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_148),
.B(n_161),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_59),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_80),
.A2(n_56),
.B1(n_54),
.B2(n_46),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_156),
.A2(n_175),
.B1(n_22),
.B2(n_78),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_84),
.B(n_42),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_70),
.B(n_30),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_173),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_98),
.A2(n_42),
.B(n_48),
.C(n_22),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_111),
.B(n_25),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_112),
.A2(n_56),
.B1(n_68),
.B2(n_57),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_153),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_114),
.B(n_25),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_49),
.Y(n_212)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_190),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_61),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_58),
.Y(n_193)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_196),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_197),
.B(n_217),
.Y(n_302)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_192),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g275 ( 
.A(n_198),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_35),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_200),
.B(n_203),
.Y(n_306)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_201),
.Y(n_278)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_202),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_48),
.Y(n_203)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_206),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_207),
.A2(n_220),
.B1(n_225),
.B2(n_230),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_146),
.A2(n_47),
.B1(n_22),
.B2(n_91),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_208),
.A2(n_209),
.B1(n_255),
.B2(n_258),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_146),
.A2(n_47),
.B1(n_118),
.B2(n_89),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g308 ( 
.A1(n_210),
.A2(n_212),
.B(n_241),
.Y(n_308)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_213),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_136),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_214),
.B(n_232),
.Y(n_282)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_128),
.Y(n_215)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_215),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_152),
.B(n_49),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_152),
.B(n_148),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_218),
.B(n_259),
.Y(n_276)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_219),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_157),
.A2(n_133),
.B1(n_167),
.B2(n_161),
.Y(n_220)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_222),
.Y(n_292)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_223),
.Y(n_274)
);

CKINVDCx12_ASAP7_75t_R g224 ( 
.A(n_134),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_224),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_129),
.Y(n_227)
);

BUFx8_ASAP7_75t_L g303 ( 
.A(n_227),
.Y(n_303)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_151),
.Y(n_228)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_158),
.Y(n_229)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_229),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_185),
.A2(n_119),
.B1(n_95),
.B2(n_93),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_231),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_136),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_133),
.A2(n_92),
.B1(n_79),
.B2(n_75),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_233),
.A2(n_240),
.B1(n_245),
.B2(n_246),
.Y(n_316)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_234),
.Y(n_293)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_122),
.Y(n_235)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_235),
.Y(n_309)
);

CKINVDCx12_ASAP7_75t_R g236 ( 
.A(n_140),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_236),
.Y(n_273)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_191),
.Y(n_237)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_237),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_129),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_243),
.Y(n_284)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_172),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_250),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_L g240 ( 
.A1(n_124),
.A2(n_71),
.B1(n_76),
.B2(n_54),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_SL g241 ( 
.A(n_137),
.B(n_52),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_167),
.B(n_50),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_242),
.B(n_248),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_160),
.B(n_33),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_135),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_244),
.B(n_249),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_159),
.A2(n_50),
.B1(n_44),
.B2(n_18),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_L g246 ( 
.A1(n_182),
.A2(n_46),
.B1(n_54),
.B2(n_33),
.Y(n_246)
);

HAxp5_ASAP7_75t_SL g247 ( 
.A(n_140),
.B(n_69),
.CON(n_247),
.SN(n_247)
);

AOI21xp33_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_254),
.B(n_180),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_150),
.B(n_44),
.Y(n_248)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_123),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_166),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_251),
.B(n_252),
.Y(n_310)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_194),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_253),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_180),
.B(n_53),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_125),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_194),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_257),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_154),
.A2(n_52),
.B1(n_51),
.B2(n_33),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_181),
.B(n_2),
.Y(n_259)
);

INVx3_ASAP7_75t_SL g260 ( 
.A(n_131),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_260),
.A2(n_263),
.B1(n_264),
.B2(n_139),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_183),
.B(n_3),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_51),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_154),
.A2(n_52),
.B1(n_51),
.B2(n_53),
.Y(n_263)
);

INVx3_ASAP7_75t_SL g264 ( 
.A(n_131),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_218),
.A2(n_261),
.B1(n_205),
.B2(n_243),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_265),
.A2(n_272),
.B1(n_297),
.B2(n_301),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_204),
.B(n_183),
.C(n_145),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_267),
.B(n_313),
.C(n_317),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_268),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_225),
.A2(n_189),
.B1(n_143),
.B2(n_132),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g358 ( 
.A1(n_269),
.A2(n_295),
.B1(n_251),
.B2(n_256),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_225),
.A2(n_210),
.B1(n_259),
.B2(n_240),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_223),
.B(n_144),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_277),
.B(n_283),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_280),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_231),
.B(n_121),
.Y(n_283)
);

OAI32xp33_ASAP7_75t_L g286 ( 
.A1(n_241),
.A2(n_189),
.A3(n_149),
.B1(n_132),
.B2(n_188),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_286),
.B(n_215),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_246),
.A2(n_143),
.B1(n_188),
.B2(n_164),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_226),
.A2(n_164),
.B1(n_142),
.B2(n_125),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_239),
.B(n_253),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_298),
.B(n_300),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_201),
.A2(n_142),
.B1(n_184),
.B2(n_149),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_260),
.A2(n_139),
.B1(n_138),
.B2(n_147),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_307),
.A2(n_312),
.B1(n_314),
.B2(n_198),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_199),
.B(n_4),
.Y(n_311)
);

AND2x2_ASAP7_75t_SL g353 ( 
.A(n_311),
.B(n_12),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_264),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_211),
.B(n_6),
.C(n_7),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_213),
.A2(n_249),
.B1(n_196),
.B2(n_255),
.Y(n_314)
);

OA22x2_ASAP7_75t_L g315 ( 
.A1(n_247),
.A2(n_7),
.B1(n_10),
.B2(n_12),
.Y(n_315)
);

NAND2x1p5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_250),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_234),
.B(n_10),
.C(n_12),
.Y(n_317)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_278),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_321),
.Y(n_385)
);

INVx2_ASAP7_75t_R g322 ( 
.A(n_308),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_322),
.B(n_331),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_302),
.B(n_235),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g397 ( 
.A(n_323),
.Y(n_397)
);

INVx8_ASAP7_75t_L g324 ( 
.A(n_266),
.Y(n_324)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_324),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_302),
.B(n_304),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_325),
.B(n_326),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_298),
.Y(n_326)
);

O2A1O1Ixp33_ASAP7_75t_L g327 ( 
.A1(n_284),
.A2(n_216),
.B(n_202),
.C(n_244),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_327),
.A2(n_350),
.B(n_352),
.Y(n_365)
);

AND2x6_ASAP7_75t_L g329 ( 
.A(n_282),
.B(n_216),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_343),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_289),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_330),
.B(n_339),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_332),
.A2(n_310),
.B(n_289),
.Y(n_380)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_271),
.Y(n_333)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

INVx8_ASAP7_75t_L g334 ( 
.A(n_266),
.Y(n_334)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_334),
.Y(n_374)
);

INVx3_ASAP7_75t_SL g336 ( 
.A(n_309),
.Y(n_336)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_336),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_296),
.Y(n_337)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_337),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_238),
.Y(n_338)
);

NAND3xp33_ASAP7_75t_L g386 ( 
.A(n_338),
.B(n_342),
.C(n_346),
.Y(n_386)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_274),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_290),
.A2(n_219),
.B1(n_206),
.B2(n_222),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_340),
.A2(n_345),
.B1(n_358),
.B2(n_360),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_273),
.B(n_227),
.Y(n_342)
);

AND2x6_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_276),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_274),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_344),
.B(n_361),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_290),
.A2(n_270),
.B1(n_316),
.B2(n_276),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_273),
.B(n_256),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_347),
.A2(n_359),
.B1(n_315),
.B2(n_305),
.Y(n_370)
);

AND2x6_ASAP7_75t_L g348 ( 
.A(n_272),
.B(n_221),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_348),
.B(n_349),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_256),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_267),
.B(n_221),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_296),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_351),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_315),
.B(n_311),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_317),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_279),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_354),
.B(n_355),
.Y(n_393)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_278),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_289),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_356),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_316),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_285),
.B(n_14),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_328),
.B(n_287),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_362),
.B(n_368),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_323),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_363),
.B(n_392),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_320),
.A2(n_300),
.B1(n_286),
.B2(n_318),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_364),
.A2(n_370),
.B1(n_378),
.B2(n_387),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_326),
.B(n_318),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_367),
.B(n_381),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_350),
.B(n_305),
.C(n_287),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_369),
.B(n_373),
.C(n_390),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_328),
.B(n_285),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_320),
.A2(n_288),
.B1(n_283),
.B2(n_277),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_380),
.B(n_322),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_357),
.B(n_299),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_341),
.A2(n_297),
.B1(n_301),
.B2(n_315),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_383),
.A2(n_347),
.B(n_275),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_331),
.A2(n_294),
.B(n_271),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_384),
.A2(n_331),
.B(n_327),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_345),
.A2(n_299),
.B1(n_309),
.B2(n_294),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_350),
.A2(n_294),
.B1(n_313),
.B2(n_293),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_389),
.A2(n_330),
.B1(n_360),
.B2(n_353),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_341),
.B(n_291),
.C(n_293),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_357),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_354),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_398),
.B(n_291),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_367),
.B(n_356),
.Y(n_400)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_400),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_396),
.Y(n_402)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_402),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_422),
.Y(n_435)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_393),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_404),
.B(n_406),
.Y(n_463)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_393),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_397),
.B(n_325),
.Y(n_407)
);

INVxp33_ASAP7_75t_L g449 ( 
.A(n_407),
.Y(n_449)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_408),
.B(n_415),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_409),
.A2(n_384),
.B(n_395),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_376),
.B(n_337),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_410),
.B(n_411),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_SL g411 ( 
.A(n_379),
.B(n_352),
.C(n_322),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_412),
.B(n_418),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_362),
.B(n_335),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_413),
.B(n_417),
.C(n_419),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_382),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_382),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_416),
.B(n_420),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_373),
.B(n_352),
.C(n_335),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_376),
.B(n_351),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_369),
.B(n_343),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_381),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_364),
.A2(n_340),
.B1(n_336),
.B2(n_351),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_421),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_388),
.Y(n_422)
);

AOI21xp33_ASAP7_75t_L g423 ( 
.A1(n_365),
.A2(n_329),
.B(n_348),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_423),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_365),
.B(n_353),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_389),
.C(n_387),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_425),
.A2(n_383),
.B1(n_391),
.B2(n_390),
.Y(n_439)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_372),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_428),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_392),
.B(n_339),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_427),
.B(n_398),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_363),
.B(n_344),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_429),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_377),
.B(n_355),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_430),
.B(n_377),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_386),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_366),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_431),
.B(n_366),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_433),
.B(n_455),
.Y(n_472)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_436),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_439),
.A2(n_458),
.B1(n_416),
.B2(n_406),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_399),
.B(n_420),
.Y(n_440)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_440),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_432),
.B(n_368),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_444),
.B(n_450),
.C(n_462),
.Y(n_476)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_446),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_399),
.B(n_378),
.Y(n_447)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_447),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_405),
.B(n_388),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_414),
.B(n_380),
.Y(n_451)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_451),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_430),
.B(n_427),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_452),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_454),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_457),
.B(n_459),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_401),
.A2(n_391),
.B1(n_375),
.B2(n_394),
.Y(n_458)
);

MAJx2_ASAP7_75t_L g459 ( 
.A(n_417),
.B(n_372),
.C(n_385),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_400),
.B(n_375),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_426),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_432),
.B(n_396),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_447),
.A2(n_401),
.B1(n_422),
.B2(n_404),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_465),
.A2(n_481),
.B1(n_439),
.B2(n_437),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_466),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_408),
.Y(n_469)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_469),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_444),
.B(n_424),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_470),
.B(n_480),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_450),
.B(n_405),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_474),
.B(n_484),
.Y(n_511)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_475),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_449),
.B(n_428),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_477),
.B(n_479),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_456),
.B(n_419),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_462),
.B(n_413),
.Y(n_480)
);

OAI22xp33_ASAP7_75t_SL g481 ( 
.A1(n_437),
.A2(n_429),
.B1(n_425),
.B2(n_414),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_441),
.B(n_409),
.Y(n_482)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_482),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_448),
.B(n_374),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_483),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_434),
.B(n_411),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_434),
.B(n_412),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_485),
.B(n_451),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_457),
.B(n_333),
.C(n_394),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_487),
.B(n_453),
.C(n_459),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_445),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_489),
.B(n_448),
.Y(n_490)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_490),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_491),
.A2(n_466),
.B1(n_478),
.B2(n_473),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_493),
.B(n_435),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_485),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_495),
.B(n_484),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_467),
.B(n_446),
.Y(n_496)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_496),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_469),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_498),
.B(n_500),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_472),
.B(n_456),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_499),
.B(n_503),
.Y(n_525)
);

INVxp33_ASAP7_75t_L g500 ( 
.A(n_482),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_486),
.B(n_455),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_471),
.B(n_445),
.Y(n_504)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_504),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_489),
.A2(n_461),
.B(n_454),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_506),
.A2(n_468),
.B(n_441),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_482),
.B(n_460),
.Y(n_508)
);

XNOR2x1_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_452),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_488),
.Y(n_509)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_509),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_510),
.B(n_474),
.C(n_464),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_512),
.A2(n_508),
.B1(n_497),
.B2(n_501),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_513),
.B(n_515),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_514),
.B(n_520),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_511),
.B(n_487),
.C(n_476),
.Y(n_515)
);

MAJx2_ASAP7_75t_L g517 ( 
.A(n_511),
.B(n_464),
.C(n_459),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_517),
.A2(n_522),
.B(n_492),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_507),
.A2(n_465),
.B1(n_458),
.B2(n_438),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_518),
.A2(n_491),
.B1(n_505),
.B2(n_506),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_495),
.B(n_470),
.C(n_480),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_519),
.B(n_527),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_526),
.B(n_443),
.Y(n_543)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_501),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_493),
.B(n_440),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_494),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_531),
.B(n_540),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_513),
.B(n_510),
.C(n_500),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_532),
.A2(n_533),
.B(n_534),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_515),
.B(n_505),
.C(n_508),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_514),
.B(n_520),
.C(n_528),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_535),
.A2(n_536),
.B1(n_523),
.B2(n_443),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_SL g536 ( 
.A1(n_529),
.A2(n_468),
.B1(n_490),
.B2(n_502),
.Y(n_536)
);

AOI21x1_ASAP7_75t_L g547 ( 
.A1(n_537),
.A2(n_516),
.B(n_517),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_521),
.Y(n_538)
);

AO21x1_ASAP7_75t_L g556 ( 
.A1(n_538),
.A2(n_453),
.B(n_371),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_512),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_539),
.B(n_541),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_518),
.A2(n_496),
.B1(n_497),
.B2(n_442),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_543),
.B(n_463),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_542),
.B(n_524),
.C(n_519),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_545),
.B(n_546),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_532),
.B(n_533),
.C(n_534),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_547),
.B(n_540),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_530),
.B(n_526),
.C(n_492),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_549),
.A2(n_554),
.B(n_371),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_544),
.B(n_525),
.Y(n_550)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_550),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_551),
.A2(n_538),
.B1(n_543),
.B2(n_535),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_530),
.B(n_463),
.C(n_435),
.Y(n_554)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_555),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_556),
.B(n_531),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_558),
.A2(n_563),
.B(n_321),
.Y(n_567)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_559),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g560 ( 
.A(n_548),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_560),
.B(n_562),
.Y(n_571)
);

CKINVDCx16_ASAP7_75t_R g564 ( 
.A(n_552),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_564),
.B(n_336),
.C(n_281),
.Y(n_570)
);

AOI322xp5_ASAP7_75t_L g566 ( 
.A1(n_557),
.A2(n_556),
.A3(n_553),
.B1(n_546),
.B2(n_554),
.C1(n_549),
.C2(n_385),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_566),
.B(n_568),
.Y(n_573)
);

AOI21x1_ASAP7_75t_L g574 ( 
.A1(n_567),
.A2(n_558),
.B(n_562),
.Y(n_574)
);

CKINVDCx14_ASAP7_75t_R g568 ( 
.A(n_561),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_570),
.B(n_324),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g572 ( 
.A(n_571),
.B(n_565),
.Y(n_572)
);

AOI322xp5_ASAP7_75t_L g576 ( 
.A1(n_572),
.A2(n_574),
.A3(n_575),
.B1(n_569),
.B2(n_568),
.C1(n_559),
.C2(n_358),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_576),
.A2(n_577),
.B(n_292),
.Y(n_578)
);

AOI322xp5_ASAP7_75t_L g577 ( 
.A1(n_573),
.A2(n_324),
.A3(n_334),
.B1(n_281),
.B2(n_292),
.C1(n_303),
.C2(n_14),
.Y(n_577)
);

BUFx24_ASAP7_75t_SL g579 ( 
.A(n_578),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_579),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_580),
.B(n_303),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g582 ( 
.A1(n_581),
.A2(n_303),
.B(n_15),
.Y(n_582)
);


endmodule