module real_aes_7374_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_1), .A2(n_136), .B(n_140), .C(n_235), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_2), .A2(n_172), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g468 ( .A(n_3), .Y(n_468) );
AOI222xp33_ASAP7_75t_L g454 ( .A1(n_4), .A2(n_455), .B1(n_736), .B2(n_739), .C1(n_742), .C2(n_743), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_5), .B(n_212), .Y(n_269) );
AOI21xp33_ASAP7_75t_L g495 ( .A1(n_6), .A2(n_172), .B(n_496), .Y(n_495) );
AND2x6_ASAP7_75t_L g136 ( .A(n_7), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g195 ( .A(n_8), .Y(n_195) );
INVx1_ASAP7_75t_L g107 ( .A(n_9), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_9), .B(n_41), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_10), .A2(n_171), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_11), .B(n_148), .Y(n_239) );
INVx1_ASAP7_75t_L g500 ( .A(n_12), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_13), .B(n_206), .Y(n_523) );
INVx1_ASAP7_75t_L g156 ( .A(n_14), .Y(n_156) );
INVx1_ASAP7_75t_L g545 ( .A(n_15), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_16), .A2(n_146), .B(n_220), .C(n_222), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_17), .B(n_212), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_18), .B(n_479), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_19), .B(n_172), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_20), .B(n_185), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_21), .A2(n_206), .B(n_207), .C(n_209), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_22), .B(n_212), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_23), .B(n_148), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_24), .A2(n_180), .B(n_222), .C(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_25), .B(n_148), .Y(n_147) );
CKINVDCx16_ASAP7_75t_R g252 ( .A(n_26), .Y(n_252) );
INVx1_ASAP7_75t_L g144 ( .A(n_27), .Y(n_144) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_28), .A2(n_102), .B1(n_113), .B2(n_746), .Y(n_101) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_29), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_30), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_31), .B(n_148), .Y(n_469) );
INVx1_ASAP7_75t_L g178 ( .A(n_32), .Y(n_178) );
INVx1_ASAP7_75t_L g490 ( .A(n_33), .Y(n_490) );
INVx2_ASAP7_75t_L g134 ( .A(n_34), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_35), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_36), .A2(n_206), .B(n_265), .C(n_267), .Y(n_264) );
INVxp67_ASAP7_75t_L g179 ( .A(n_37), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_38), .A2(n_140), .B(n_143), .C(n_151), .Y(n_139) );
CKINVDCx14_ASAP7_75t_R g263 ( .A(n_39), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_40), .A2(n_136), .B(n_140), .C(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_41), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g489 ( .A(n_42), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_43), .A2(n_193), .B(n_194), .C(n_196), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_44), .B(n_148), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_45), .A2(n_48), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_45), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_46), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_47), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_48), .Y(n_122) );
INVx1_ASAP7_75t_L g204 ( .A(n_49), .Y(n_204) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_50), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_51), .B(n_172), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_52), .A2(n_140), .B1(n_209), .B2(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_53), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g465 ( .A(n_54), .Y(n_465) );
CKINVDCx14_ASAP7_75t_R g191 ( .A(n_55), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_56), .A2(n_193), .B(n_267), .C(n_499), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_57), .Y(n_538) );
INVx1_ASAP7_75t_L g497 ( .A(n_58), .Y(n_497) );
INVx1_ASAP7_75t_L g137 ( .A(n_59), .Y(n_137) );
INVx1_ASAP7_75t_L g155 ( .A(n_60), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_61), .A2(n_90), .B1(n_737), .B2(n_738), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_61), .Y(n_737) );
INVx1_ASAP7_75t_SL g266 ( .A(n_62), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_63), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_64), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_65), .B(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g255 ( .A(n_66), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_SL g478 ( .A1(n_67), .A2(n_267), .B(n_479), .C(n_480), .Y(n_478) );
INVxp67_ASAP7_75t_L g481 ( .A(n_68), .Y(n_481) );
INVx1_ASAP7_75t_L g112 ( .A(n_69), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_70), .A2(n_172), .B(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_71), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_72), .A2(n_172), .B(n_217), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_73), .Y(n_493) );
INVx1_ASAP7_75t_L g532 ( .A(n_74), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_75), .A2(n_171), .B(n_173), .Y(n_170) );
CKINVDCx16_ASAP7_75t_R g138 ( .A(n_76), .Y(n_138) );
INVx1_ASAP7_75t_L g218 ( .A(n_77), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_78), .A2(n_136), .B(n_140), .C(n_534), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_79), .A2(n_172), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g221 ( .A(n_80), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_81), .B(n_145), .Y(n_514) );
INVx2_ASAP7_75t_L g153 ( .A(n_82), .Y(n_153) );
INVx1_ASAP7_75t_L g236 ( .A(n_83), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_84), .B(n_479), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_85), .A2(n_136), .B(n_140), .C(n_467), .Y(n_466) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_86), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g445 ( .A(n_86), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g733 ( .A(n_86), .Y(n_733) );
OR2x2_ASAP7_75t_L g735 ( .A(n_86), .B(n_447), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_87), .A2(n_140), .B(n_254), .C(n_257), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_88), .B(n_152), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_89), .Y(n_472) );
CKINVDCx14_ASAP7_75t_R g738 ( .A(n_90), .Y(n_738) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_91), .A2(n_136), .B(n_140), .C(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_92), .Y(n_527) );
INVx1_ASAP7_75t_L g477 ( .A(n_93), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g542 ( .A(n_94), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_95), .B(n_145), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_96), .B(n_160), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_97), .B(n_160), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g208 ( .A(n_99), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_100), .A2(n_172), .B(n_476), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx5_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
CKINVDCx9p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
BUFx4f_ASAP7_75t_SL g746 ( .A(n_105), .Y(n_746) );
OR2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
AND2x2_ASAP7_75t_L g447 ( .A(n_109), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_453), .Y(n_113) );
BUFx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g745 ( .A(n_117), .Y(n_745) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_442), .B(n_449), .Y(n_119) );
XNOR2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_124), .Y(n_120) );
INVx1_ASAP7_75t_SL g734 ( .A(n_124), .Y(n_734) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_124), .A2(n_457), .B1(n_730), .B2(n_740), .Y(n_739) );
OR5x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_336), .C(n_400), .D(n_416), .E(n_431), .Y(n_124) );
NAND4xp25_ASAP7_75t_L g125 ( .A(n_126), .B(n_270), .C(n_297), .D(n_320), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_213), .B(n_224), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_162), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx3_ASAP7_75t_SL g247 ( .A(n_129), .Y(n_247) );
AND2x4_ASAP7_75t_L g283 ( .A(n_129), .B(n_272), .Y(n_283) );
OR2x2_ASAP7_75t_L g293 ( .A(n_129), .B(n_249), .Y(n_293) );
OR2x2_ASAP7_75t_L g339 ( .A(n_129), .B(n_165), .Y(n_339) );
AND2x2_ASAP7_75t_L g353 ( .A(n_129), .B(n_248), .Y(n_353) );
AND2x2_ASAP7_75t_L g396 ( .A(n_129), .B(n_286), .Y(n_396) );
AND2x2_ASAP7_75t_L g403 ( .A(n_129), .B(n_260), .Y(n_403) );
AND2x2_ASAP7_75t_L g422 ( .A(n_129), .B(n_312), .Y(n_422) );
AND2x2_ASAP7_75t_L g440 ( .A(n_129), .B(n_282), .Y(n_440) );
OR2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_157), .Y(n_129) );
O2A1O1Ixp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_138), .B(n_139), .C(n_152), .Y(n_130) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_131), .A2(n_233), .B(n_234), .Y(n_232) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_131), .A2(n_252), .B(n_253), .Y(n_251) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_131), .A2(n_465), .B(n_466), .Y(n_464) );
OAI22xp33_ASAP7_75t_L g486 ( .A1(n_131), .A2(n_182), .B1(n_487), .B2(n_491), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_131), .A2(n_532), .B(n_533), .Y(n_531) );
NAND2x1p5_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
AND2x4_ASAP7_75t_L g172 ( .A(n_132), .B(n_136), .Y(n_172) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx1_ASAP7_75t_L g150 ( .A(n_133), .Y(n_150) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g141 ( .A(n_134), .Y(n_141) );
INVx1_ASAP7_75t_L g210 ( .A(n_134), .Y(n_210) );
INVx1_ASAP7_75t_L g142 ( .A(n_135), .Y(n_142) );
INVx3_ASAP7_75t_L g146 ( .A(n_135), .Y(n_146) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_135), .Y(n_148) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_135), .Y(n_181) );
INVx1_ASAP7_75t_L g479 ( .A(n_135), .Y(n_479) );
BUFx3_ASAP7_75t_L g151 ( .A(n_136), .Y(n_151) );
INVx4_ASAP7_75t_SL g182 ( .A(n_136), .Y(n_182) );
INVx5_ASAP7_75t_L g175 ( .A(n_140), .Y(n_175) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
BUFx3_ASAP7_75t_L g197 ( .A(n_141), .Y(n_197) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_141), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_147), .C(n_149), .Y(n_143) );
OAI22xp33_ASAP7_75t_L g177 ( .A1(n_145), .A2(n_178), .B1(n_179), .B2(n_180), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_145), .A2(n_468), .B(n_469), .C(n_470), .Y(n_467) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_146), .B(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_146), .B(n_481), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_146), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g193 ( .A(n_148), .Y(n_193) );
INVx4_ASAP7_75t_L g206 ( .A(n_148), .Y(n_206) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_150), .B(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_152), .A2(n_189), .B(n_198), .Y(n_188) );
INVx1_ASAP7_75t_L g231 ( .A(n_152), .Y(n_231) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_152), .A2(n_540), .B(n_546), .Y(n_539) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AND2x2_ASAP7_75t_L g161 ( .A(n_153), .B(n_154), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
INVx3_ASAP7_75t_L g212 ( .A(n_159), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_159), .B(n_242), .Y(n_241) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_159), .A2(n_251), .B(n_258), .Y(n_250) );
NOR2xp33_ASAP7_75t_SL g516 ( .A(n_159), .B(n_517), .Y(n_516) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_160), .Y(n_201) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_160), .A2(n_475), .B(n_482), .Y(n_474) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g168 ( .A(n_161), .Y(n_168) );
INVx1_ASAP7_75t_L g405 ( .A(n_162), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_187), .Y(n_162) );
AND2x2_ASAP7_75t_L g315 ( .A(n_163), .B(n_248), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_163), .B(n_335), .Y(n_334) );
AOI32xp33_ASAP7_75t_L g348 ( .A1(n_163), .A2(n_349), .A3(n_352), .B1(n_354), .B2(n_358), .Y(n_348) );
AND2x2_ASAP7_75t_L g418 ( .A(n_163), .B(n_312), .Y(n_418) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g282 ( .A(n_165), .B(n_249), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_165), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g324 ( .A(n_165), .B(n_271), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_165), .B(n_403), .Y(n_402) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_169), .B(n_183), .Y(n_165) );
INVx1_ASAP7_75t_L g287 ( .A(n_166), .Y(n_287) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_166), .A2(n_531), .B(n_537), .Y(n_530) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_SL g510 ( .A1(n_167), .A2(n_511), .B(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AO21x2_ASAP7_75t_L g463 ( .A1(n_168), .A2(n_464), .B(n_471), .Y(n_463) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_168), .A2(n_486), .B(n_492), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_168), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OA21x2_ASAP7_75t_L g286 ( .A1(n_170), .A2(n_184), .B(n_287), .Y(n_286) );
BUFx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_175), .B(n_176), .C(n_182), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_SL g190 ( .A1(n_175), .A2(n_182), .B(n_191), .C(n_192), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_SL g203 ( .A1(n_175), .A2(n_182), .B(n_204), .C(n_205), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_SL g217 ( .A1(n_175), .A2(n_182), .B(n_218), .C(n_219), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_175), .A2(n_182), .B(n_263), .C(n_264), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_175), .A2(n_182), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_175), .A2(n_182), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_175), .A2(n_182), .B(n_542), .C(n_543), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_180), .B(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_180), .B(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_180), .B(n_545), .Y(n_544) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g238 ( .A(n_181), .Y(n_238) );
OAI22xp5_ASAP7_75t_SL g488 ( .A1(n_181), .A2(n_238), .B1(n_489), .B2(n_490), .Y(n_488) );
INVx1_ASAP7_75t_L g257 ( .A(n_182), .Y(n_257) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_186), .B(n_259), .Y(n_258) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_186), .A2(n_519), .B(n_526), .Y(n_518) );
AND2x2_ASAP7_75t_L g289 ( .A(n_187), .B(n_228), .Y(n_289) );
AND2x2_ASAP7_75t_L g365 ( .A(n_187), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g437 ( .A(n_187), .Y(n_437) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_199), .Y(n_187) );
OR2x2_ASAP7_75t_L g227 ( .A(n_188), .B(n_200), .Y(n_227) );
AND2x2_ASAP7_75t_L g244 ( .A(n_188), .B(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_188), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g296 ( .A(n_188), .Y(n_296) );
AND2x2_ASAP7_75t_L g323 ( .A(n_188), .B(n_200), .Y(n_323) );
BUFx3_ASAP7_75t_L g326 ( .A(n_188), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_188), .B(n_301), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_188), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g240 ( .A(n_196), .Y(n_240) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g222 ( .A(n_197), .Y(n_222) );
INVx2_ASAP7_75t_L g277 ( .A(n_199), .Y(n_277) );
AND2x2_ASAP7_75t_L g295 ( .A(n_199), .B(n_275), .Y(n_295) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g306 ( .A(n_200), .B(n_215), .Y(n_306) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_200), .Y(n_319) );
OA21x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_211), .Y(n_200) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_201), .A2(n_216), .B(n_223), .Y(n_215) );
OA21x2_ASAP7_75t_L g260 ( .A1(n_201), .A2(n_261), .B(n_269), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_206), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g470 ( .A(n_209), .Y(n_470) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_212), .A2(n_495), .B(n_501), .Y(n_494) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_214), .B(n_326), .Y(n_376) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_SL g245 ( .A(n_215), .Y(n_245) );
NAND3xp33_ASAP7_75t_L g294 ( .A(n_215), .B(n_295), .C(n_296), .Y(n_294) );
OR2x2_ASAP7_75t_L g302 ( .A(n_215), .B(n_275), .Y(n_302) );
AND2x2_ASAP7_75t_L g322 ( .A(n_215), .B(n_275), .Y(n_322) );
AND2x2_ASAP7_75t_L g366 ( .A(n_215), .B(n_230), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_243), .B(n_246), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_226), .B(n_228), .Y(n_225) );
AND2x2_ASAP7_75t_L g441 ( .A(n_226), .B(n_366), .Y(n_441) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_227), .A2(n_339), .B1(n_381), .B2(n_383), .Y(n_380) );
OR2x2_ASAP7_75t_L g387 ( .A(n_227), .B(n_302), .Y(n_387) );
OR2x2_ASAP7_75t_L g411 ( .A(n_227), .B(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_227), .B(n_331), .Y(n_424) );
AND2x2_ASAP7_75t_L g317 ( .A(n_228), .B(n_318), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_228), .A2(n_390), .B(n_405), .Y(n_404) );
AOI32xp33_ASAP7_75t_L g425 ( .A1(n_228), .A2(n_315), .A3(n_426), .B1(n_428), .B2(n_429), .Y(n_425) );
OR2x2_ASAP7_75t_L g436 ( .A(n_228), .B(n_437), .Y(n_436) );
CKINVDCx16_ASAP7_75t_R g228 ( .A(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g304 ( .A(n_229), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_229), .B(n_318), .Y(n_383) );
BUFx3_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx4_ASAP7_75t_L g275 ( .A(n_230), .Y(n_275) );
AND2x2_ASAP7_75t_L g341 ( .A(n_230), .B(n_306), .Y(n_341) );
AND3x2_ASAP7_75t_L g350 ( .A(n_230), .B(n_244), .C(n_351), .Y(n_350) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_241), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_231), .B(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_231), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_231), .B(n_538), .Y(n_537) );
O2A1O1Ixp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_239), .C(n_240), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_237), .A2(n_240), .B(n_255), .C(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_240), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_240), .A2(n_535), .B(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g276 ( .A(n_245), .B(n_277), .Y(n_276) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_245), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_245), .B(n_275), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
AND2x2_ASAP7_75t_L g271 ( .A(n_247), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g311 ( .A(n_247), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g329 ( .A(n_247), .B(n_260), .Y(n_329) );
AND2x2_ASAP7_75t_L g347 ( .A(n_247), .B(n_249), .Y(n_347) );
OR2x2_ASAP7_75t_L g361 ( .A(n_247), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g407 ( .A(n_247), .B(n_335), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_248), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_260), .Y(n_248) );
AND2x2_ASAP7_75t_L g308 ( .A(n_249), .B(n_286), .Y(n_308) );
OR2x2_ASAP7_75t_L g362 ( .A(n_249), .B(n_286), .Y(n_362) );
AND2x2_ASAP7_75t_L g415 ( .A(n_249), .B(n_272), .Y(n_415) );
INVx2_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
BUFx2_ASAP7_75t_L g313 ( .A(n_250), .Y(n_313) );
AND2x2_ASAP7_75t_L g335 ( .A(n_250), .B(n_260), .Y(n_335) );
INVx2_ASAP7_75t_L g272 ( .A(n_260), .Y(n_272) );
INVx1_ASAP7_75t_L g292 ( .A(n_260), .Y(n_292) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_268), .Y(n_524) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_273), .B(n_278), .C(n_290), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_271), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g434 ( .A(n_271), .Y(n_434) );
AND2x2_ASAP7_75t_L g312 ( .A(n_272), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_275), .B(n_276), .Y(n_284) );
INVx1_ASAP7_75t_L g369 ( .A(n_275), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_275), .B(n_296), .Y(n_393) );
AND2x2_ASAP7_75t_L g409 ( .A(n_275), .B(n_323), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_276), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g300 ( .A(n_277), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_284), .B1(n_285), .B2(n_288), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_281), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_282), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g307 ( .A(n_283), .B(n_308), .Y(n_307) );
AOI221xp5_ASAP7_75t_SL g372 ( .A1(n_283), .A2(n_325), .B1(n_373), .B2(n_378), .C(n_380), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_283), .B(n_346), .Y(n_379) );
INVx1_ASAP7_75t_L g439 ( .A(n_285), .Y(n_439) );
BUFx3_ASAP7_75t_L g346 ( .A(n_286), .Y(n_346) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AOI21xp33_ASAP7_75t_SL g290 ( .A1(n_291), .A2(n_293), .B(n_294), .Y(n_290) );
INVx1_ASAP7_75t_L g355 ( .A(n_292), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_292), .B(n_346), .Y(n_399) );
INVx1_ASAP7_75t_L g356 ( .A(n_293), .Y(n_356) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_293), .B(n_346), .Y(n_357) );
INVxp67_ASAP7_75t_L g377 ( .A(n_295), .Y(n_377) );
AND2x2_ASAP7_75t_L g318 ( .A(n_296), .B(n_319), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_303), .B(n_307), .C(n_309), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_SL g332 ( .A(n_300), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_301), .B(n_332), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_301), .B(n_323), .Y(n_374) );
INVx2_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_304), .A2(n_310), .B1(n_314), .B2(n_316), .Y(n_309) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g325 ( .A(n_306), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g370 ( .A(n_306), .B(n_371), .Y(n_370) );
OAI21xp33_ASAP7_75t_L g373 ( .A1(n_308), .A2(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_312), .A2(n_321), .B1(n_324), .B2(n_325), .C(n_327), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_312), .B(n_346), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_312), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g428 ( .A(n_318), .Y(n_428) );
INVxp67_ASAP7_75t_L g351 ( .A(n_319), .Y(n_351) );
INVx1_ASAP7_75t_L g358 ( .A(n_321), .Y(n_358) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x2_ASAP7_75t_L g397 ( .A(n_322), .B(n_326), .Y(n_397) );
INVx1_ASAP7_75t_L g371 ( .A(n_326), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_326), .B(n_341), .Y(n_401) );
OAI32xp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_330), .A3(n_332), .B1(n_333), .B2(n_334), .Y(n_327) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_SL g340 ( .A(n_335), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_335), .B(n_367), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_335), .B(n_396), .Y(n_427) );
NAND2x1p5_ASAP7_75t_L g435 ( .A(n_335), .B(n_346), .Y(n_435) );
NAND5xp2_ASAP7_75t_L g336 ( .A(n_337), .B(n_359), .C(n_372), .D(n_384), .E(n_385), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_341), .B1(n_342), .B2(n_344), .C(n_348), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp33_ASAP7_75t_SL g363 ( .A(n_343), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_346), .B(n_415), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_347), .A2(n_360), .B1(n_363), .B2(n_367), .Y(n_359) );
INVx2_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
OAI211xp5_ASAP7_75t_SL g354 ( .A1(n_350), .A2(n_355), .B(n_356), .C(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_SL g382 ( .A(n_362), .Y(n_382) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_371), .B(n_420), .Y(n_430) );
OR2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI222xp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_388), .B1(n_390), .B2(n_394), .C1(n_397), .C2(n_398), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_404), .B2(n_406), .C(n_408), .Y(n_400) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
OAI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B(n_413), .Y(n_408) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g420 ( .A(n_412), .Y(n_420) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .B1(n_421), .B2(n_423), .C(n_425), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
A2O1A1Ixp33_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_435), .B(n_436), .C(n_438), .Y(n_431) );
INVxp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI21xp33_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g452 ( .A(n_445), .Y(n_452) );
NOR2x2_ASAP7_75t_L g743 ( .A(n_446), .B(n_733), .Y(n_743) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g732 ( .A(n_447), .B(n_733), .Y(n_732) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_449), .B(n_454), .C(n_744), .Y(n_453) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_456), .A2(n_730), .B1(n_734), .B2(n_735), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR4x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_619), .C(n_679), .D(n_706), .Y(n_457) );
NAND4xp25_ASAP7_75t_SL g458 ( .A(n_459), .B(n_567), .C(n_598), .D(n_615), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_502), .B(n_504), .C(n_547), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_483), .Y(n_460) );
INVx1_ASAP7_75t_L g609 ( .A(n_461), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_461), .A2(n_650), .B1(n_698), .B2(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_473), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_462), .B(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g560 ( .A(n_462), .B(n_485), .Y(n_560) );
AND2x2_ASAP7_75t_L g602 ( .A(n_462), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_462), .B(n_503), .Y(n_614) );
INVx1_ASAP7_75t_L g654 ( .A(n_462), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_462), .B(n_708), .Y(n_707) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g582 ( .A(n_463), .B(n_485), .Y(n_582) );
INVx3_ASAP7_75t_L g586 ( .A(n_463), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_463), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g673 ( .A(n_473), .B(n_494), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_473), .B(n_586), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_473), .B(n_701), .Y(n_700) );
INVx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g503 ( .A(n_474), .B(n_485), .Y(n_503) );
INVx1_ASAP7_75t_L g555 ( .A(n_474), .Y(n_555) );
BUFx2_ASAP7_75t_L g559 ( .A(n_474), .Y(n_559) );
AND2x2_ASAP7_75t_L g603 ( .A(n_474), .B(n_484), .Y(n_603) );
OR2x2_ASAP7_75t_L g642 ( .A(n_474), .B(n_484), .Y(n_642) );
AND2x2_ASAP7_75t_L g667 ( .A(n_474), .B(n_494), .Y(n_667) );
AND2x2_ASAP7_75t_L g726 ( .A(n_474), .B(n_556), .Y(n_726) );
INVx1_ASAP7_75t_L g701 ( .A(n_483), .Y(n_701) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_494), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_484), .B(n_494), .Y(n_587) );
AND2x2_ASAP7_75t_L g597 ( .A(n_484), .B(n_586), .Y(n_597) );
BUFx2_ASAP7_75t_L g608 ( .A(n_484), .Y(n_608) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g630 ( .A(n_485), .B(n_494), .Y(n_630) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_485), .Y(n_685) );
AND2x2_ASAP7_75t_SL g502 ( .A(n_494), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_SL g556 ( .A(n_494), .Y(n_556) );
BUFx2_ASAP7_75t_L g581 ( .A(n_494), .Y(n_581) );
INVx2_ASAP7_75t_L g600 ( .A(n_494), .Y(n_600) );
AND2x2_ASAP7_75t_L g662 ( .A(n_494), .B(n_586), .Y(n_662) );
AOI321xp33_ASAP7_75t_L g681 ( .A1(n_502), .A2(n_682), .A3(n_683), .B1(n_684), .B2(n_686), .C(n_687), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_503), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_503), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g675 ( .A(n_503), .B(n_654), .Y(n_675) );
AND2x2_ASAP7_75t_L g708 ( .A(n_503), .B(n_600), .Y(n_708) );
INVx1_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_528), .Y(n_505) );
OR2x2_ASAP7_75t_L g610 ( .A(n_506), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_518), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx3_ASAP7_75t_L g562 ( .A(n_509), .Y(n_562) );
AND2x2_ASAP7_75t_L g572 ( .A(n_509), .B(n_530), .Y(n_572) );
AND2x2_ASAP7_75t_L g577 ( .A(n_509), .B(n_552), .Y(n_577) );
INVx1_ASAP7_75t_L g594 ( .A(n_509), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_509), .B(n_575), .Y(n_613) );
AND2x2_ASAP7_75t_L g618 ( .A(n_509), .B(n_551), .Y(n_618) );
OR2x2_ASAP7_75t_L g650 ( .A(n_509), .B(n_639), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_509), .B(n_563), .Y(n_689) );
AND2x2_ASAP7_75t_L g723 ( .A(n_509), .B(n_549), .Y(n_723) );
OR2x6_ASAP7_75t_L g509 ( .A(n_510), .B(n_516), .Y(n_509) );
INVx1_ASAP7_75t_L g550 ( .A(n_518), .Y(n_550) );
INVx2_ASAP7_75t_L g565 ( .A(n_518), .Y(n_565) );
AND2x2_ASAP7_75t_L g605 ( .A(n_518), .B(n_576), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_518), .B(n_552), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_525), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_524), .Y(n_521) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g711 ( .A(n_529), .B(n_562), .Y(n_711) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_539), .Y(n_529) );
INVx2_ASAP7_75t_L g552 ( .A(n_530), .Y(n_552) );
AND2x2_ASAP7_75t_L g705 ( .A(n_530), .B(n_565), .Y(n_705) );
AND2x2_ASAP7_75t_L g551 ( .A(n_539), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g566 ( .A(n_539), .Y(n_566) );
INVx1_ASAP7_75t_L g576 ( .A(n_539), .Y(n_576) );
OAI22xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_553), .B1(n_557), .B2(n_561), .Y(n_547) );
OAI22xp33_ASAP7_75t_L g702 ( .A1(n_548), .A2(n_666), .B1(n_703), .B2(n_704), .Y(n_702) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g617 ( .A(n_550), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_551), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g612 ( .A(n_552), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_552), .B(n_565), .Y(n_639) );
INVx1_ASAP7_75t_L g655 ( .A(n_552), .Y(n_655) );
AND2x2_ASAP7_75t_L g596 ( .A(n_554), .B(n_597), .Y(n_596) );
INVx3_ASAP7_75t_SL g635 ( .A(n_554), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_554), .B(n_560), .Y(n_712) );
AND2x4_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g721 ( .A(n_557), .Y(n_721) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_558), .B(n_654), .Y(n_696) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx3_ASAP7_75t_SL g601 ( .A(n_560), .Y(n_601) );
NAND2x1_ASAP7_75t_SL g561 ( .A(n_562), .B(n_563), .Y(n_561) );
AND2x2_ASAP7_75t_L g622 ( .A(n_562), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g629 ( .A(n_562), .B(n_566), .Y(n_629) );
AND2x2_ASAP7_75t_L g634 ( .A(n_562), .B(n_575), .Y(n_634) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_562), .Y(n_683) );
OAI311xp33_ASAP7_75t_L g706 ( .A1(n_563), .A2(n_707), .A3(n_709), .B1(n_710), .C1(n_720), .Y(n_706) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g719 ( .A(n_564), .B(n_592), .Y(n_719) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AND2x2_ASAP7_75t_L g575 ( .A(n_565), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g623 ( .A(n_565), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g678 ( .A(n_565), .Y(n_678) );
INVx1_ASAP7_75t_L g571 ( .A(n_566), .Y(n_571) );
INVx1_ASAP7_75t_L g591 ( .A(n_566), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_566), .B(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g624 ( .A(n_566), .Y(n_624) );
AOI221xp5_ASAP7_75t_SL g567 ( .A1(n_568), .A2(n_570), .B1(n_578), .B2(n_583), .C(n_588), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_573), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx4_ASAP7_75t_L g592 ( .A(n_572), .Y(n_592) );
AND2x2_ASAP7_75t_L g686 ( .A(n_572), .B(n_605), .Y(n_686) );
AND2x2_ASAP7_75t_L g693 ( .A(n_572), .B(n_575), .Y(n_693) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_575), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g604 ( .A(n_577), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_580), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g729 ( .A(n_582), .B(n_673), .Y(n_729) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g714 ( .A(n_586), .B(n_642), .Y(n_714) );
OAI211xp5_ASAP7_75t_L g679 ( .A1(n_587), .A2(n_680), .B(n_681), .C(n_694), .Y(n_679) );
AOI21xp33_ASAP7_75t_SL g588 ( .A1(n_589), .A2(n_593), .B(n_595), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NOR2xp67_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g658 ( .A(n_592), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g687 ( .A1(n_593), .A2(n_688), .B1(n_689), .B2(n_690), .C(n_691), .Y(n_687) );
AND2x2_ASAP7_75t_L g664 ( .A(n_594), .B(n_605), .Y(n_664) );
AND2x2_ASAP7_75t_L g717 ( .A(n_594), .B(n_612), .Y(n_717) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_597), .B(n_635), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_602), .B(n_604), .C(n_606), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
AND2x2_ASAP7_75t_L g645 ( .A(n_600), .B(n_603), .Y(n_645) );
OR2x2_ASAP7_75t_L g688 ( .A(n_600), .B(n_642), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_601), .B(n_667), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_601), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g632 ( .A(n_602), .Y(n_632) );
INVx1_ASAP7_75t_L g698 ( .A(n_605), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_610), .B1(n_613), .B2(n_614), .Y(n_606) );
INVx1_ASAP7_75t_L g621 ( .A(n_607), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_608), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g684 ( .A(n_609), .B(n_685), .Y(n_684) );
INVxp67_ASAP7_75t_L g670 ( .A(n_611), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_612), .B(n_698), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g671 ( .A1(n_613), .A2(n_672), .B1(n_674), .B2(n_676), .Y(n_671) );
INVx1_ASAP7_75t_L g680 ( .A(n_616), .Y(n_680) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AND2x2_ASAP7_75t_L g722 ( .A(n_617), .B(n_717), .Y(n_722) );
AOI222xp33_ASAP7_75t_L g651 ( .A1(n_618), .A2(n_652), .B1(n_655), .B2(n_656), .C1(n_659), .C2(n_660), .Y(n_651) );
NAND4xp25_ASAP7_75t_SL g619 ( .A(n_620), .B(n_640), .C(n_651), .D(n_663), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_625), .B2(n_630), .C(n_631), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_623), .B(n_658), .Y(n_657) );
INVxp67_ASAP7_75t_L g649 ( .A(n_624), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_625), .A2(n_695), .B1(n_697), .B2(n_699), .C(n_702), .Y(n_694) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g637 ( .A(n_629), .B(n_638), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g691 ( .A1(n_630), .A2(n_692), .B(n_693), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B1(n_635), .B2(n_636), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B(n_646), .Y(n_640) );
INVxp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g682 ( .A(n_653), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_654), .B(n_673), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_654), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_658), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g690 ( .A(n_662), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_668), .B2(n_670), .C(n_671), .Y(n_663) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI222xp33_ASAP7_75t_L g710 ( .A1(n_673), .A2(n_711), .B1(n_712), .B2(n_713), .C1(n_715), .C2(n_718), .Y(n_710) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_677), .B(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g709 ( .A(n_683), .Y(n_709) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVxp33_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_723), .B2(n_724), .C(n_727), .Y(n_720) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g741 ( .A(n_735), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_736), .Y(n_742) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
endmodule