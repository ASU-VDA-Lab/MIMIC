module fake_jpeg_31714_n_76 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_75;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_14),
.B(n_2),
.Y(n_21)
);

OAI21xp33_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_15),
.B(n_19),
.Y(n_33)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_17),
.Y(n_24)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_28),
.Y(n_29)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_10),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

AO22x1_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_30),
.A2(n_37),
.B1(n_38),
.B2(n_28),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_15),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_12),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_27),
.C(n_23),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_49),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_12),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_48),
.B(n_31),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_13),
.B1(n_18),
.B2(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_37),
.Y(n_49)
);

NOR3xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_34),
.C(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_16),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_39),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_44),
.C(n_10),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_11),
.B1(n_34),
.B2(n_8),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_49),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_60),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_47),
.B(n_48),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_61),
.B(n_62),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_9),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_63),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_SL g69 ( 
.A1(n_67),
.A2(n_50),
.B(n_60),
.C(n_53),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_69),
.B(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_52),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_67),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_57),
.C(n_9),
.Y(n_75)
);

MAJx2_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_73),
.C(n_11),
.Y(n_76)
);


endmodule