module real_jpeg_6752_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_205;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx8_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_1),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_2),
.B(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_2),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_2),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_2),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_3),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_3),
.B(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_3),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_4),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_4),
.B(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_4),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_4),
.A2(n_138),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_4),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_4),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_4),
.B(n_186),
.Y(n_212)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_5),
.Y(n_139)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_7),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_7),
.B(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_7),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_7),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_7),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_7),
.B(n_174),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_7),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_8),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_9),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_9),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_9),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_9),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_10),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_10),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_10),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_10),
.B(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_10),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_11),
.Y(n_137)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_13),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_14),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_14),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_14),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_15),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_15),
.B(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_15),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_161),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_160),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_20),
.B(n_106),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_67),
.C(n_89),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_21),
.B(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_39),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_22),
.B(n_50),
.C(n_66),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_24),
.B(n_30),
.C(n_34),
.Y(n_130)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_28),
.Y(n_153)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_28),
.Y(n_177)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_32),
.Y(n_192)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_38),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_50),
.B1(n_65),
.B2(n_66),
.Y(n_39)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_41),
.B(n_47),
.Y(n_128)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_45),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_48),
.Y(n_182)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_48),
.Y(n_203)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_49),
.Y(n_211)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.C(n_60),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_51),
.A2(n_52),
.B1(n_60),
.B2(n_61),
.Y(n_227)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_56),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_57),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_58),
.Y(n_196)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_67),
.A2(n_89),
.B1(n_90),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_67),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_77),
.B1(n_78),
.B2(n_88),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_72),
.B2(n_76),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_69),
.B(n_76),
.C(n_77),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_83),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_83),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_83),
.Y(n_98)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_87),
.Y(n_205)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_90),
.B(n_224),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_90),
.B(n_225),
.C(n_226),
.Y(n_233)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_96),
.CI(n_99),
.CON(n_90),
.SN(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_100),
.A2(n_102),
.B1(n_103),
.B2(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_100),
.Y(n_188)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_131),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_126),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_125),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_159),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_144),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_138),
.B(n_142),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_135),
.B(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_155),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_150),
.B1(n_151),
.B2(n_154),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_146),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_229),
.B(n_234),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_221),
.B(n_228),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_197),
.B(n_220),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_189),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_165),
.B(n_189),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_178),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_166),
.B(n_179),
.C(n_187),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_172),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_167),
.B(n_173),
.C(n_175),
.Y(n_225)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_187),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_183),
.Y(n_190)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.C(n_193),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_193),
.B1(n_194),
.B2(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_214),
.B(n_219),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_207),
.B(n_213),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_206),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_206),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_204),
.Y(n_215)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_216),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_223),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_233),
.Y(n_234)
);


endmodule