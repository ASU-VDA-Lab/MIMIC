module fake_ariane_3196_n_111 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_10, n_111);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_111;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_40;
wire n_106;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_109;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_108;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVxp67_ASAP7_75t_SL g21 ( 
.A(n_18),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_1),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_32),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_21),
.Y(n_49)
);

AO22x2_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_47),
.B1(n_36),
.B2(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

AOI22x1_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

AND2x6_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_25),
.Y(n_57)
);

AOI222xp33_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_39),
.B1(n_44),
.B2(n_47),
.C1(n_41),
.C2(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_38),
.B(n_29),
.C(n_27),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_38),
.B(n_39),
.C(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_37),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_43),
.Y(n_63)
);

OAI21x1_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_51),
.B(n_56),
.Y(n_64)
);

AND2x4_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_57),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_45),
.B1(n_57),
.B2(n_50),
.Y(n_66)
);

OAI21x1_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_51),
.B(n_54),
.Y(n_67)
);

OAI21x1_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_57),
.B(n_50),
.Y(n_68)
);

OAI21x1_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_57),
.B(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

OR2x6_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_63),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_61),
.B1(n_45),
.B2(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_65),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_65),
.B1(n_68),
.B2(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

AND2x4_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_70),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NOR2xp67_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_72),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_75),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_76),
.C(n_70),
.Y(n_88)
);

OAI332xp33_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_7),
.B3(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_75),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_67),
.B(n_68),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_88),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

NAND5xp2_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_89),
.C(n_76),
.D(n_75),
.E(n_9),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_4),
.B(n_7),
.C(n_8),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_97),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_95),
.B1(n_78),
.B2(n_67),
.Y(n_103)
);

AND2x4_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_78),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_102),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_R g106 ( 
.A(n_104),
.B(n_99),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_103),
.B1(n_98),
.B2(n_106),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_108),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_101),
.B1(n_78),
.B2(n_24),
.Y(n_110)
);

AOI221xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_19),
.B1(n_24),
.B2(n_46),
.C(n_109),
.Y(n_111)
);


endmodule