module fake_jpeg_11512_n_540 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_540);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_540;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_56),
.Y(n_146)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_58),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_59),
.Y(n_169)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_60),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_27),
.B(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_62),
.B(n_63),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_27),
.B(n_9),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_65),
.Y(n_151)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_66),
.Y(n_156)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_67),
.Y(n_160)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_18),
.B1(n_9),
.B2(n_11),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_35),
.B1(n_50),
.B2(n_31),
.Y(n_110)
);

NAND2x1_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_8),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_73),
.A2(n_35),
.B(n_12),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_23),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_74),
.B(n_78),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_29),
.B(n_8),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_44),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_29),
.B(n_8),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_83),
.B(n_86),
.Y(n_162)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_28),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_84),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_23),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_89),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_31),
.B(n_32),
.C(n_45),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_104),
.B(n_106),
.Y(n_171)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_73),
.A2(n_50),
.B1(n_35),
.B2(n_48),
.Y(n_108)
);

AO22x1_ASAP7_75t_SL g214 ( 
.A1(n_108),
.A2(n_152),
.B1(n_25),
.B2(n_39),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_110),
.A2(n_117),
.B1(n_166),
.B2(n_36),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_47),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_112),
.B(n_127),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_65),
.A2(n_42),
.B1(n_49),
.B2(n_25),
.Y(n_117)
);

BUFx2_ASAP7_75t_R g123 ( 
.A(n_84),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_123),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_47),
.Y(n_127)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_143),
.Y(n_217)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_157),
.Y(n_185)
);

BUFx12_ASAP7_75t_L g147 ( 
.A(n_55),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_55),
.A2(n_31),
.B1(n_48),
.B2(n_49),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_152),
.A2(n_50),
.B1(n_81),
.B2(n_85),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_46),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_172),
.Y(n_183)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_54),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_158),
.B(n_36),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_51),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_56),
.A2(n_41),
.B1(n_32),
.B2(n_45),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_66),
.B(n_46),
.Y(n_172)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_67),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_121),
.A2(n_48),
.B1(n_31),
.B2(n_71),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_178),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_179),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_117),
.A2(n_102),
.B1(n_98),
.B2(n_100),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_180),
.A2(n_196),
.B1(n_229),
.B2(n_230),
.Y(n_275)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_181),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_148),
.A2(n_71),
.B1(n_64),
.B2(n_60),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_184),
.A2(n_210),
.B1(n_216),
.B2(n_221),
.Y(n_262)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_187),
.Y(n_260)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_188),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_149),
.Y(n_189)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_189),
.Y(n_266)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_191),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_108),
.A2(n_75),
.B1(n_77),
.B2(n_88),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_193),
.A2(n_197),
.B1(n_201),
.B2(n_211),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_194),
.Y(n_281)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_114),
.Y(n_195)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_195),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_108),
.A2(n_96),
.B1(n_95),
.B2(n_90),
.Y(n_196)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_198),
.Y(n_276)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_200),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_138),
.B1(n_111),
.B2(n_162),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_202),
.Y(n_269)
);

INVx4_ASAP7_75t_SL g203 ( 
.A(n_125),
.Y(n_203)
);

INVx13_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_204),
.Y(n_270)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_205),
.Y(n_253)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_207),
.Y(n_257)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_208),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_209),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_116),
.A2(n_64),
.B1(n_79),
.B2(n_69),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_171),
.A2(n_93),
.B1(n_61),
.B2(n_59),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_138),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_212),
.B(n_220),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_58),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_213),
.B(n_227),
.C(n_231),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_214),
.A2(n_218),
.B1(n_235),
.B2(n_175),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_133),
.Y(n_215)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_131),
.A2(n_49),
.B1(n_42),
.B2(n_40),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_111),
.A2(n_40),
.B1(n_39),
.B2(n_37),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_120),
.Y(n_219)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_219),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_162),
.B(n_128),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_165),
.A2(n_40),
.B1(n_39),
.B2(n_37),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_124),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_222),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_137),
.B(n_37),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_236),
.Y(n_241)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_134),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_224),
.B(n_233),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_226),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_147),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_109),
.B(n_0),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_153),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_232),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_164),
.A2(n_36),
.B1(n_25),
.B2(n_20),
.Y(n_230)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_118),
.B(n_0),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_129),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_125),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_136),
.B(n_20),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_234),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_139),
.A2(n_20),
.B1(n_19),
.B2(n_26),
.Y(n_235)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_115),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_126),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_238),
.Y(n_247)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_167),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_183),
.C(n_206),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_242),
.B(n_265),
.C(n_283),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_211),
.B(n_119),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_249),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_229),
.A2(n_173),
.B1(n_146),
.B2(n_126),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_251),
.A2(n_255),
.B1(n_264),
.B2(n_268),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_209),
.A2(n_144),
.B(n_132),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_252),
.A2(n_2),
.B(n_6),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_214),
.A2(n_142),
.B1(n_150),
.B2(n_156),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_183),
.B(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_256),
.B(n_278),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_259),
.B(n_249),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_214),
.A2(n_156),
.B1(n_146),
.B2(n_169),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_213),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_223),
.A2(n_115),
.B1(n_19),
.B2(n_24),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_227),
.B(n_0),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_227),
.B(n_0),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_279),
.B(n_287),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_213),
.A2(n_19),
.B1(n_26),
.B2(n_24),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_282),
.A2(n_286),
.B1(n_2),
.B2(n_5),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_209),
.B(n_26),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_224),
.A2(n_185),
.B1(n_238),
.B2(n_188),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_284),
.A2(n_204),
.B1(n_205),
.B2(n_189),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_202),
.A2(n_26),
.B1(n_24),
.B2(n_3),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_217),
.B(n_1),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_244),
.A2(n_222),
.B1(n_187),
.B2(n_177),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_290),
.A2(n_297),
.B1(n_310),
.B2(n_318),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_291),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_192),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_292),
.B(n_293),
.C(n_315),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_182),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_186),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_295),
.B(n_298),
.Y(n_356)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_247),
.Y(n_296)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_296),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_244),
.A2(n_176),
.B1(n_237),
.B2(n_207),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_240),
.B(n_261),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_252),
.Y(n_299)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_299),
.Y(n_350)
);

MAJx3_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_283),
.C(n_289),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_300),
.A2(n_321),
.B(n_327),
.Y(n_369)
);

AO21x2_ASAP7_75t_L g301 ( 
.A1(n_241),
.A2(n_198),
.B(n_200),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_301),
.A2(n_308),
.B1(n_320),
.B2(n_322),
.Y(n_361)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_303),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_288),
.B(n_194),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_258),
.B(n_195),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_305),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_329),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_275),
.A2(n_176),
.B1(n_228),
.B2(n_191),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_274),
.A2(n_276),
.B1(n_262),
.B2(n_251),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_309),
.A2(n_314),
.B(n_266),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_274),
.A2(n_189),
.B(n_236),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_311),
.A2(n_273),
.B(n_269),
.Y(n_360)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_247),
.Y(n_312)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_312),
.Y(n_362)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_239),
.Y(n_313)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_313),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_276),
.A2(n_181),
.B1(n_190),
.B2(n_232),
.Y(n_314)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_242),
.B(n_203),
.C(n_208),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_277),
.B(n_219),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_317),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_259),
.A2(n_179),
.B1(n_199),
.B2(n_26),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_199),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_319),
.B(n_260),
.C(n_245),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_249),
.A2(n_24),
.B1(n_12),
.B2(n_3),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_SL g321 ( 
.A1(n_241),
.A2(n_199),
.B(n_24),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_249),
.A2(n_11),
.B1(n_16),
.B2(n_5),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_1),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_323),
.B(n_325),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_254),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_324),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_278),
.B(n_2),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_268),
.B(n_2),
.Y(n_326)
);

NAND2x1_ASAP7_75t_L g351 ( 
.A(n_326),
.B(n_310),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_248),
.Y(n_327)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_250),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_332),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_284),
.A2(n_279),
.B1(n_253),
.B2(n_257),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_331),
.A2(n_308),
.B1(n_306),
.B2(n_312),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_246),
.B(n_2),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_333),
.B(n_243),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_334),
.A2(n_367),
.B1(n_347),
.B2(n_350),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_302),
.A2(n_286),
.B1(n_272),
.B2(n_250),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_336),
.A2(n_347),
.B1(n_365),
.B2(n_367),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_310),
.A2(n_272),
.B1(n_246),
.B2(n_271),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_338),
.A2(n_363),
.B1(n_366),
.B2(n_301),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_340),
.B(n_343),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_243),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_299),
.A2(n_271),
.B(n_248),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_302),
.A2(n_267),
.B1(n_270),
.B2(n_263),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_351),
.Y(n_402)
);

AND2x6_ASAP7_75t_L g353 ( 
.A(n_300),
.B(n_263),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_353),
.B(n_357),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_293),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_358),
.C(n_319),
.Y(n_375)
);

OAI32xp33_ASAP7_75t_L g357 ( 
.A1(n_296),
.A2(n_270),
.A3(n_260),
.B1(n_245),
.B2(n_269),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_360),
.A2(n_364),
.B(n_368),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_297),
.A2(n_267),
.B1(n_273),
.B2(n_11),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_316),
.B(n_332),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_290),
.A2(n_17),
.B1(n_7),
.B2(n_13),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_301),
.A2(n_6),
.B1(n_7),
.B2(n_14),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_311),
.A2(n_6),
.B(n_14),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g371 ( 
.A(n_300),
.B(n_14),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_322),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_356),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_372),
.B(n_377),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_348),
.A2(n_301),
.B1(n_331),
.B2(n_328),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_373),
.A2(n_390),
.B1(n_404),
.B2(n_341),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_374),
.A2(n_384),
.B(n_399),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_375),
.B(n_380),
.C(n_383),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_356),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_379),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_355),
.B(n_354),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_363),
.Y(n_381)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_381),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_354),
.B(n_292),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_350),
.A2(n_343),
.B(n_364),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_370),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_385),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_342),
.B(n_313),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g407 ( 
.A(n_386),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_358),
.B(n_315),
.C(n_294),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_388),
.B(n_397),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_342),
.B(n_333),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_389),
.B(n_391),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_348),
.A2(n_301),
.B1(n_294),
.B2(n_320),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_335),
.B(n_303),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_395),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_361),
.A2(n_318),
.B1(n_326),
.B2(n_307),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_394),
.A2(n_396),
.B1(n_403),
.B2(n_366),
.Y(n_406)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_370),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_361),
.A2(n_326),
.B1(n_307),
.B2(n_323),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_369),
.B(n_291),
.C(n_325),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_327),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_398),
.B(n_400),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_343),
.A2(n_330),
.B(n_16),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_338),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_359),
.B(n_15),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_401),
.B(n_349),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_365),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_362),
.A2(n_16),
.B1(n_17),
.B2(n_337),
.Y(n_404)
);

OAI22x1_ASAP7_75t_L g405 ( 
.A1(n_353),
.A2(n_337),
.B1(n_334),
.B2(n_369),
.Y(n_405)
);

AOI22x1_ASAP7_75t_L g414 ( 
.A1(n_405),
.A2(n_364),
.B1(n_352),
.B2(n_336),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_406),
.A2(n_393),
.B1(n_378),
.B2(n_381),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_410),
.A2(n_416),
.B1(n_424),
.B2(n_387),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_386),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_412),
.B(n_413),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_392),
.A2(n_374),
.B1(n_394),
.B2(n_396),
.Y(n_413)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_414),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_402),
.A2(n_352),
.B1(n_359),
.B2(n_341),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_398),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_417),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_389),
.B(n_335),
.Y(n_418)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_418),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_391),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_419),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_404),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_421),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_388),
.B(n_380),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_422),
.B(n_420),
.Y(n_455)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_423),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_373),
.A2(n_341),
.B1(n_352),
.B2(n_345),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_357),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_426),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_380),
.B(n_340),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_429),
.B(n_433),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_372),
.B(n_346),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_432),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_375),
.B(n_339),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_377),
.B(n_346),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_434),
.B(n_385),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_390),
.B(n_339),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_435),
.B(n_406),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_383),
.C(n_397),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_436),
.B(n_437),
.C(n_459),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_427),
.B(n_383),
.C(n_384),
.Y(n_437)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_441),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_442),
.A2(n_446),
.B1(n_449),
.B2(n_407),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_405),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_443),
.B(n_444),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_405),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_445),
.B(n_457),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_410),
.A2(n_378),
.B1(n_392),
.B2(n_379),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_448),
.A2(n_425),
.B1(n_409),
.B2(n_426),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_435),
.A2(n_381),
.B1(n_376),
.B2(n_403),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_433),
.B(n_376),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_450),
.B(n_455),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_425),
.A2(n_382),
.B(n_399),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_420),
.B(n_351),
.C(n_382),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_351),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_460),
.B(n_461),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_434),
.B(n_371),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_437),
.C(n_455),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_464),
.B(n_470),
.C(n_472),
.Y(n_493)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_441),
.Y(n_465)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_465),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_451),
.A2(n_424),
.B(n_416),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_466),
.A2(n_457),
.B(n_453),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_418),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_467),
.B(n_349),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_468),
.A2(n_473),
.B1(n_475),
.B2(n_449),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_SL g469 ( 
.A1(n_442),
.A2(n_430),
.B1(n_409),
.B2(n_431),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_469),
.A2(n_479),
.B1(n_454),
.B2(n_459),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_440),
.B(n_413),
.C(n_414),
.Y(n_470)
);

OA21x2_ASAP7_75t_SL g471 ( 
.A1(n_438),
.A2(n_408),
.B(n_415),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_471),
.B(n_481),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_436),
.B(n_414),
.C(n_417),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_448),
.A2(n_415),
.B1(n_408),
.B2(n_430),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_452),
.A2(n_421),
.B1(n_419),
.B2(n_412),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_441),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_477),
.B(n_478),
.Y(n_483)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_451),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_450),
.B(n_411),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_481),
.B(n_445),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_486),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_462),
.B(n_439),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_487),
.A2(n_488),
.B(n_466),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_472),
.A2(n_453),
.B(n_458),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_462),
.B(n_456),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_489),
.B(n_475),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_490),
.A2(n_482),
.B1(n_477),
.B2(n_465),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_491),
.A2(n_468),
.B1(n_470),
.B2(n_478),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_473),
.A2(n_446),
.B1(n_443),
.B2(n_444),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_492),
.A2(n_474),
.B1(n_360),
.B2(n_428),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_496),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_460),
.C(n_461),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_498),
.C(n_480),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_479),
.B(n_423),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_463),
.B(n_411),
.C(n_428),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_499),
.B(n_507),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_500),
.B(n_509),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_501),
.A2(n_490),
.B1(n_492),
.B2(n_487),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_498),
.B(n_464),
.C(n_482),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_502),
.B(n_505),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_503),
.B(n_508),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_493),
.B(n_495),
.C(n_491),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_476),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_493),
.A2(n_471),
.B(n_480),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_488),
.B(n_476),
.C(n_474),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_510),
.B(n_511),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_506),
.B(n_484),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_515),
.B(n_521),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_517),
.Y(n_528)
);

BUFx24_ASAP7_75t_SL g518 ( 
.A(n_504),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_518),
.B(n_520),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_484),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_502),
.B(n_486),
.Y(n_521)
);

AOI21x1_ASAP7_75t_SL g522 ( 
.A1(n_514),
.A2(n_489),
.B(n_516),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_522),
.A2(n_523),
.B(n_524),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_508),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_519),
.A2(n_505),
.B(n_500),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_519),
.A2(n_483),
.B(n_510),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_527),
.A2(n_499),
.B1(n_501),
.B2(n_497),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_529),
.A2(n_530),
.B(n_531),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_526),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_513),
.Y(n_531)
);

A2O1A1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_532),
.A2(n_528),
.B(n_523),
.C(n_483),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_513),
.B(n_507),
.Y(n_535)
);

O2A1O1Ixp33_ASAP7_75t_SL g537 ( 
.A1(n_535),
.A2(n_536),
.B(n_503),
.C(n_395),
.Y(n_537)
);

BUFx24_ASAP7_75t_SL g536 ( 
.A(n_533),
.Y(n_536)
);

AO21x2_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_368),
.B(n_401),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_538),
.B(n_344),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_344),
.Y(n_540)
);


endmodule