module fake_jpeg_16649_n_348 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_45),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_18),
.B(n_8),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_21),
.Y(n_57)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_38),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_37),
.B1(n_24),
.B2(n_38),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_53),
.A2(n_31),
.B1(n_26),
.B2(n_30),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_24),
.B1(n_37),
.B2(n_25),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_56),
.B1(n_19),
.B2(n_18),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_37),
.B1(n_25),
.B2(n_24),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_57),
.B(n_29),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_62),
.B(n_45),
.Y(n_108)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_36),
.C(n_20),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_67),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_20),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_35),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_72),
.Y(n_112)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_34),
.B(n_48),
.C(n_20),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_73),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_51),
.A2(n_24),
.B1(n_44),
.B2(n_38),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_74),
.A2(n_78),
.B1(n_81),
.B2(n_85),
.Y(n_116)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_47),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_86),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_25),
.B1(n_18),
.B2(n_21),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_19),
.B(n_44),
.C(n_20),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_80),
.A2(n_107),
.B(n_17),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_38),
.B1(n_43),
.B2(n_42),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_82),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_29),
.B1(n_43),
.B2(n_42),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_105),
.B1(n_59),
.B2(n_81),
.Y(n_111)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_61),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_21),
.B1(n_22),
.B2(n_32),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_47),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_90),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_63),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_92),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_19),
.C(n_31),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_108),
.C(n_17),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_40),
.B1(n_32),
.B2(n_22),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_91),
.B1(n_98),
.B2(n_101),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_22),
.B1(n_32),
.B2(n_29),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_95),
.Y(n_127)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_102),
.Y(n_136)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_33),
.B1(n_26),
.B2(n_30),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_104),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_53),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_59),
.A2(n_35),
.B1(n_33),
.B2(n_40),
.Y(n_105)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_109),
.B(n_110),
.Y(n_114)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_115),
.B1(n_94),
.B2(n_84),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_106),
.A2(n_59),
.B1(n_65),
.B2(n_67),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_117),
.A2(n_132),
.B1(n_124),
.B2(n_125),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_107),
.B1(n_71),
.B2(n_74),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_128),
.B(n_133),
.Y(n_144)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_36),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_70),
.B(n_61),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_131),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_61),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_45),
.C(n_39),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_135),
.C(n_140),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_0),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_80),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_27),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_98),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_72),
.B(n_62),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_143),
.B(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_147),
.B(n_152),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_112),
.A2(n_75),
.B(n_23),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_148),
.A2(n_156),
.B(n_167),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_149),
.A2(n_169),
.B1(n_170),
.B2(n_137),
.Y(n_178)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_127),
.B(n_75),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_99),
.B1(n_103),
.B2(n_109),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_161),
.B1(n_143),
.B2(n_162),
.Y(n_180)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_155),
.Y(n_189)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_76),
.B(n_39),
.C(n_110),
.D(n_100),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_126),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_159),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_122),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_97),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_162),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_100),
.B1(n_11),
.B2(n_16),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_17),
.Y(n_162)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_163),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_112),
.B(n_17),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_118),
.Y(n_172)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_166),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_0),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_168),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_116),
.A2(n_102),
.B1(n_79),
.B2(n_23),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_158),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_148),
.A2(n_140),
.B(n_131),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_173),
.A2(n_199),
.B(n_201),
.Y(n_231)
);

OAI22x1_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_116),
.B1(n_140),
.B2(n_118),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_175),
.A2(n_177),
.B1(n_178),
.B2(n_147),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_165),
.A2(n_119),
.B1(n_140),
.B2(n_118),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_180),
.A2(n_202),
.B1(n_169),
.B2(n_150),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_117),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_187),
.C(n_190),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_155),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_186),
.B(n_192),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_119),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_136),
.C(n_139),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_145),
.B(n_133),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_133),
.Y(n_196)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_144),
.B(n_160),
.C(n_151),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_187),
.C(n_190),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_167),
.A2(n_111),
.B1(n_134),
.B2(n_136),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_142),
.B(n_127),
.Y(n_200)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_144),
.A2(n_120),
.B(n_134),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_153),
.A2(n_130),
.B1(n_138),
.B2(n_122),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_201),
.A2(n_161),
.B(n_167),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_203),
.A2(n_4),
.B(n_5),
.Y(n_259)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_154),
.Y(n_205)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_205),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_120),
.Y(n_206)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_208),
.A2(n_202),
.B1(n_196),
.B2(n_191),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_176),
.B(n_198),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_221),
.Y(n_251)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_226),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_163),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_228),
.C(n_234),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_218),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_219),
.B1(n_224),
.B2(n_232),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_166),
.Y(n_216)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_137),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_217),
.Y(n_243)
);

AO22x1_ASAP7_75t_L g218 ( 
.A1(n_175),
.A2(n_164),
.B1(n_82),
.B2(n_23),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_177),
.A2(n_200),
.B1(n_182),
.B2(n_193),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_179),
.B(n_9),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_220),
.B(n_222),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_173),
.B(n_16),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_180),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_225),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_172),
.B(n_1),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_182),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_230),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_3),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_194),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_233),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_184),
.B(n_10),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_215),
.A2(n_213),
.B1(n_225),
.B2(n_207),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_235),
.A2(n_252),
.B1(n_230),
.B2(n_210),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_214),
.B1(n_224),
.B2(n_216),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_176),
.C(n_184),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_244),
.C(n_249),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_199),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_192),
.C(n_186),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_185),
.C(n_189),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_255),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_207),
.A2(n_185),
.B1(n_181),
.B2(n_5),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_209),
.B(n_181),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_212),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_218),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_3),
.C(n_4),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_226),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_259),
.A2(n_221),
.B(n_203),
.Y(n_263)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_257),
.Y(n_260)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_261),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_223),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_265),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_263),
.A2(n_251),
.B(n_259),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_231),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_269),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_223),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_253),
.A2(n_231),
.B(n_245),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_266),
.A2(n_279),
.B(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_273),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_234),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_250),
.C(n_249),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_253),
.B1(n_241),
.B2(n_258),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_276),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_247),
.B(n_232),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_238),
.B(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_236),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_240),
.A2(n_218),
.B1(n_5),
.B2(n_6),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_278),
.A2(n_12),
.B1(n_16),
.B2(n_14),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_248),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_235),
.Y(n_280)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_286),
.C(n_292),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_274),
.C(n_264),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_236),
.Y(n_290)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_290),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_291),
.B(n_272),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_239),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_239),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_299),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_294),
.A2(n_263),
.B(n_260),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_270),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_242),
.C(n_251),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_10),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_11),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_300),
.A2(n_308),
.B(n_291),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_302),
.A2(n_305),
.B1(n_311),
.B2(n_299),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_297),
.B(n_278),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_307),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_261),
.B(n_267),
.Y(n_305)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_11),
.Y(n_307)
);

MAJx2_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_10),
.C(n_12),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_296),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_284),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_313),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_287),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_307),
.Y(n_324)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_316),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_295),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_319),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_281),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_285),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_320),
.A2(n_321),
.B1(n_306),
.B2(n_289),
.Y(n_329)
);

INVx11_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_322),
.A2(n_308),
.B1(n_303),
.B2(n_288),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_325),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_323),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_331),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_318),
.A2(n_300),
.B(n_303),
.Y(n_328)
);

OAI31xp33_ASAP7_75t_SL g336 ( 
.A1(n_328),
.A2(n_333),
.A3(n_334),
.B(n_321),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_324),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_315),
.A2(n_293),
.B(n_292),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_315),
.A2(n_309),
.B(n_286),
.Y(n_334)
);

AOI21x1_ASAP7_75t_L g343 ( 
.A1(n_336),
.A2(n_298),
.B(n_12),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_320),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_337),
.B(n_338),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_327),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_339),
.B(n_340),
.C(n_332),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_309),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_341),
.A2(n_343),
.B(n_337),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_342),
.B1(n_335),
.B2(n_14),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_345),
.A2(n_13),
.B(n_14),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_13),
.Y(n_347)
);

FAx1_ASAP7_75t_SL g348 ( 
.A(n_347),
.B(n_6),
.CI(n_345),
.CON(n_348),
.SN(n_348)
);


endmodule