module fake_jpeg_15507_n_297 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_107;
wire n_39;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_9),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_44),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_16),
.B(n_0),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_53),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_54),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_15),
.B(n_1),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_1),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_1),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_58),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_19),
.B(n_2),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_63),
.Y(n_89)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_18),
.B(n_2),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_5),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_70),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_21),
.B(n_5),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_21),
.B(n_41),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_41),
.Y(n_98)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_37),
.B1(n_26),
.B2(n_33),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_86),
.A2(n_101),
.B1(n_120),
.B2(n_10),
.Y(n_158)
);

AND2x4_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_32),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_87),
.A2(n_27),
.B(n_32),
.C(n_25),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_40),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_100),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_33),
.B1(n_26),
.B2(n_32),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_29),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_105),
.B(n_106),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_29),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_51),
.B(n_24),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_107),
.B(n_110),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_55),
.B(n_40),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_109),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_28),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_39),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_48),
.B(n_28),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_24),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_60),
.A2(n_26),
.B1(n_38),
.B2(n_30),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_116),
.B1(n_34),
.B2(n_32),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_50),
.A2(n_39),
.B1(n_38),
.B2(n_30),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_56),
.B(n_20),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_89),
.Y(n_141)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_66),
.A2(n_32),
.B1(n_25),
.B2(n_23),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_20),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_111),
.Y(n_165)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_34),
.C(n_25),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_124),
.B(n_139),
.C(n_96),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_87),
.A2(n_27),
.B1(n_76),
.B2(n_73),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_125),
.A2(n_158),
.B1(n_124),
.B2(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_94),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_132),
.B(n_136),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_86),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_95),
.A2(n_34),
.B1(n_23),
.B2(n_32),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_134),
.A2(n_79),
.B(n_90),
.Y(n_181)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_123),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_141),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_138),
.A2(n_156),
.B1(n_145),
.B2(n_139),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_81),
.B(n_72),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_143),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_82),
.B(n_5),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_102),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_85),
.B(n_6),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g147 ( 
.A(n_96),
.Y(n_147)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_7),
.Y(n_150)
);

BUFx24_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_94),
.B(n_13),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_153),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_13),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_8),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_161),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_90),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_159),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_104),
.A2(n_119),
.B1(n_100),
.B2(n_88),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_13),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_95),
.B(n_103),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_162),
.B(n_118),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_165),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_163),
.A2(n_84),
.B1(n_97),
.B2(n_83),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_166),
.A2(n_189),
.B1(n_164),
.B2(n_132),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_127),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_172),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_181),
.B(n_188),
.Y(n_198)
);

AOI32xp33_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_88),
.A3(n_83),
.B1(n_118),
.B2(n_79),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_174),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_196),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_79),
.B(n_90),
.C(n_133),
.Y(n_188)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_160),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_160),
.C(n_149),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_126),
.B(n_130),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_136),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_139),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_134),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_200),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_142),
.Y(n_201)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g202 ( 
.A(n_167),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_202),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_140),
.C(n_144),
.Y(n_204)
);

OAI211xp5_ASAP7_75t_L g230 ( 
.A1(n_204),
.A2(n_185),
.B(n_173),
.C(n_178),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_146),
.Y(n_206)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_158),
.Y(n_207)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_170),
.A2(n_148),
.B1(n_162),
.B2(n_135),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_220),
.B1(n_222),
.B2(n_183),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_175),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_210),
.A2(n_174),
.B(n_169),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_175),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_213),
.A2(n_217),
.B1(n_219),
.B2(n_221),
.Y(n_235)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_157),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_172),
.A2(n_164),
.B1(n_147),
.B2(n_148),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_170),
.A2(n_189),
.B1(n_186),
.B2(n_193),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_171),
.B1(n_196),
.B2(n_184),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_SL g254 ( 
.A1(n_224),
.A2(n_227),
.B(n_242),
.C(n_180),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_222),
.A2(n_181),
.B1(n_188),
.B2(n_182),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_226),
.B(n_231),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_203),
.A2(n_209),
.B1(n_200),
.B2(n_220),
.Y(n_227)
);

AOI221xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_214),
.B1(n_203),
.B2(n_208),
.C(n_199),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_206),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_198),
.A2(n_166),
.B1(n_176),
.B2(n_177),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_185),
.B(n_176),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_234),
.A2(n_228),
.B(n_232),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_177),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_203),
.C(n_210),
.Y(n_246)
);

OA21x2_ASAP7_75t_L g242 ( 
.A1(n_201),
.A2(n_180),
.B(n_190),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_257),
.B(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_247),
.C(n_252),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_205),
.C(n_219),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_232),
.A2(n_221),
.B(n_215),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_253),
.B(n_231),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_236),
.Y(n_249)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_218),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_250),
.B(n_255),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_235),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_256),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_205),
.C(n_211),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_254),
.A2(n_225),
.B(n_234),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_218),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_147),
.Y(n_257)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_259),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_260),
.B(n_224),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_227),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_265),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_239),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_241),
.C(n_233),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_254),
.C(n_155),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_249),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_271),
.B(n_273),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_258),
.C(n_245),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_275),
.Y(n_281)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_261),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_276),
.Y(n_279)
);

AOI322xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_248),
.A3(n_254),
.B1(n_226),
.B2(n_223),
.C1(n_178),
.C2(n_168),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_278),
.B(n_266),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_285),
.Y(n_287)
);

OAI31xp33_ASAP7_75t_L g283 ( 
.A1(n_278),
.A2(n_259),
.A3(n_269),
.B(n_262),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_283),
.A2(n_151),
.B(n_168),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_263),
.C(n_274),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_264),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_279),
.C(n_151),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_265),
.B(n_151),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_288),
.A2(n_289),
.B(n_290),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_287),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_292),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_291),
.C(n_129),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_294),
.Y(n_297)
);


endmodule