module fake_jpeg_7841_n_59 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_3),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

AO21x1_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_6),
.B(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_35),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

A2O1A1O1Ixp25_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_21),
.B(n_24),
.C(n_14),
.D(n_20),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_41),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_24),
.B1(n_25),
.B2(n_21),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_39),
.B1(n_40),
.B2(n_10),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_13),
.B1(n_17),
.B2(n_7),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_5),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_44),
.B(n_45),
.Y(n_46)
);

FAx1_ASAP7_75t_SL g45 ( 
.A(n_30),
.B(n_6),
.CI(n_19),
.CON(n_45),
.SN(n_45)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_50),
.C(n_51),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_43),
.B(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_11),
.C(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_53),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_48),
.B1(n_46),
.B2(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_49),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_54),
.B1(n_36),
.B2(n_44),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_52),
.Y(n_59)
);


endmodule