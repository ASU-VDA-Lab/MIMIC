module real_aes_8963_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_283;
wire n_252;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g431 ( .A(n_0), .Y(n_431) );
INVx1_ASAP7_75t_L g530 ( .A(n_1), .Y(n_530) );
INVx1_ASAP7_75t_L g183 ( .A(n_2), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_3), .A2(n_39), .B1(n_145), .B2(n_472), .Y(n_489) );
AOI21xp33_ASAP7_75t_L g124 ( .A1(n_4), .A2(n_125), .B(n_132), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_5), .B(n_118), .Y(n_521) );
AND2x6_ASAP7_75t_L g130 ( .A(n_6), .B(n_131), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_7), .A2(n_224), .B(n_225), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_8), .B(n_41), .Y(n_432) );
INVx1_ASAP7_75t_L g142 ( .A(n_9), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_10), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g123 ( .A(n_11), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_12), .B(n_155), .Y(n_467) );
INVx1_ASAP7_75t_L g230 ( .A(n_13), .Y(n_230) );
INVx1_ASAP7_75t_L g525 ( .A(n_14), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_15), .B(n_119), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_16), .A2(n_741), .B1(n_742), .B2(n_745), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_16), .Y(n_745) );
AO32x2_ASAP7_75t_L g487 ( .A1(n_17), .A2(n_118), .A3(n_152), .B1(n_488), .B2(n_492), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_18), .B(n_145), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_19), .B(n_171), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_20), .B(n_119), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_21), .A2(n_52), .B1(n_145), .B2(n_472), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_22), .B(n_125), .Y(n_195) );
AOI22xp33_ASAP7_75t_SL g500 ( .A1(n_23), .A2(n_78), .B1(n_145), .B2(n_155), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_24), .B(n_145), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_25), .B(n_116), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_26), .A2(n_228), .B(n_229), .C(n_231), .Y(n_227) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_27), .A2(n_76), .B1(n_743), .B2(n_744), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_27), .Y(n_744) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_28), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_29), .B(n_148), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_30), .B(n_140), .Y(n_185) );
INVx1_ASAP7_75t_L g161 ( .A(n_31), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_32), .B(n_148), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_33), .B(n_427), .Y(n_436) );
INVx2_ASAP7_75t_L g128 ( .A(n_34), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_35), .B(n_145), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_36), .B(n_148), .Y(n_473) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_37), .A2(n_64), .B1(n_107), .B2(n_108), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_37), .Y(n_107) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_38), .A2(n_130), .B(n_135), .C(n_197), .Y(n_196) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_40), .A2(n_447), .B1(n_739), .B2(n_740), .C1(n_746), .C2(n_750), .Y(n_446) );
INVx1_ASAP7_75t_L g159 ( .A(n_42), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_43), .B(n_140), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_44), .B(n_145), .Y(n_515) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_45), .A2(n_103), .B1(n_437), .B2(n_445), .C1(n_753), .C2(n_758), .Y(n_102) );
OAI321xp33_ASAP7_75t_L g103 ( .A1(n_45), .A2(n_104), .A3(n_427), .B1(n_433), .B2(n_434), .C(n_436), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g433 ( .A(n_45), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_46), .A2(n_88), .B1(n_202), .B2(n_472), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_47), .B(n_145), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_48), .B(n_145), .Y(n_526) );
CKINVDCx16_ASAP7_75t_R g162 ( .A(n_49), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_50), .B(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_51), .B(n_125), .Y(n_218) );
AOI22xp33_ASAP7_75t_SL g510 ( .A1(n_53), .A2(n_62), .B1(n_145), .B2(n_155), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_54), .A2(n_135), .B1(n_155), .B2(n_157), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_55), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_56), .B(n_145), .Y(n_466) );
CKINVDCx16_ASAP7_75t_R g180 ( .A(n_57), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_58), .B(n_145), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g138 ( .A1(n_59), .A2(n_139), .B(n_141), .C(n_144), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_60), .Y(n_248) );
INVx1_ASAP7_75t_L g133 ( .A(n_61), .Y(n_133) );
INVx1_ASAP7_75t_L g131 ( .A(n_63), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_64), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_65), .B(n_145), .Y(n_531) );
INVx1_ASAP7_75t_L g122 ( .A(n_66), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_67), .Y(n_441) );
AO32x2_ASAP7_75t_L g497 ( .A1(n_68), .A2(n_118), .A3(n_210), .B1(n_492), .B2(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g542 ( .A(n_69), .Y(n_542) );
INVx1_ASAP7_75t_L g480 ( .A(n_70), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_SL g170 ( .A1(n_71), .A2(n_144), .B(n_171), .C(n_172), .Y(n_170) );
INVxp67_ASAP7_75t_L g173 ( .A(n_72), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_73), .B(n_155), .Y(n_481) );
INVx1_ASAP7_75t_L g444 ( .A(n_74), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_75), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_76), .Y(n_743) );
INVx1_ASAP7_75t_L g241 ( .A(n_77), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_79), .A2(n_130), .B(n_135), .C(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_80), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_81), .B(n_155), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_82), .B(n_184), .Y(n_198) );
INVx2_ASAP7_75t_L g120 ( .A(n_83), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_84), .B(n_171), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_85), .B(n_155), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_86), .A2(n_130), .B(n_135), .C(n_182), .Y(n_181) );
OR2x2_ASAP7_75t_L g428 ( .A(n_87), .B(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g452 ( .A(n_87), .B(n_430), .Y(n_452) );
INVx2_ASAP7_75t_L g455 ( .A(n_87), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_89), .A2(n_101), .B1(n_155), .B2(n_156), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_90), .B(n_148), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_91), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_92), .A2(n_130), .B(n_135), .C(n_213), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_93), .Y(n_220) );
INVx1_ASAP7_75t_L g169 ( .A(n_94), .Y(n_169) );
CKINVDCx16_ASAP7_75t_R g226 ( .A(n_95), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_96), .B(n_184), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_97), .B(n_155), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_98), .B(n_118), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_99), .A2(n_125), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_100), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_104), .B(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_106), .B1(n_109), .B2(n_426), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_109), .A2(n_457), .B1(n_748), .B2(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g426 ( .A(n_110), .Y(n_426) );
AND3x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_348), .C(n_393), .Y(n_110) );
NOR4xp25_ASAP7_75t_L g111 ( .A(n_112), .B(n_271), .C(n_312), .D(n_329), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_175), .B(n_191), .C(n_233), .Y(n_112) );
OR2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_149), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_114), .B(n_176), .Y(n_175) );
NOR4xp25_ASAP7_75t_L g295 ( .A(n_114), .B(n_289), .C(n_296), .D(n_302), .Y(n_295) );
AND2x2_ASAP7_75t_L g368 ( .A(n_114), .B(n_257), .Y(n_368) );
AND2x2_ASAP7_75t_L g387 ( .A(n_114), .B(n_333), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_114), .B(n_382), .Y(n_396) );
AND2x2_ASAP7_75t_L g409 ( .A(n_114), .B(n_190), .Y(n_409) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g254 ( .A(n_115), .Y(n_254) );
AND2x2_ASAP7_75t_L g261 ( .A(n_115), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g311 ( .A(n_115), .B(n_150), .Y(n_311) );
AND2x2_ASAP7_75t_SL g322 ( .A(n_115), .B(n_257), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_115), .B(n_150), .Y(n_326) );
AND2x2_ASAP7_75t_L g335 ( .A(n_115), .B(n_260), .Y(n_335) );
BUFx2_ASAP7_75t_L g358 ( .A(n_115), .Y(n_358) );
AND2x2_ASAP7_75t_L g362 ( .A(n_115), .B(n_166), .Y(n_362) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_124), .B(n_147), .Y(n_115) );
INVx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_SL g204 ( .A(n_117), .B(n_205), .Y(n_204) );
NAND3xp33_ASAP7_75t_L g507 ( .A(n_117), .B(n_492), .C(n_508), .Y(n_507) );
AO21x1_ASAP7_75t_L g545 ( .A1(n_117), .A2(n_508), .B(n_546), .Y(n_545) );
INVx4_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_118), .A2(n_167), .B(n_174), .Y(n_166) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_118), .A2(n_513), .B(n_521), .Y(n_512) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g152 ( .A(n_119), .Y(n_152) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
AND2x2_ASAP7_75t_SL g148 ( .A(n_120), .B(n_121), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
BUFx2_ASAP7_75t_L g224 ( .A(n_125), .Y(n_224) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_130), .Y(n_125) );
NAND2x1p5_ASAP7_75t_L g163 ( .A(n_126), .B(n_130), .Y(n_163) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
INVx1_ASAP7_75t_L g520 ( .A(n_127), .Y(n_520) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g136 ( .A(n_128), .Y(n_136) );
INVx1_ASAP7_75t_L g156 ( .A(n_128), .Y(n_156) );
INVx1_ASAP7_75t_L g137 ( .A(n_129), .Y(n_137) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_129), .Y(n_140) );
INVx3_ASAP7_75t_L g143 ( .A(n_129), .Y(n_143) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_129), .Y(n_158) );
INVx1_ASAP7_75t_L g171 ( .A(n_129), .Y(n_171) );
INVx4_ASAP7_75t_SL g146 ( .A(n_130), .Y(n_146) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_130), .A2(n_465), .B(n_469), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_130), .A2(n_479), .B(n_482), .Y(n_478) );
BUFx3_ASAP7_75t_L g492 ( .A(n_130), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_130), .A2(n_514), .B(n_517), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_130), .A2(n_524), .B(n_528), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_134), .B(n_138), .C(n_146), .Y(n_132) );
O2A1O1Ixp33_ASAP7_75t_L g168 ( .A1(n_134), .A2(n_146), .B(n_169), .C(n_170), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_134), .A2(n_146), .B(n_226), .C(n_227), .Y(n_225) );
INVx5_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_136), .Y(n_145) );
BUFx3_ASAP7_75t_L g202 ( .A(n_136), .Y(n_202) );
INVx1_ASAP7_75t_L g472 ( .A(n_136), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_139), .A2(n_470), .B(n_471), .Y(n_469) );
O2A1O1Ixp5_ASAP7_75t_L g541 ( .A1(n_139), .A2(n_529), .B(n_542), .C(n_543), .Y(n_541) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx4_ASAP7_75t_L g216 ( .A(n_140), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_140), .A2(n_489), .B1(n_490), .B2(n_491), .Y(n_488) );
OAI22xp5_ASAP7_75t_SL g498 ( .A1(n_140), .A2(n_143), .B1(n_499), .B2(n_500), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_140), .A2(n_490), .B1(n_509), .B2(n_510), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_143), .B(n_173), .Y(n_172) );
INVx5_ASAP7_75t_L g184 ( .A(n_143), .Y(n_184) );
O2A1O1Ixp5_ASAP7_75t_SL g479 ( .A1(n_144), .A2(n_184), .B(n_480), .C(n_481), .Y(n_479) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
HB1xp67_ASAP7_75t_L g217 ( .A(n_145), .Y(n_217) );
OAI22xp33_ASAP7_75t_L g153 ( .A1(n_146), .A2(n_154), .B1(n_162), .B2(n_163), .Y(n_153) );
INVx1_ASAP7_75t_L g189 ( .A(n_148), .Y(n_189) );
INVx2_ASAP7_75t_L g210 ( .A(n_148), .Y(n_210) );
OA21x2_ASAP7_75t_L g222 ( .A1(n_148), .A2(n_223), .B(n_232), .Y(n_222) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_148), .A2(n_464), .B(n_473), .Y(n_463) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_148), .A2(n_478), .B(n_485), .Y(n_477) );
OR2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_166), .Y(n_149) );
AND2x2_ASAP7_75t_L g190 ( .A(n_150), .B(n_166), .Y(n_190) );
BUFx2_ASAP7_75t_L g264 ( .A(n_150), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_150), .A2(n_297), .B1(n_299), .B2(n_300), .Y(n_296) );
OR2x2_ASAP7_75t_L g318 ( .A(n_150), .B(n_178), .Y(n_318) );
AND2x2_ASAP7_75t_L g382 ( .A(n_150), .B(n_260), .Y(n_382) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g250 ( .A(n_151), .B(n_178), .Y(n_250) );
AND2x2_ASAP7_75t_L g257 ( .A(n_151), .B(n_166), .Y(n_257) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_151), .Y(n_299) );
OR2x2_ASAP7_75t_L g334 ( .A(n_151), .B(n_177), .Y(n_334) );
AO21x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_164), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_152), .B(n_165), .Y(n_164) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_152), .A2(n_179), .B(n_187), .Y(n_178) );
INVx2_ASAP7_75t_L g203 ( .A(n_152), .Y(n_203) );
INVx2_ASAP7_75t_L g186 ( .A(n_155), .Y(n_186) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OAI22xp5_ASAP7_75t_SL g157 ( .A1(n_158), .A2(n_159), .B1(n_160), .B2(n_161), .Y(n_157) );
INVx2_ASAP7_75t_L g160 ( .A(n_158), .Y(n_160) );
INVx4_ASAP7_75t_L g228 ( .A(n_158), .Y(n_228) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_163), .A2(n_180), .B(n_181), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_163), .A2(n_241), .B(n_242), .Y(n_240) );
INVx1_ASAP7_75t_L g253 ( .A(n_166), .Y(n_253) );
INVx3_ASAP7_75t_L g262 ( .A(n_166), .Y(n_262) );
BUFx2_ASAP7_75t_L g286 ( .A(n_166), .Y(n_286) );
AND2x2_ASAP7_75t_L g319 ( .A(n_166), .B(n_254), .Y(n_319) );
INVx1_ASAP7_75t_L g468 ( .A(n_171), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_175), .A2(n_405), .B1(n_406), .B2(n_407), .Y(n_404) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_190), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_177), .B(n_262), .Y(n_266) );
INVx1_ASAP7_75t_L g294 ( .A(n_177), .Y(n_294) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx3_ASAP7_75t_L g260 ( .A(n_178), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_185), .C(n_186), .Y(n_182) );
INVx2_ASAP7_75t_L g490 ( .A(n_184), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_184), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_184), .A2(n_539), .B(n_540), .Y(n_538) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_186), .A2(n_525), .B(n_526), .C(n_527), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_189), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_189), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g272 ( .A(n_190), .Y(n_272) );
NAND2x1_ASAP7_75t_SL g191 ( .A(n_192), .B(n_206), .Y(n_191) );
AND2x2_ASAP7_75t_L g270 ( .A(n_192), .B(n_221), .Y(n_270) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_192), .Y(n_344) );
AND2x2_ASAP7_75t_L g371 ( .A(n_192), .B(n_291), .Y(n_371) );
AND2x2_ASAP7_75t_L g379 ( .A(n_192), .B(n_341), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_192), .B(n_236), .Y(n_406) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g237 ( .A(n_193), .B(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g255 ( .A(n_193), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g276 ( .A(n_193), .Y(n_276) );
INVx1_ASAP7_75t_L g282 ( .A(n_193), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_193), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g315 ( .A(n_193), .B(n_239), .Y(n_315) );
OR2x2_ASAP7_75t_L g353 ( .A(n_193), .B(n_308), .Y(n_353) );
AOI32xp33_ASAP7_75t_L g365 ( .A1(n_193), .A2(n_366), .A3(n_369), .B1(n_370), .B2(n_371), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_193), .B(n_341), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_193), .B(n_301), .Y(n_416) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_204), .Y(n_193) );
AOI21xp5_ASAP7_75t_SL g194 ( .A1(n_195), .A2(n_196), .B(n_203), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_200), .A2(n_244), .B(n_245), .Y(n_243) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g231 ( .A(n_202), .Y(n_231) );
INVx1_ASAP7_75t_L g246 ( .A(n_203), .Y(n_246) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_203), .A2(n_523), .B(n_532), .Y(n_522) );
OA21x2_ASAP7_75t_L g536 ( .A1(n_203), .A2(n_537), .B(n_544), .Y(n_536) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
OR2x2_ASAP7_75t_L g327 ( .A(n_207), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_221), .Y(n_207) );
INVx1_ASAP7_75t_L g289 ( .A(n_208), .Y(n_289) );
AND2x2_ASAP7_75t_L g291 ( .A(n_208), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_208), .B(n_238), .Y(n_308) );
AND2x2_ASAP7_75t_L g341 ( .A(n_208), .B(n_317), .Y(n_341) );
AND2x2_ASAP7_75t_L g378 ( .A(n_208), .B(n_239), .Y(n_378) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g236 ( .A(n_209), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_209), .B(n_238), .Y(n_268) );
AND2x2_ASAP7_75t_L g275 ( .A(n_209), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g316 ( .A(n_209), .B(n_317), .Y(n_316) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_219), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_218), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_217), .Y(n_213) );
INVx2_ASAP7_75t_L g292 ( .A(n_221), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_221), .B(n_238), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_221), .B(n_283), .Y(n_364) );
INVx1_ASAP7_75t_L g386 ( .A(n_221), .Y(n_386) );
INVx1_ASAP7_75t_L g403 ( .A(n_221), .Y(n_403) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g256 ( .A(n_222), .B(n_238), .Y(n_256) );
AND2x2_ASAP7_75t_L g278 ( .A(n_222), .B(n_239), .Y(n_278) );
INVx1_ASAP7_75t_L g317 ( .A(n_222), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_228), .B(n_230), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_228), .A2(n_483), .B(n_484), .Y(n_482) );
INVx1_ASAP7_75t_L g527 ( .A(n_228), .Y(n_527) );
AOI221x1_ASAP7_75t_SL g233 ( .A1(n_234), .A2(n_249), .B1(n_255), .B2(n_257), .C(n_258), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_234), .A2(n_322), .B1(n_389), .B2(n_390), .Y(n_388) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
AND2x2_ASAP7_75t_L g280 ( .A(n_235), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g375 ( .A(n_235), .B(n_255), .Y(n_375) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g331 ( .A(n_236), .B(n_256), .Y(n_331) );
INVx1_ASAP7_75t_L g343 ( .A(n_237), .Y(n_343) );
AND2x2_ASAP7_75t_L g354 ( .A(n_237), .B(n_341), .Y(n_354) );
AND2x2_ASAP7_75t_L g421 ( .A(n_237), .B(n_316), .Y(n_421) );
INVx2_ASAP7_75t_L g283 ( .A(n_238), .Y(n_283) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_246), .B(n_247), .Y(n_239) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_250), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g373 ( .A(n_250), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_251), .B(n_334), .Y(n_337) );
INVx3_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_252), .A2(n_373), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NOR2xp33_ASAP7_75t_SL g395 ( .A(n_255), .B(n_281), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_256), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g347 ( .A(n_256), .B(n_275), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_256), .B(n_282), .Y(n_424) );
AND2x2_ASAP7_75t_L g293 ( .A(n_257), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g360 ( .A(n_257), .Y(n_360) );
AOI21xp33_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_263), .B(n_267), .Y(n_258) );
NAND2x1_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_260), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g309 ( .A(n_260), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_SL g321 ( .A(n_260), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_260), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g345 ( .A(n_261), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_261), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_261), .B(n_264), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
AOI211xp5_ASAP7_75t_L g332 ( .A1(n_264), .A2(n_303), .B(n_333), .C(n_335), .Y(n_332) );
AOI221xp5_ASAP7_75t_L g350 ( .A1(n_264), .A2(n_351), .B1(n_354), .B2(n_355), .C(n_359), .Y(n_350) );
AND2x2_ASAP7_75t_L g346 ( .A(n_265), .B(n_299), .Y(n_346) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g306 ( .A(n_270), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g377 ( .A(n_270), .B(n_378), .Y(n_377) );
OAI211xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_273), .B(n_279), .C(n_304), .Y(n_271) );
NAND3xp33_ASAP7_75t_SL g390 ( .A(n_272), .B(n_391), .C(n_392), .Y(n_390) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_277), .Y(n_273) );
OR2x2_ASAP7_75t_L g363 ( .A(n_274), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_284), .B1(n_287), .B2(n_293), .C(n_295), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_281), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_281), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g303 ( .A(n_286), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_286), .A2(n_343), .B1(n_344), .B2(n_345), .Y(n_342) );
OR2x2_ASAP7_75t_L g423 ( .A(n_286), .B(n_334), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVxp67_ASAP7_75t_L g397 ( .A(n_289), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_291), .B(n_412), .Y(n_411) );
INVxp67_ASAP7_75t_L g298 ( .A(n_292), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_294), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_294), .B(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_294), .B(n_361), .Y(n_400) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_298), .Y(n_324) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g414 ( .A(n_303), .B(n_334), .Y(n_414) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g392 ( .A(n_309), .Y(n_392) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OAI322xp33_ASAP7_75t_SL g312 ( .A1(n_313), .A2(n_318), .A3(n_319), .B1(n_320), .B2(n_323), .C1(n_325), .C2(n_327), .Y(n_312) );
OAI322xp33_ASAP7_75t_L g394 ( .A1(n_313), .A2(n_395), .A3(n_396), .B1(n_397), .B2(n_398), .C1(n_399), .C2(n_401), .Y(n_394) );
CKINVDCx16_ASAP7_75t_R g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx4_ASAP7_75t_L g328 ( .A(n_315), .Y(n_328) );
AND2x2_ASAP7_75t_L g389 ( .A(n_315), .B(n_341), .Y(n_389) );
AND2x2_ASAP7_75t_L g402 ( .A(n_315), .B(n_403), .Y(n_402) );
CKINVDCx16_ASAP7_75t_R g413 ( .A(n_318), .Y(n_413) );
INVx1_ASAP7_75t_L g391 ( .A(n_319), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
OR2x2_ASAP7_75t_L g325 ( .A(n_321), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g408 ( .A(n_321), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_321), .B(n_362), .Y(n_419) );
OR2x2_ASAP7_75t_L g352 ( .A(n_324), .B(n_353), .Y(n_352) );
INVxp33_ASAP7_75t_L g369 ( .A(n_324), .Y(n_369) );
OAI221xp5_ASAP7_75t_SL g329 ( .A1(n_328), .A2(n_330), .B1(n_332), .B2(n_336), .C(n_338), .Y(n_329) );
NOR2xp67_ASAP7_75t_L g385 ( .A(n_328), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g412 ( .A(n_328), .Y(n_412) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
INVx3_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
AOI322xp5_ASAP7_75t_L g376 ( .A1(n_335), .A2(n_360), .A3(n_377), .B1(n_379), .B2(n_380), .C1(n_383), .C2(n_387), .Y(n_376) );
INVxp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .B1(n_346), .B2(n_347), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_372), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_350), .B(n_365), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_353), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
NAND2xp33_ASAP7_75t_SL g370 ( .A(n_356), .B(n_367), .Y(n_370) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
OAI322xp33_ASAP7_75t_L g410 ( .A1(n_358), .A2(n_411), .A3(n_413), .B1(n_414), .B2(n_415), .C1(n_417), .C2(n_420), .Y(n_410) );
AOI21xp33_ASAP7_75t_SL g359 ( .A1(n_360), .A2(n_361), .B(n_363), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_368), .B(n_416), .Y(n_425) );
OAI211xp5_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_374), .B(n_376), .C(n_388), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR4xp25_ASAP7_75t_L g393 ( .A(n_394), .B(n_404), .C(n_410), .D(n_422), .Y(n_393) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
CKINVDCx14_ASAP7_75t_R g420 ( .A(n_421), .Y(n_420) );
OAI21xp5_ASAP7_75t_SL g422 ( .A1(n_423), .A2(n_424), .B(n_425), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_426), .A2(n_449), .B1(n_453), .B2(n_456), .Y(n_448) );
INVx1_ASAP7_75t_L g435 ( .A(n_427), .Y(n_435) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g757 ( .A(n_428), .Y(n_757) );
BUFx2_ASAP7_75t_L g760 ( .A(n_428), .Y(n_760) );
NOR2x2_ASAP7_75t_L g752 ( .A(n_429), .B(n_455), .Y(n_752) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g454 ( .A(n_430), .B(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_442), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_SL g755 ( .A(n_441), .B(n_443), .Y(n_755) );
OA21x2_ASAP7_75t_L g759 ( .A1(n_441), .A2(n_442), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVxp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g748 ( .A(n_452), .Y(n_748) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx6_ASAP7_75t_L g749 ( .A(n_454), .Y(n_749) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_661), .Y(n_457) );
NAND5xp2_ASAP7_75t_L g458 ( .A(n_459), .B(n_580), .C(n_595), .D(n_621), .E(n_643), .Y(n_458) );
NOR2xp33_ASAP7_75t_SL g459 ( .A(n_460), .B(n_560), .Y(n_459) );
OAI221xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_501), .B1(n_533), .B2(n_549), .C(n_550), .Y(n_460) );
NOR2xp33_ASAP7_75t_SL g461 ( .A(n_462), .B(n_493), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_462), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_SL g737 ( .A(n_462), .Y(n_737) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_474), .Y(n_462) );
INVx1_ASAP7_75t_L g577 ( .A(n_463), .Y(n_577) );
AND2x2_ASAP7_75t_L g579 ( .A(n_463), .B(n_487), .Y(n_579) );
AND2x2_ASAP7_75t_L g589 ( .A(n_463), .B(n_486), .Y(n_589) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_463), .Y(n_607) );
INVx1_ASAP7_75t_L g617 ( .A(n_463), .Y(n_617) );
OR2x2_ASAP7_75t_L g655 ( .A(n_463), .B(n_554), .Y(n_655) );
INVx2_ASAP7_75t_L g705 ( .A(n_463), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_463), .B(n_553), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B(n_468), .Y(n_465) );
NOR2xp67_ASAP7_75t_L g474 ( .A(n_475), .B(n_486), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_476), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_476), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_SL g637 ( .A(n_476), .B(n_577), .Y(n_637) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_477), .Y(n_495) );
INVx2_ASAP7_75t_L g554 ( .A(n_477), .Y(n_554) );
OR2x2_ASAP7_75t_L g616 ( .A(n_477), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g555 ( .A(n_486), .B(n_497), .Y(n_555) );
AND2x2_ASAP7_75t_L g572 ( .A(n_486), .B(n_552), .Y(n_572) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g496 ( .A(n_487), .B(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g575 ( .A(n_487), .Y(n_575) );
AND2x2_ASAP7_75t_L g704 ( .A(n_487), .B(n_705), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_490), .A2(n_518), .B(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_490), .A2(n_529), .B(n_530), .C(n_531), .Y(n_528) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_492), .A2(n_538), .B(n_541), .Y(n_537) );
INVx1_ASAP7_75t_L g549 ( .A(n_493), .Y(n_549) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_496), .Y(n_493) );
AND2x2_ASAP7_75t_L g667 ( .A(n_494), .B(n_555), .Y(n_667) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g668 ( .A(n_495), .B(n_579), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_L g635 ( .A1(n_496), .A2(n_636), .B(n_638), .C(n_640), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_496), .B(n_636), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_496), .A2(n_566), .B1(n_709), .B2(n_710), .C(n_712), .Y(n_708) );
INVx1_ASAP7_75t_L g552 ( .A(n_497), .Y(n_552) );
INVx1_ASAP7_75t_L g588 ( .A(n_497), .Y(n_588) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_497), .Y(n_597) );
INVx1_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_511), .Y(n_502) );
AND2x2_ASAP7_75t_L g614 ( .A(n_503), .B(n_559), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_503), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_504), .B(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g706 ( .A(n_504), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g738 ( .A(n_504), .Y(n_738) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g568 ( .A(n_505), .Y(n_568) );
AND2x2_ASAP7_75t_L g594 ( .A(n_505), .B(n_548), .Y(n_594) );
NOR2x1_ASAP7_75t_L g603 ( .A(n_505), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g610 ( .A(n_505), .B(n_611), .Y(n_610) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g546 ( .A(n_506), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_511), .B(n_650), .Y(n_685) );
INVx1_ASAP7_75t_SL g689 ( .A(n_511), .Y(n_689) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_522), .Y(n_511) );
INVx3_ASAP7_75t_L g548 ( .A(n_512), .Y(n_548) );
AND2x2_ASAP7_75t_L g559 ( .A(n_512), .B(n_536), .Y(n_559) );
AND2x2_ASAP7_75t_L g581 ( .A(n_512), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g626 ( .A(n_512), .B(n_620), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_512), .B(n_558), .Y(n_707) );
INVx2_ASAP7_75t_L g529 ( .A(n_520), .Y(n_529) );
AND2x2_ASAP7_75t_L g547 ( .A(n_522), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g558 ( .A(n_522), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_522), .B(n_536), .Y(n_583) );
AND2x2_ASAP7_75t_L g619 ( .A(n_522), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_547), .Y(n_534) );
INVx1_ASAP7_75t_L g599 ( .A(n_535), .Y(n_599) );
AND2x2_ASAP7_75t_L g641 ( .A(n_535), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_535), .B(n_562), .Y(n_647) );
AOI21xp5_ASAP7_75t_SL g721 ( .A1(n_535), .A2(n_553), .B(n_576), .Y(n_721) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_545), .Y(n_535) );
OR2x2_ASAP7_75t_L g564 ( .A(n_536), .B(n_545), .Y(n_564) );
AND2x2_ASAP7_75t_L g611 ( .A(n_536), .B(n_548), .Y(n_611) );
INVx2_ASAP7_75t_L g620 ( .A(n_536), .Y(n_620) );
INVx1_ASAP7_75t_L g726 ( .A(n_536), .Y(n_726) );
AND2x2_ASAP7_75t_L g650 ( .A(n_545), .B(n_620), .Y(n_650) );
INVx1_ASAP7_75t_L g675 ( .A(n_545), .Y(n_675) );
AND2x2_ASAP7_75t_L g584 ( .A(n_547), .B(n_568), .Y(n_584) );
AND2x2_ASAP7_75t_L g596 ( .A(n_547), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_SL g714 ( .A(n_547), .Y(n_714) );
INVx2_ASAP7_75t_L g604 ( .A(n_548), .Y(n_604) );
AND2x2_ASAP7_75t_L g642 ( .A(n_548), .B(n_558), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_548), .B(n_726), .Y(n_725) );
OAI21xp33_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_555), .B(n_556), .Y(n_550) );
AND2x2_ASAP7_75t_L g657 ( .A(n_551), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g711 ( .A(n_551), .Y(n_711) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx1_ASAP7_75t_L g631 ( .A(n_552), .Y(n_631) );
BUFx2_ASAP7_75t_L g730 ( .A(n_552), .Y(n_730) );
BUFx2_ASAP7_75t_L g601 ( .A(n_553), .Y(n_601) );
AND2x2_ASAP7_75t_L g703 ( .A(n_553), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g686 ( .A(n_554), .Y(n_686) );
AND2x4_ASAP7_75t_L g613 ( .A(n_555), .B(n_576), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_555), .B(n_637), .Y(n_649) );
AOI32xp33_ASAP7_75t_L g573 ( .A1(n_556), .A2(n_574), .A3(n_576), .B1(n_578), .B2(n_579), .Y(n_573) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
INVx3_ASAP7_75t_L g562 ( .A(n_557), .Y(n_562) );
OR2x2_ASAP7_75t_L g698 ( .A(n_557), .B(n_654), .Y(n_698) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g567 ( .A(n_558), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g674 ( .A(n_558), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g566 ( .A(n_559), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g578 ( .A(n_559), .B(n_568), .Y(n_578) );
INVx1_ASAP7_75t_L g699 ( .A(n_559), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_559), .B(n_674), .Y(n_732) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_565), .B(n_569), .C(n_573), .Y(n_560) );
OAI322xp33_ASAP7_75t_L g669 ( .A1(n_561), .A2(n_606), .A3(n_670), .B1(n_672), .B2(n_676), .C1(n_677), .C2(n_681), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVxp67_ASAP7_75t_L g634 ( .A(n_562), .Y(n_634) );
INVx1_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g688 ( .A(n_564), .B(n_689), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_564), .B(n_604), .Y(n_735) );
INVxp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g627 ( .A(n_567), .Y(n_627) );
OR2x2_ASAP7_75t_L g713 ( .A(n_568), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_571), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g622 ( .A(n_572), .B(n_601), .Y(n_622) );
AND2x2_ASAP7_75t_L g693 ( .A(n_572), .B(n_606), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_572), .B(n_680), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g580 ( .A1(n_574), .A2(n_581), .B1(n_584), .B2(n_585), .C(n_590), .Y(n_580) );
OR2x2_ASAP7_75t_L g591 ( .A(n_574), .B(n_587), .Y(n_591) );
AND2x2_ASAP7_75t_L g679 ( .A(n_574), .B(n_680), .Y(n_679) );
AOI32xp33_ASAP7_75t_L g718 ( .A1(n_574), .A2(n_604), .A3(n_719), .B1(n_720), .B2(n_723), .Y(n_718) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_575), .B(n_611), .C(n_634), .Y(n_652) );
AND2x2_ASAP7_75t_L g678 ( .A(n_575), .B(n_671), .Y(n_678) );
INVxp67_ASAP7_75t_L g658 ( .A(n_576), .Y(n_658) );
BUFx3_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_579), .B(n_631), .Y(n_687) );
INVx2_ASAP7_75t_L g697 ( .A(n_579), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_579), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g666 ( .A(n_582), .Y(n_666) );
OR2x2_ASAP7_75t_L g592 ( .A(n_583), .B(n_593), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_585), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_588), .Y(n_671) );
AND2x2_ASAP7_75t_L g630 ( .A(n_589), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g676 ( .A(n_589), .Y(n_676) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_589), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AOI21xp33_ASAP7_75t_SL g615 ( .A1(n_591), .A2(n_616), .B(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g709 ( .A(n_594), .B(n_619), .Y(n_709) );
AOI211xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_598), .B(n_608), .C(n_615), .Y(n_595) );
AND2x2_ASAP7_75t_L g639 ( .A(n_597), .B(n_607), .Y(n_639) );
INVx2_ASAP7_75t_L g654 ( .A(n_597), .Y(n_654) );
OR2x2_ASAP7_75t_L g692 ( .A(n_597), .B(n_655), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_597), .B(n_735), .Y(n_734) );
AOI211xp5_ASAP7_75t_SL g598 ( .A1(n_599), .A2(n_600), .B(n_602), .C(n_605), .Y(n_598) );
INVxp67_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_601), .B(n_639), .Y(n_638) );
OAI211xp5_ASAP7_75t_L g720 ( .A1(n_602), .A2(n_697), .B(n_721), .C(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2x1p5_ASAP7_75t_L g618 ( .A(n_603), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g660 ( .A(n_604), .B(n_650), .Y(n_660) );
INVx1_ASAP7_75t_L g665 ( .A(n_604), .Y(n_665) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_609), .B(n_612), .Y(n_608) );
INVxp33_ASAP7_75t_L g716 ( .A(n_610), .Y(n_716) );
AND2x2_ASAP7_75t_L g695 ( .A(n_611), .B(n_674), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_616), .A2(n_678), .B(n_679), .Y(n_677) );
OAI322xp33_ASAP7_75t_L g696 ( .A1(n_618), .A2(n_697), .A3(n_698), .B1(n_699), .B2(n_700), .C1(n_702), .C2(n_706), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_623), .B1(n_628), .B2(n_632), .C(n_635), .Y(n_621) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g673 ( .A(n_626), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g717 ( .A(n_630), .Y(n_717) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_633), .B(n_653), .Y(n_719) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g682 ( .A(n_642), .B(n_650), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_646), .B1(n_648), .B2(n_650), .C(n_651), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_646), .A2(n_663), .B1(n_667), .B2(n_668), .C(n_669), .Y(n_662) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVxp67_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_650), .B(n_665), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_656), .B2(n_659), .Y(n_651) );
OR2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx2_ASAP7_75t_SL g680 ( .A(n_655), .Y(n_680) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND5xp2_ASAP7_75t_L g661 ( .A(n_662), .B(n_683), .C(n_708), .D(n_718), .E(n_728), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_664), .B(n_666), .Y(n_663) );
NOR4xp25_ASAP7_75t_L g736 ( .A(n_665), .B(n_671), .C(n_737), .D(n_738), .Y(n_736) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_668), .A2(n_729), .B1(n_731), .B2(n_733), .C(n_736), .Y(n_728) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g727 ( .A(n_674), .Y(n_727) );
OAI322xp33_ASAP7_75t_L g684 ( .A1(n_678), .A2(n_685), .A3(n_686), .B1(n_687), .B2(n_688), .C1(n_690), .C2(n_694), .Y(n_684) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_696), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g729 ( .A(n_704), .B(n_730), .Y(n_729) );
OAI22xp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_715), .B1(n_716), .B2(n_717), .Y(n_712) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_727), .Y(n_724) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
NAND2xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_759), .Y(n_758) );
endmodule