module real_jpeg_29484_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_0),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_0),
.A2(n_49),
.B1(n_50),
.B2(n_70),
.Y(n_79)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_3),
.A2(n_27),
.B1(n_92),
.B2(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_3),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_3),
.A2(n_27),
.B1(n_49),
.B2(n_50),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_5),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_6),
.A2(n_36),
.B1(n_49),
.B2(n_50),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_7),
.A2(n_49),
.B1(n_50),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_7),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_9),
.A2(n_49),
.B1(n_50),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_9),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_59),
.Y(n_104)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_11),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_11),
.B(n_24),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_11),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_11),
.A2(n_24),
.B(n_76),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_94),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_11),
.A2(n_50),
.B(n_63),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_11),
.B(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_11),
.A2(n_47),
.B1(n_86),
.B2(n_162),
.Y(n_164)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_14),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_67),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_14),
.A2(n_49),
.B1(n_50),
.B2(n_67),
.Y(n_148)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_15),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_116),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_114),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_81),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_19),
.B(n_81),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_60),
.C(n_72),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_20),
.A2(n_21),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_37),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_22),
.B(n_38),
.C(n_44),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_23),
.A2(n_28),
.B1(n_31),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_24),
.A2(n_25),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_24),
.B(n_41),
.Y(n_90)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI32xp33_ASAP7_75t_L g73 ( 
.A1(n_25),
.A2(n_32),
.A3(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_25),
.A2(n_90),
.B1(n_91),
.B2(n_95),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_28),
.A2(n_31),
.B1(n_35),
.B2(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_31),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_32),
.A2(n_33),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_33),
.B(n_75),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_33),
.A2(n_64),
.B(n_94),
.C(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_40),
.A2(n_91),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_40),
.A2(n_41),
.B(n_92),
.C(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_41),
.B(n_92),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_48),
.B(n_53),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_48),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_46),
.B(n_79),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_46),
.A2(n_54),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_58),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_47),
.A2(n_86),
.B1(n_154),
.B2(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_47),
.B(n_94),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_55),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_50),
.B1(n_63),
.B2(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_49),
.B(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_60),
.B(n_72),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_66),
.B(n_68),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_61),
.A2(n_102),
.B(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_61),
.A2(n_65),
.B1(n_66),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_61),
.A2(n_65),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_61),
.A2(n_65),
.B1(n_126),
.B2(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_65),
.B(n_94),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_71),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_78),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_78),
.Y(n_120)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_98),
.B1(n_99),
.B2(n_113),
.Y(n_81)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_96),
.B2(n_97),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_86),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

HAxp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_94),
.CON(n_91),
.SN(n_91)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_109),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_101),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_130),
.B(n_176),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_127),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_118),
.B(n_127),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.C(n_124),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_119),
.A2(n_120),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_170),
.B(n_175),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_150),
.B(n_169),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_133),
.B(n_140),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_138),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_135),
.B1(n_138),
.B2(n_157),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_138),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_147),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_146),
.C(n_147),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_148),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_158),
.B(n_168),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_156),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_152),
.B(n_156),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_163),
.B(n_167),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_160),
.B(n_161),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_171),
.B(n_172),
.Y(n_175)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);


endmodule