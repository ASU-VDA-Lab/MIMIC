module real_jpeg_51_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_215;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_216;
wire n_128;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_1),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_4),
.A2(n_29),
.B1(n_32),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_4),
.A2(n_41),
.B1(n_45),
.B2(n_56),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_56),
.Y(n_109)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_7),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_7),
.A2(n_34),
.B1(n_41),
.B2(n_45),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_7),
.B(n_23),
.C(n_29),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_7),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_7),
.B(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_7),
.B(n_41),
.C(n_59),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_7),
.B(n_44),
.C(n_48),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_7),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_7),
.B(n_85),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_7),
.B(n_46),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_8),
.A2(n_41),
.B1(n_45),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_8),
.A2(n_29),
.B1(n_32),
.B2(n_53),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_93),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_92),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_68),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_15),
.B(n_68),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_65),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_35),
.B2(n_36),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_19),
.A2(n_20),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_19),
.A2(n_81),
.B(n_91),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_19),
.A2(n_20),
.B1(n_83),
.B2(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_19),
.B(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_19),
.A2(n_20),
.B1(n_75),
.B2(n_113),
.Y(n_125)
);

AOI211xp5_ASAP7_75t_SL g139 ( 
.A1(n_19),
.A2(n_111),
.B(n_115),
.C(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_19),
.A2(n_20),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_37),
.C(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_20),
.B(n_75),
.Y(n_115)
);

AO21x2_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_28),
.B(n_33),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_25),
.B(n_129),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_28),
.Y(n_161)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_29),
.A2(n_32),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_29),
.B(n_175),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_36)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_37),
.A2(n_63),
.B1(n_66),
.B2(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_51),
.B(n_52),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_38),
.A2(n_51),
.B1(n_78),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_39),
.A2(n_46),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_39),
.A2(n_46),
.B(n_90),
.Y(n_111)
);

NOR2x1_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_40)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

OA22x2_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_45),
.B1(n_59),
.B2(n_60),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_41),
.B(n_186),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AO22x1_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_85),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_48),
.B(n_197),
.Y(n_196)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_57),
.B1(n_61),
.B2(n_67),
.Y(n_66)
);

AO21x2_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_61),
.B(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_59),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_61),
.Y(n_192)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.C(n_80),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_73),
.B1(n_74),
.B2(n_97),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_75),
.B(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_75),
.B(n_136),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_75),
.A2(n_111),
.B1(n_113),
.B2(n_136),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_75),
.B(n_131),
.C(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_75),
.A2(n_113),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_82),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_83),
.A2(n_88),
.B1(n_91),
.B2(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_88),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_116),
.B(n_237),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_95),
.B(n_98),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.C(n_104),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_99),
.Y(n_234)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_104),
.A2(n_105),
.B1(n_233),
.B2(n_235),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_112),
.B(n_114),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_106),
.A2(n_124),
.B1(n_125),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_106),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_111),
.B1(n_136),
.B2(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_107),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_132),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_134)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_135),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_111),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_111),
.A2(n_136),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_111),
.A2(n_136),
.B1(n_184),
.B2(n_185),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_111),
.A2(n_113),
.B(n_140),
.C(n_207),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_111),
.A2(n_136),
.B1(n_172),
.B2(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_114),
.B(n_126),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_112),
.A2(n_114),
.B(n_145),
.Y(n_219)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21x1_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_230),
.B(n_236),
.Y(n_117)
);

AOI21x1_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_216),
.B(n_229),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_163),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_149),
.B(n_162),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_SL g163 ( 
.A(n_121),
.B(n_164),
.C(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_141),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_141),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_134),
.C(n_138),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_133),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_124),
.A2(n_125),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_130),
.A2(n_131),
.B1(n_160),
.B2(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_130),
.A2(n_131),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_130),
.B(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_130),
.A2(n_131),
.B1(n_173),
.B2(n_174),
.Y(n_207)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_131),
.B(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_131),
.B(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_131),
.B(n_136),
.C(n_191),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_134),
.A2(n_138),
.B1(n_139),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_135),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_168),
.C(n_172),
.Y(n_167)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_142),
.B(n_144),
.C(n_147),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_153),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_158),
.C(n_159),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_154),
.A2(n_155),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_156),
.A2(n_157),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_179),
.B(n_215),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_176),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_167),
.B(n_176),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_209),
.B(n_214),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_203),
.B(n_208),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_193),
.B(n_202),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_187),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_200),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_205),
.Y(n_208)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_211),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_217),
.B(n_218),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_228),
.Y(n_218)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_226),
.C(n_228),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_232),
.Y(n_236)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);


endmodule