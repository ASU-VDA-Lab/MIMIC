module fake_jpeg_3803_n_252 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_18),
.Y(n_32)
);

AO22x1_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_18),
.B1(n_27),
.B2(n_15),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_1),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_24),
.B1(n_21),
.B2(n_27),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_30),
.B1(n_16),
.B2(n_29),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_47),
.B1(n_51),
.B2(n_58),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_42),
.A2(n_30),
.B1(n_16),
.B2(n_29),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_48),
.B1(n_55),
.B2(n_63),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_30),
.B1(n_26),
.B2(n_29),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_17),
.B1(n_28),
.B2(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_23),
.B1(n_28),
.B2(n_20),
.Y(n_51)
);

AO22x1_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_40),
.B1(n_38),
.B2(n_33),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_17),
.B1(n_28),
.B2(n_20),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_57),
.Y(n_75)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_32),
.A2(n_23),
.B1(n_17),
.B2(n_25),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_27),
.B1(n_15),
.B2(n_22),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_37),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_33),
.A2(n_25),
.B1(n_24),
.B2(n_21),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_74),
.Y(n_88)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_21),
.B1(n_31),
.B2(n_33),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_45),
.B1(n_47),
.B2(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_80),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_40),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_60),
.B(n_61),
.Y(n_91)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_31),
.B1(n_3),
.B2(n_4),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_78),
.Y(n_92)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_57),
.A2(n_31),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_82),
.Y(n_96)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_56),
.B1(n_53),
.B2(n_49),
.Y(n_106)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_101),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_69),
.B1(n_75),
.B2(n_80),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_44),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_95),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_73),
.B(n_67),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_54),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_54),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_61),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_22),
.Y(n_127)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_78),
.Y(n_102)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_105),
.A2(n_68),
.B1(n_74),
.B2(n_83),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_70),
.B1(n_96),
.B2(n_97),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_107),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_127),
.B(n_95),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_109),
.B(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_112),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_116),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_121),
.B1(n_106),
.B2(n_96),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_125),
.B1(n_92),
.B2(n_105),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_84),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_92),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_59),
.B1(n_77),
.B2(n_53),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_150),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_147),
.B(n_27),
.Y(n_164)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_135),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_134),
.B1(n_114),
.B2(n_102),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_128),
.A2(n_85),
.B1(n_101),
.B2(n_94),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_143),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_142),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_118),
.B1(n_120),
.B2(n_112),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_101),
.C(n_104),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_148),
.C(n_114),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_126),
.B(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_43),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_107),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_102),
.B1(n_77),
.B2(n_83),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_145),
.A2(n_111),
.B1(n_110),
.B2(n_77),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_108),
.A2(n_43),
.B(n_33),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_50),
.C(n_38),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_153),
.B1(n_165),
.B2(n_167),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_155),
.B(n_158),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_159),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_148),
.C(n_147),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_171),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_149),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_162),
.A2(n_103),
.B1(n_90),
.B2(n_27),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_169),
.B(n_130),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_144),
.A2(n_136),
.B1(n_140),
.B2(n_132),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_50),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_40),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_103),
.B1(n_40),
.B2(n_38),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_27),
.B(n_15),
.Y(n_169)
);

NOR2x1_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_134),
.Y(n_171)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_180),
.C(n_191),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_189),
.B(n_5),
.Y(n_205)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_185),
.Y(n_198)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

XNOR2x1_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_38),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_169),
.C(n_166),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_2),
.Y(n_188)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_164),
.A2(n_90),
.B(n_103),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_2),
.Y(n_190)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_90),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_156),
.B1(n_162),
.B2(n_157),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_194),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_176),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_175),
.A2(n_172),
.B1(n_167),
.B2(n_14),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_181),
.Y(n_219)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_202),
.B(n_203),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_178),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_2),
.B(n_5),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_204),
.A2(n_205),
.B(n_188),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_14),
.C(n_7),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_190),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_219),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_200),
.A2(n_175),
.B1(n_174),
.B2(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_186),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_213),
.C(n_216),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_189),
.B1(n_184),
.B2(n_179),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_211),
.A2(n_193),
.B1(n_201),
.B2(n_183),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_198),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_193),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_173),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_215),
.A2(n_217),
.B(n_204),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_180),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_195),
.C(n_206),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_207),
.B(n_173),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

AO22x1_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_197),
.B1(n_205),
.B2(n_196),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_208),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_225),
.C(n_213),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_228),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_199),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_235),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_232),
.A2(n_233),
.B(n_228),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_183),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_218),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_237),
.C(n_8),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_210),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_227),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_238),
.A2(n_240),
.B(n_242),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_224),
.B(n_222),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_243),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_6),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_238),
.A2(n_234),
.B1(n_10),
.B2(n_11),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

AOI322xp5_ASAP7_75t_L g247 ( 
.A1(n_241),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_239),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_246),
.C(n_244),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_248),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_9),
.Y(n_252)
);


endmodule