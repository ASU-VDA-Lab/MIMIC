module fake_jpeg_16771_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_SL g7 ( 
.A(n_6),
.B(n_1),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_6),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_11),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_9),
.A2(n_2),
.B(n_3),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_23),
.C(n_18),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_2),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVxp33_ASAP7_75t_SL g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_31),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_13),
.B1(n_8),
.B2(n_14),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_26),
.A2(n_28),
.B(n_32),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_13),
.B1(n_14),
.B2(n_12),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_12),
.C(n_3),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_35),
.C(n_36),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_5),
.B(n_31),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_28),
.C(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_39),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_27),
.C(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_34),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_44),
.B(n_27),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_40),
.B(n_24),
.Y(n_46)
);


endmodule