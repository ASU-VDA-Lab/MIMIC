module real_jpeg_6209_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_1),
.A2(n_118),
.B1(n_122),
.B2(n_125),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_1),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_1),
.A2(n_125),
.B1(n_199),
.B2(n_202),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_2),
.Y(n_112)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_2),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_2),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_3),
.A2(n_167),
.B1(n_172),
.B2(n_176),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_3),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_3),
.A2(n_176),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_4),
.A2(n_199),
.B1(n_219),
.B2(n_222),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_4),
.Y(n_222)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_5),
.A2(n_50),
.B1(n_81),
.B2(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_5),
.B(n_257),
.C(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_5),
.B(n_77),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_5),
.B(n_161),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_5),
.B(n_105),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_5),
.B(n_321),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_6),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_6),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_6),
.A2(n_100),
.B1(n_167),
.B2(n_262),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_6),
.A2(n_100),
.B1(n_138),
.B2(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_7),
.A2(n_30),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_7),
.A2(n_57),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_7),
.A2(n_57),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_7),
.A2(n_57),
.B1(n_113),
.B2(n_162),
.Y(n_264)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_9),
.Y(n_161)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_9),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_10),
.A2(n_167),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_10),
.Y(n_183)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_11),
.Y(n_151)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_13),
.A2(n_90),
.B1(n_94),
.B2(n_95),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_13),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_13),
.A2(n_29),
.B1(n_95),
.B2(n_234),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_13),
.A2(n_95),
.B1(n_251),
.B2(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_13),
.A2(n_95),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_15),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_15),
.Y(n_116)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_15),
.Y(n_136)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_242),
.B1(n_243),
.B2(n_361),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_18),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_241),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_205),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_20),
.B(n_205),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_140),
.C(n_187),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_21),
.B(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_62),
.B2(n_139),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_22),
.B(n_63),
.C(n_103),
.Y(n_225)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_45),
.B(n_54),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_24),
.B(n_56),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_35),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_36),
.B1(n_39),
.B2(n_43),
.Y(n_35)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_37),
.B(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_40),
.Y(n_193)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_41),
.Y(n_323)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_42),
.Y(n_154)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_42),
.Y(n_195)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_44),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_50),
.B(n_51),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_49),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_50),
.B(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_50),
.A2(n_157),
.B(n_263),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_SL g317 ( 
.A1(n_50),
.A2(n_318),
.B(n_319),
.Y(n_317)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_51),
.A2(n_144),
.A3(n_147),
.B1(n_149),
.B2(n_152),
.Y(n_143)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_61),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_60),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_61),
.Y(n_204)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_103),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_89),
.B1(n_96),
.B2(n_97),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_64),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_77),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_68),
.B1(n_71),
.B2(n_75),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_70),
.Y(n_332)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_77),
.Y(n_96)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_84),
.B2(n_87),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_80),
.Y(n_336)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_83),
.Y(n_339)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_86),
.Y(n_213)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_86),
.Y(n_272)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_89),
.A2(n_96),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_96),
.B(n_191),
.Y(n_240)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_97),
.Y(n_239)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_117),
.B(n_126),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_104),
.A2(n_117),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_104),
.A2(n_209),
.B1(n_268),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_105),
.B(n_127),
.Y(n_253)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_106),
.A2(n_126),
.B(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_113),
.B2(n_115),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_130),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_134),
.B1(n_137),
.B2(n_138),
.Y(n_131)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_133),
.B(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_136),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_140),
.A2(n_141),
.B1(n_187),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_155),
.B2(n_156),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_143),
.B(n_155),
.Y(n_229)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_153),
.Y(n_318)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_165),
.B1(n_177),
.B2(n_181),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_157),
.A2(n_261),
.B(n_263),
.Y(n_260)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_158),
.A2(n_160),
.B1(n_166),
.B2(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_158),
.A2(n_182),
.B1(n_217),
.B2(n_223),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_158),
.B(n_264),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_158),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

INVx3_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_161),
.Y(n_224)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_170),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_174),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx8_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_175),
.Y(n_288)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_180),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_184),
.B(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_187),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_197),
.C(n_203),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_188),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_196),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_196),
.A2(n_239),
.B(n_240),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_196),
.A2(n_240),
.B(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_197),
.B(n_203),
.Y(n_352)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_198),
.Y(n_326)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_199),
.Y(n_284)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_233),
.B(n_236),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_228),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_216),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_209),
.A2(n_250),
.B(n_253),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_209),
.A2(n_253),
.B(n_312),
.Y(n_349)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_212),
.Y(n_314)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_224),
.A2(n_292),
.B(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_237),
.B2(n_238),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI21x1_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_355),
.B(n_360),
.Y(n_243)
);

AO21x1_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_344),
.B(n_354),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_306),
.B(n_343),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_275),
.B(n_305),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_259),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_248),
.B(n_259),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_249),
.A2(n_254),
.B1(n_255),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_249),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_265),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_260),
.B(n_266),
.C(n_274),
.Y(n_307)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_273),
.B2(n_274),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_271),
.Y(n_333)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_295),
.B(n_304),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_281),
.B(n_294),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_293),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_293),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_289),
.B(n_292),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_302),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_302),
.Y(n_304)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_308),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_324),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_315),
.B2(n_316),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_311),
.B(n_315),
.C(n_324),
.Y(n_345)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

AOI32xp33_ASAP7_75t_L g327 ( 
.A1(n_320),
.A2(n_328),
.A3(n_333),
.B1(n_334),
.B2(n_337),
.Y(n_327)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_327),
.Y(n_350)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx5_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx8_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx6_ASAP7_75t_L g342 ( 
.A(n_336),
.Y(n_342)
);

NAND2xp33_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_340),
.Y(n_337)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_345),
.B(n_346),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_351),
.B2(n_353),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_350),
.C(n_353),
.Y(n_356)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_351),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_356),
.B(n_357),
.Y(n_360)
);


endmodule