module real_aes_3738_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_592;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_417;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_552;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_859;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1161;
wire n_686;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1162;
wire n_762;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_414;
wire n_776;
wire n_1138;
wire n_890;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1289;
wire n_937;
wire n_773;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_816;
wire n_625;
wire n_953;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1050;
wire n_426;
wire n_1134;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1060;
wire n_1154;
wire n_632;
wire n_714;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1033;
wire n_1028;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_974;
wire n_857;
wire n_376;
wire n_491;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1198;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_698;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_483;
wire n_1280;
wire n_394;
wire n_729;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g609 ( .A(n_0), .Y(n_609) );
INVx1_ASAP7_75t_L g697 ( .A(n_1), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_2), .A2(n_361), .B1(n_526), .B2(n_857), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_3), .A2(n_308), .B1(n_741), .B2(n_851), .Y(n_850) );
AOI21xp33_ASAP7_75t_SL g893 ( .A1(n_4), .A2(n_894), .B(n_895), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_5), .A2(n_359), .B1(n_565), .B2(n_567), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_6), .A2(n_188), .B1(n_605), .B2(n_857), .Y(n_1248) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_7), .A2(n_203), .B1(n_539), .B2(n_540), .Y(n_955) );
AO22x1_ASAP7_75t_L g930 ( .A1(n_8), .A2(n_234), .B1(n_536), .B2(n_537), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_9), .A2(n_275), .B1(n_513), .B2(n_819), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_10), .A2(n_318), .B1(n_513), .B2(n_514), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_11), .A2(n_311), .B1(n_450), .B2(n_526), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_12), .A2(n_209), .B1(n_558), .B2(n_567), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_13), .A2(n_131), .B1(n_485), .B2(n_552), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_14), .A2(n_28), .B1(n_536), .B2(n_537), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_15), .A2(n_44), .B1(n_598), .B2(n_599), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_16), .A2(n_344), .B1(n_623), .B2(n_911), .Y(n_910) );
AOI21xp33_ASAP7_75t_SL g977 ( .A1(n_17), .A2(n_619), .B(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g621 ( .A(n_18), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g939 ( .A1(n_19), .A2(n_221), .B1(n_446), .B2(n_539), .Y(n_939) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_20), .B(n_404), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_21), .A2(n_179), .B1(n_502), .B2(n_982), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_22), .A2(n_313), .B1(n_666), .B2(n_667), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_23), .A2(n_192), .B1(n_477), .B2(n_513), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_24), .A2(n_129), .B1(n_558), .B2(n_561), .Y(n_576) );
OAI22x1_ASAP7_75t_L g747 ( .A1(n_25), .A2(n_748), .B1(n_779), .B2(n_780), .Y(n_747) );
INVx1_ASAP7_75t_L g780 ( .A(n_25), .Y(n_780) );
AOI21xp33_ASAP7_75t_L g948 ( .A1(n_26), .A2(n_705), .B(n_949), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_27), .A2(n_341), .B1(n_517), .B2(n_775), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g1283 ( .A1(n_29), .A2(n_302), .B1(n_450), .B2(n_526), .Y(n_1283) );
AOI221xp5_ASAP7_75t_L g1273 ( .A1(n_30), .A2(n_294), .B1(n_1274), .B2(n_1275), .C(n_1276), .Y(n_1273) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_31), .Y(n_404) );
INVx1_ASAP7_75t_L g690 ( .A(n_32), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_33), .A2(n_96), .B1(n_539), .B2(n_797), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_34), .A2(n_360), .B1(n_443), .B2(n_446), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_35), .A2(n_126), .B1(n_770), .B2(n_772), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g1017 ( .A1(n_36), .A2(n_271), .B1(n_1018), .B2(n_1020), .Y(n_1017) );
AO22x1_ASAP7_75t_L g647 ( .A1(n_37), .A2(n_156), .B1(n_489), .B2(n_648), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_38), .A2(n_41), .B1(n_428), .B2(n_905), .Y(n_987) );
INVx1_ASAP7_75t_L g950 ( .A(n_39), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_40), .A2(n_151), .B1(n_522), .B2(n_718), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g1035 ( .A1(n_42), .A2(n_196), .B1(n_1018), .B2(n_1020), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_43), .B(n_701), .Y(n_960) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_45), .A2(n_351), .B1(n_1022), .B2(n_1028), .Y(n_1027) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_46), .A2(n_159), .B1(n_450), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_47), .A2(n_94), .B1(n_598), .B2(n_866), .Y(n_865) );
AO22x2_ASAP7_75t_L g595 ( .A1(n_48), .A2(n_596), .B1(n_606), .B2(n_634), .Y(n_595) );
INVxp33_ASAP7_75t_SL g633 ( .A(n_48), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_49), .A2(n_207), .B1(n_1005), .B2(n_1009), .Y(n_1004) );
INVx1_ASAP7_75t_L g487 ( .A(n_50), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_51), .A2(n_152), .B1(n_398), .B2(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_52), .A2(n_61), .B1(n_1012), .B2(n_1015), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_53), .A2(n_214), .B1(n_518), .B2(n_603), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g1284 ( .A1(n_54), .A2(n_357), .B1(n_603), .B2(n_1285), .Y(n_1284) );
INVx1_ASAP7_75t_L g559 ( .A(n_55), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_56), .A2(n_107), .B1(n_398), .B2(n_601), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_57), .A2(n_643), .B(n_647), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_58), .A2(n_242), .B1(n_450), .B2(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_59), .B(n_872), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_60), .A2(n_326), .B1(n_517), .B2(n_599), .Y(n_840) );
AOI22xp33_ASAP7_75t_SL g653 ( .A1(n_62), .A2(n_73), .B1(n_654), .B2(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g554 ( .A(n_63), .Y(n_554) );
OA22x2_ASAP7_75t_L g410 ( .A1(n_64), .A2(n_160), .B1(n_404), .B2(n_408), .Y(n_410) );
INVx1_ASAP7_75t_L g438 ( .A(n_64), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g942 ( .A1(n_65), .A2(n_117), .B1(n_454), .B2(n_943), .Y(n_942) );
AOI22xp5_ASAP7_75t_L g842 ( .A1(n_66), .A2(n_223), .B1(n_450), .B2(n_526), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_67), .A2(n_374), .B1(n_398), .B2(n_598), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_68), .A2(n_135), .B1(n_868), .B2(n_1246), .Y(n_1245) );
AOI22xp5_ASAP7_75t_L g1021 ( .A1(n_69), .A2(n_290), .B1(n_1022), .B2(n_1023), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_70), .A2(n_78), .B1(n_463), .B2(n_623), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g1282 ( .A1(n_71), .A2(n_113), .B1(n_398), .B2(n_423), .Y(n_1282) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_72), .A2(n_171), .B1(n_658), .B2(n_659), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_74), .A2(n_137), .B1(n_428), .B2(n_431), .Y(n_727) );
INVx1_ASAP7_75t_L g979 ( .A(n_75), .Y(n_979) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_76), .A2(n_353), .B1(n_536), .B2(n_537), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g1286 ( .A1(n_77), .A2(n_194), .B1(n_428), .B2(n_601), .Y(n_1286) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_79), .A2(n_237), .B1(n_651), .B2(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_80), .A2(n_248), .B1(n_536), .B2(n_537), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_81), .A2(n_174), .B1(n_539), .B2(n_540), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_82), .A2(n_285), .B1(n_502), .B2(n_982), .Y(n_1255) );
INVx1_ASAP7_75t_L g1139 ( .A(n_83), .Y(n_1139) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_84), .A2(n_231), .B1(n_540), .B2(n_544), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_85), .A2(n_139), .B1(n_474), .B2(n_477), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_86), .A2(n_372), .B1(n_543), .B2(n_544), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_87), .A2(n_306), .B1(n_398), .B2(n_524), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_88), .B(n_177), .Y(n_385) );
INVx1_ASAP7_75t_L g407 ( .A(n_88), .Y(n_407) );
OAI21xp33_ASAP7_75t_L g439 ( .A1(n_88), .A2(n_160), .B(n_440), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_89), .A2(n_230), .B1(n_543), .B2(n_547), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_90), .A2(n_243), .B1(n_428), .B2(n_431), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_91), .A2(n_358), .B1(n_474), .B2(n_477), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g871 ( .A1(n_92), .A2(n_872), .B(n_873), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_93), .A2(n_363), .B1(n_630), .B2(n_631), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_95), .A2(n_249), .B1(n_775), .B2(n_776), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_97), .A2(n_224), .B1(n_539), .B2(n_546), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_98), .B(n_848), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_99), .A2(n_181), .B1(n_428), .B2(n_603), .Y(n_602) );
INVxp33_ASAP7_75t_L g1054 ( .A(n_100), .Y(n_1054) );
AND2x4_ASAP7_75t_L g1008 ( .A(n_101), .B(n_276), .Y(n_1008) );
INVx1_ASAP7_75t_L g1014 ( .A(n_101), .Y(n_1014) );
INVx1_ASAP7_75t_L g760 ( .A(n_102), .Y(n_760) );
INVx1_ASAP7_75t_L g814 ( .A(n_103), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_104), .A2(n_218), .B1(n_546), .B2(n_547), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g927 ( .A1(n_105), .A2(n_332), .B1(n_539), .B2(n_540), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_106), .A2(n_267), .B1(n_558), .B2(n_561), .Y(n_921) );
AOI21xp5_ASAP7_75t_L g1252 ( .A1(n_108), .A2(n_460), .B(n_1253), .Y(n_1252) );
OAI22xp5_ASAP7_75t_L g1268 ( .A1(n_109), .A2(n_1269), .B1(n_1270), .B2(n_1287), .Y(n_1268) );
INVx1_ASAP7_75t_L g1287 ( .A(n_109), .Y(n_1287) );
INVx1_ASAP7_75t_L g674 ( .A(n_110), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g989 ( .A1(n_111), .A2(n_286), .B1(n_768), .B2(n_868), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_112), .A2(n_331), .B1(n_460), .B2(n_630), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_114), .A2(n_253), .B1(n_460), .B2(n_463), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g799 ( .A1(n_115), .A2(n_301), .B1(n_485), .B2(n_552), .C(n_800), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g965 ( .A1(n_116), .A2(n_258), .B1(n_565), .B2(n_567), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_118), .B(n_485), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_119), .A2(n_162), .B1(n_502), .B2(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g1007 ( .A(n_120), .Y(n_1007) );
AND2x4_ASAP7_75t_L g1010 ( .A(n_120), .B(n_381), .Y(n_1010) );
INVx1_ASAP7_75t_SL g1019 ( .A(n_120), .Y(n_1019) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_121), .A2(n_150), .B1(n_524), .B2(n_718), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_122), .A2(n_278), .B1(n_661), .B2(n_662), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_123), .A2(n_322), .B1(n_598), .B2(n_718), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g1039 ( .A1(n_124), .A2(n_239), .B1(n_1022), .B2(n_1023), .Y(n_1039) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_125), .A2(n_250), .B1(n_565), .B2(n_680), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_127), .A2(n_314), .B1(n_428), .B2(n_905), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_128), .A2(n_342), .B1(n_565), .B2(n_567), .Y(n_803) );
INVx1_ASAP7_75t_L g801 ( .A(n_130), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_132), .A2(n_169), .B1(n_650), .B2(n_651), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g1257 ( .A1(n_133), .A2(n_282), .B1(n_652), .B2(n_984), .Y(n_1257) );
XOR2x2_ASAP7_75t_L g639 ( .A(n_134), .B(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_134), .A2(n_281), .B1(n_1005), .B2(n_1009), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_136), .A2(n_187), .B1(n_868), .B2(n_869), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_138), .A2(n_315), .B1(n_443), .B2(n_518), .Y(n_900) );
XNOR2x1_ASAP7_75t_L g394 ( .A(n_140), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g735 ( .A(n_141), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g1247 ( .A1(n_142), .A2(n_355), .B1(n_863), .B2(n_991), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_143), .A2(n_144), .B1(n_546), .B2(n_547), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_145), .A2(n_254), .B1(n_428), .B2(n_720), .Y(n_719) );
AO22x1_ASAP7_75t_L g928 ( .A1(n_146), .A2(n_291), .B1(n_546), .B2(n_547), .Y(n_928) );
INVx1_ASAP7_75t_L g852 ( .A(n_147), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_148), .A2(n_352), .B1(n_546), .B2(n_547), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_149), .A2(n_297), .B1(n_659), .B2(n_662), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_153), .A2(n_316), .B1(n_450), .B2(n_454), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_154), .A2(n_202), .B1(n_454), .B2(n_795), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_155), .A2(n_369), .B1(n_1012), .B2(n_1015), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_157), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g422 ( .A(n_158), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_158), .B(n_215), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_158), .B(n_436), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_160), .B(n_289), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_161), .A2(n_210), .B1(n_536), .B2(n_537), .Y(n_583) );
AOI21xp33_ASAP7_75t_L g507 ( .A1(n_163), .A2(n_508), .B(n_509), .Y(n_507) );
AOI22xp5_ASAP7_75t_L g1038 ( .A1(n_164), .A2(n_168), .B1(n_1018), .B2(n_1020), .Y(n_1038) );
AOI221xp5_ASAP7_75t_L g479 ( .A1(n_165), .A2(n_337), .B1(n_480), .B2(n_483), .C(n_486), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_166), .A2(n_310), .B1(n_524), .B2(n_599), .Y(n_826) );
INVx1_ASAP7_75t_L g703 ( .A(n_167), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_170), .A2(n_339), .B1(n_630), .B2(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g936 ( .A(n_172), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_173), .A2(n_340), .B1(n_546), .B2(n_547), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_175), .B(n_631), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_176), .A2(n_208), .B1(n_654), .B2(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_177), .B(n_414), .Y(n_413) );
AO22x1_ASAP7_75t_L g929 ( .A1(n_178), .A2(n_317), .B1(n_543), .B2(n_544), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_180), .A2(n_324), .B1(n_520), .B2(n_522), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_182), .B(n_872), .Y(n_1256) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_183), .A2(n_259), .B1(n_443), .B2(n_518), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_184), .B(n_645), .Y(n_892) );
AOI21xp33_ASAP7_75t_L g962 ( .A1(n_185), .A2(n_705), .B(n_963), .Y(n_962) );
XOR2x2_ASAP7_75t_L g721 ( .A(n_186), .B(n_722), .Y(n_721) );
AOI21xp33_ASAP7_75t_SL g820 ( .A1(n_189), .A2(n_508), .B(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g730 ( .A(n_190), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_191), .A2(n_338), .B1(n_543), .B2(n_544), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_193), .A2(n_364), .B1(n_450), .B2(n_605), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_195), .A2(n_354), .B1(n_477), .B2(n_502), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g922 ( .A1(n_197), .A2(n_552), .B(n_923), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_198), .A2(n_269), .B1(n_1028), .B2(n_1059), .Y(n_1141) );
NAND2xp5_ASAP7_75t_SL g823 ( .A(n_199), .B(n_758), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_200), .B(n_701), .Y(n_947) );
AOI22xp33_ASAP7_75t_SL g1036 ( .A1(n_201), .A2(n_277), .B1(n_1022), .B2(n_1023), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_204), .A2(n_349), .B1(n_477), .B2(n_623), .Y(n_824) );
NAND2xp33_ASAP7_75t_L g677 ( .A(n_205), .B(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_206), .A2(n_280), .B1(n_718), .B2(n_768), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_211), .A2(n_238), .B1(n_857), .B2(n_858), .Y(n_856) );
AOI22xp33_ASAP7_75t_SL g577 ( .A1(n_212), .A2(n_236), .B1(n_565), .B2(n_567), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_213), .A2(n_279), .B1(n_614), .B2(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g405 ( .A(n_215), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g1029 ( .A1(n_216), .A2(n_217), .B1(n_1018), .B2(n_1020), .Y(n_1029) );
OAI22x1_ASAP7_75t_L g1242 ( .A1(n_216), .A2(n_1243), .B1(n_1249), .B2(n_1258), .Y(n_1242) );
NAND5xp2_ASAP7_75t_SL g1243 ( .A(n_216), .B(n_1244), .C(n_1245), .D(n_1247), .E(n_1248), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1266 ( .A1(n_216), .A2(n_1267), .B1(n_1288), .B2(n_1291), .Y(n_1266) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_219), .A2(n_268), .B1(n_765), .B2(n_766), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_220), .A2(n_346), .B1(n_450), .B2(n_526), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_222), .A2(n_246), .B1(n_543), .B2(n_544), .Y(n_542) );
INVx1_ASAP7_75t_L g822 ( .A(n_225), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_226), .A2(n_293), .B1(n_423), .B2(n_718), .Y(n_903) );
INVx1_ASAP7_75t_L g617 ( .A(n_227), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_228), .A2(n_266), .B1(n_518), .B2(n_598), .Y(n_1244) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_229), .A2(n_233), .B1(n_605), .B2(n_857), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_232), .A2(n_257), .B1(n_398), .B2(n_423), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_235), .A2(n_325), .B1(n_652), .B2(n_984), .Y(n_983) );
CKINVDCx14_ASAP7_75t_R g571 ( .A(n_239), .Y(n_571) );
XNOR2x2_ASAP7_75t_L g916 ( .A(n_240), .B(n_917), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_241), .B(n_630), .Y(n_711) );
INVx1_ASAP7_75t_L g734 ( .A(n_244), .Y(n_734) );
AOI21xp5_ASAP7_75t_SL g551 ( .A1(n_245), .A2(n_552), .B(n_553), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_247), .A2(n_303), .B1(n_558), .B2(n_561), .Y(n_804) );
INVx1_ASAP7_75t_L g612 ( .A(n_251), .Y(n_612) );
INVx1_ASAP7_75t_L g1140 ( .A(n_252), .Y(n_1140) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_255), .A2(n_284), .B1(n_450), .B2(n_454), .Y(n_449) );
INVx1_ASAP7_75t_L g973 ( .A(n_256), .Y(n_973) );
AOI221xp5_ASAP7_75t_L g755 ( .A1(n_260), .A2(n_370), .B1(n_756), .B2(n_757), .C(n_759), .Y(n_755) );
CKINVDCx5p33_ASAP7_75t_R g896 ( .A(n_261), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_262), .A2(n_328), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_263), .A2(n_295), .B1(n_611), .B2(n_1280), .Y(n_1279) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_264), .A2(n_368), .B1(n_428), .B2(n_601), .Y(n_843) );
INVx1_ASAP7_75t_L g875 ( .A(n_265), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_270), .A2(n_343), .B1(n_619), .B2(n_880), .Y(n_879) );
AOI22xp5_ASAP7_75t_SL g961 ( .A1(n_272), .A2(n_367), .B1(n_558), .B2(n_561), .Y(n_961) );
INVx1_ASAP7_75t_L g731 ( .A(n_273), .Y(n_731) );
INVx1_ASAP7_75t_L g966 ( .A(n_274), .Y(n_966) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_276), .Y(n_386) );
AND2x4_ASAP7_75t_L g1013 ( .A(n_276), .B(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_SL g531 ( .A(n_277), .Y(n_531) );
INVx1_ASAP7_75t_L g556 ( .A(n_283), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_287), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g737 ( .A(n_288), .Y(n_737) );
INVx1_ASAP7_75t_L g420 ( .A(n_289), .Y(n_420) );
INVxp67_ASAP7_75t_L g472 ( .A(n_289), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_290), .A2(n_499), .B1(n_527), .B2(n_528), .Y(n_498) );
INVxp67_ASAP7_75t_L g528 ( .A(n_290), .Y(n_528) );
OAI21x1_ASAP7_75t_L g791 ( .A1(n_292), .A2(n_792), .B(n_808), .Y(n_791) );
NAND4xp25_ASAP7_75t_L g808 ( .A(n_292), .B(n_793), .C(n_798), .D(n_805), .Y(n_808) );
INVxp67_ASAP7_75t_R g888 ( .A(n_296), .Y(n_888) );
INVx1_ASAP7_75t_L g914 ( .A(n_296), .Y(n_914) );
INVx2_ASAP7_75t_L g381 ( .A(n_298), .Y(n_381) );
INVx1_ASAP7_75t_L g563 ( .A(n_299), .Y(n_563) );
XOR2x2_ASAP7_75t_L g853 ( .A(n_300), .B(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g709 ( .A(n_304), .Y(n_709) );
INVx1_ASAP7_75t_L g1056 ( .A(n_305), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_307), .B(n_567), .Y(n_566) );
XNOR2x1_ASAP7_75t_L g691 ( .A(n_309), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g924 ( .A(n_312), .Y(n_924) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_319), .A2(n_348), .B1(n_546), .B2(n_547), .Y(n_684) );
INVx1_ASAP7_75t_L g625 ( .A(n_320), .Y(n_625) );
INVx1_ASAP7_75t_L g1254 ( .A(n_321), .Y(n_1254) );
INVx1_ASAP7_75t_L g964 ( .A(n_323), .Y(n_964) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_327), .A2(n_334), .B1(n_539), .B2(n_540), .Y(n_683) );
INVx1_ASAP7_75t_L g1060 ( .A(n_329), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_330), .A2(n_335), .B1(n_863), .B2(n_864), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_333), .B(n_489), .Y(n_578) );
AOI21xp33_ASAP7_75t_L g695 ( .A1(n_336), .A2(n_513), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g706 ( .A(n_345), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_347), .A2(n_356), .B1(n_518), .B2(n_991), .Y(n_990) );
INVx1_ASAP7_75t_L g550 ( .A(n_350), .Y(n_550) );
INVx1_ASAP7_75t_L g510 ( .A(n_362), .Y(n_510) );
AOI21xp33_ASAP7_75t_SL g688 ( .A1(n_365), .A2(n_552), .B(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_366), .A2(n_373), .B1(n_508), .B2(n_909), .Y(n_908) );
CKINVDCx20_ASAP7_75t_R g1277 ( .A(n_371), .Y(n_1277) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_387), .B(n_997), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
BUFx4_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
NAND3xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_382), .C(n_386), .Y(n_378) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_379), .B(n_1264), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_379), .B(n_1265), .Y(n_1290) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OA21x2_ASAP7_75t_L g1292 ( .A1(n_380), .A2(n_1019), .B(n_1293), .Y(n_1292) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_381), .B(n_1007), .Y(n_1006) );
AND3x4_ASAP7_75t_L g1018 ( .A(n_381), .B(n_1013), .C(n_1019), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1264 ( .A(n_382), .B(n_1265), .Y(n_1264) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_383), .A2(n_492), .B(n_493), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g1265 ( .A(n_386), .Y(n_1265) );
XNOR2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_784), .Y(n_387) );
XNOR2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_591), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_495), .B1(n_589), .B2(n_590), .Y(n_390) );
INVx1_ASAP7_75t_L g590 ( .A(n_391), .Y(n_590) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND4xp75_ASAP7_75t_L g395 ( .A(n_396), .B(n_441), .C(n_458), .D(n_479), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_427), .Y(n_396) );
BUFx2_ASAP7_75t_SL g666 ( .A(n_398), .Y(n_666) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx12f_ASAP7_75t_L g718 ( .A(n_399), .Y(n_718) );
BUFx6f_ASAP7_75t_L g868 ( .A(n_399), .Y(n_868) );
AND2x4_ASAP7_75t_L g399 ( .A(n_400), .B(n_411), .Y(n_399) );
AND2x4_ASAP7_75t_L g424 ( .A(n_400), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g451 ( .A(n_400), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g455 ( .A(n_400), .B(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g536 ( .A(n_400), .B(n_452), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_400), .B(n_456), .Y(n_537) );
AND2x4_ASAP7_75t_L g543 ( .A(n_400), .B(n_411), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_400), .B(n_445), .Y(n_544) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_409), .Y(n_400) );
AND2x2_ASAP7_75t_L g462 ( .A(n_401), .B(n_410), .Y(n_462) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g430 ( .A(n_402), .B(n_410), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_406), .Y(n_402) );
NAND2xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
INVx2_ASAP7_75t_L g408 ( .A(n_404), .Y(n_408) );
INVx3_ASAP7_75t_L g414 ( .A(n_404), .Y(n_414) );
NAND2xp33_ASAP7_75t_L g421 ( .A(n_404), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g440 ( .A(n_404), .Y(n_440) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_404), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_405), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_407), .A2(n_440), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g470 ( .A(n_410), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g429 ( .A(n_411), .B(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_L g433 ( .A(n_411), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g521 ( .A(n_411), .B(n_430), .Y(n_521) );
AND2x4_ASAP7_75t_L g546 ( .A(n_411), .B(n_430), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_411), .B(n_434), .Y(n_547) );
AND2x4_ASAP7_75t_L g411 ( .A(n_412), .B(n_416), .Y(n_411) );
OR2x2_ASAP7_75t_L g426 ( .A(n_412), .B(n_417), .Y(n_426) );
AND2x4_ASAP7_75t_L g452 ( .A(n_412), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g457 ( .A(n_412), .Y(n_457) );
AND2x2_ASAP7_75t_L g466 ( .A(n_412), .B(n_467), .Y(n_466) );
AND2x4_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_414), .B(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g436 ( .A(n_414), .Y(n_436) );
NAND3xp33_ASAP7_75t_L g493 ( .A(n_415), .B(n_435), .C(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g453 ( .A(n_418), .Y(n_453) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
BUFx3_ASAP7_75t_L g658 ( .A(n_423), .Y(n_658) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_424), .Y(n_524) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_424), .Y(n_598) );
BUFx6f_ASAP7_75t_L g768 ( .A(n_424), .Y(n_768) );
AND2x4_ASAP7_75t_L g448 ( .A(n_425), .B(n_434), .Y(n_448) );
AND2x4_ASAP7_75t_L g539 ( .A(n_425), .B(n_430), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_425), .B(n_434), .Y(n_540) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g445 ( .A(n_426), .Y(n_445) );
BUFx3_ASAP7_75t_L g661 ( .A(n_428), .Y(n_661) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx8_ASAP7_75t_L g863 ( .A(n_429), .Y(n_863) );
AND2x4_ASAP7_75t_L g444 ( .A(n_430), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g476 ( .A(n_430), .B(n_452), .Y(n_476) );
AND2x2_ASAP7_75t_L g485 ( .A(n_430), .B(n_456), .Y(n_485) );
AND2x2_ASAP7_75t_L g506 ( .A(n_430), .B(n_456), .Y(n_506) );
AND2x4_ASAP7_75t_L g565 ( .A(n_430), .B(n_452), .Y(n_565) );
INVx4_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g522 ( .A(n_432), .Y(n_522) );
INVx4_ASAP7_75t_L g601 ( .A(n_432), .Y(n_601) );
INVx2_ASAP7_75t_L g668 ( .A(n_432), .Y(n_668) );
INVx2_ASAP7_75t_SL g720 ( .A(n_432), .Y(n_720) );
INVx1_ASAP7_75t_L g777 ( .A(n_432), .Y(n_777) );
INVx1_ASAP7_75t_L g869 ( .A(n_432), .Y(n_869) );
INVx2_ASAP7_75t_L g905 ( .A(n_432), .Y(n_905) );
INVx4_ASAP7_75t_L g1246 ( .A(n_432), .Y(n_1246) );
INVx8_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g478 ( .A(n_434), .B(n_456), .Y(n_478) );
AND2x4_ASAP7_75t_L g561 ( .A(n_434), .B(n_456), .Y(n_561) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_439), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_449), .Y(n_441) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx12f_ASAP7_75t_L g517 ( .A(n_444), .Y(n_517) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_444), .Y(n_603) );
BUFx3_ASAP7_75t_L g864 ( .A(n_444), .Y(n_864) );
BUFx6f_ASAP7_75t_L g991 ( .A(n_444), .Y(n_991) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx5_ASAP7_75t_L g599 ( .A(n_447), .Y(n_599) );
INVx3_ASAP7_75t_L g797 ( .A(n_447), .Y(n_797) );
INVx1_ASAP7_75t_L g866 ( .A(n_447), .Y(n_866) );
INVx2_ASAP7_75t_L g1285 ( .A(n_447), .Y(n_1285) );
INVx6_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx12f_ASAP7_75t_L g518 ( .A(n_448), .Y(n_518) );
BUFx12f_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g771 ( .A(n_451), .Y(n_771) );
BUFx6f_ASAP7_75t_L g857 ( .A(n_451), .Y(n_857) );
AND2x4_ASAP7_75t_L g461 ( .A(n_452), .B(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g558 ( .A(n_452), .B(n_462), .Y(n_558) );
AND2x4_ASAP7_75t_L g456 ( .A(n_453), .B(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_455), .Y(n_526) );
BUFx5_ASAP7_75t_L g605 ( .A(n_455), .Y(n_605) );
INVx1_ASAP7_75t_L g861 ( .A(n_455), .Y(n_861) );
AND2x4_ASAP7_75t_L g482 ( .A(n_456), .B(n_462), .Y(n_482) );
AND2x2_ASAP7_75t_L g552 ( .A(n_456), .B(n_462), .Y(n_552) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_473), .Y(n_458) );
BUFx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx3_ASAP7_75t_L g513 ( .A(n_461), .Y(n_513) );
INVx1_ASAP7_75t_L g620 ( .A(n_461), .Y(n_620) );
BUFx6f_ASAP7_75t_L g1274 ( .A(n_461), .Y(n_1274) );
INVx4_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g648 ( .A(n_464), .Y(n_648) );
INVx3_ASAP7_75t_L g756 ( .A(n_464), .Y(n_756) );
INVx2_ASAP7_75t_L g911 ( .A(n_464), .Y(n_911) );
INVx2_ASAP7_75t_L g982 ( .A(n_464), .Y(n_982) );
INVx5_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g514 ( .A(n_465), .Y(n_514) );
BUFx4f_ASAP7_75t_L g630 ( .A(n_465), .Y(n_630) );
BUFx2_ASAP7_75t_L g819 ( .A(n_465), .Y(n_819) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_470), .Y(n_465) );
AND2x4_ASAP7_75t_L g567 ( .A(n_466), .B(n_470), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g492 ( .A(n_468), .Y(n_492) );
INVx1_ASAP7_75t_L g710 ( .A(n_474), .Y(n_710) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx6f_ASAP7_75t_L g881 ( .A(n_475), .Y(n_881) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx3_ASAP7_75t_L g502 ( .A(n_476), .Y(n_502) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_476), .Y(n_623) );
INVx3_ASAP7_75t_L g707 ( .A(n_477), .Y(n_707) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx3_ASAP7_75t_L g615 ( .A(n_478), .Y(n_615) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_478), .Y(n_652) );
INVx2_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_SL g984 ( .A(n_481), .Y(n_984) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_482), .Y(n_508) );
BUFx3_ASAP7_75t_L g611 ( .A(n_482), .Y(n_611) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_482), .Y(n_705) );
INVx2_ASAP7_75t_L g849 ( .A(n_482), .Y(n_849) );
BUFx8_ASAP7_75t_SL g878 ( .A(n_482), .Y(n_878) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI21xp33_ASAP7_75t_L g549 ( .A1(n_484), .A2(n_550), .B(n_551), .Y(n_549) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_485), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx2_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_SL g489 ( .A(n_490), .Y(n_489) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_490), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_490), .B(n_554), .Y(n_553) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_490), .Y(n_632) );
INVx2_ASAP7_75t_L g699 ( .A(n_490), .Y(n_699) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g743 ( .A(n_491), .Y(n_743) );
INVx2_ASAP7_75t_L g589 ( .A(n_495), .Y(n_589) );
OAI22x1_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B1(n_568), .B2(n_587), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
XOR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_529), .Y(n_497) );
INVx1_ASAP7_75t_L g527 ( .A(n_499), .Y(n_527) );
NOR2xp67_ASAP7_75t_L g499 ( .A(n_500), .B(n_515), .Y(n_499) );
NAND4xp25_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .C(n_507), .D(n_512), .Y(n_500) );
BUFx2_ASAP7_75t_L g655 ( .A(n_502), .Y(n_655) );
INVx2_ASAP7_75t_L g732 ( .A(n_502), .Y(n_732) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g701 ( .A(n_505), .Y(n_701) );
INVx2_ASAP7_75t_L g739 ( .A(n_505), .Y(n_739) );
INVx2_ASAP7_75t_L g1275 ( .A(n_505), .Y(n_1275) );
INVx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g628 ( .A(n_506), .Y(n_628) );
BUFx3_ASAP7_75t_L g851 ( .A(n_506), .Y(n_851) );
BUFx3_ASAP7_75t_L g650 ( .A(n_508), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
BUFx2_ASAP7_75t_L g654 ( .A(n_513), .Y(n_654) );
NAND4xp25_ASAP7_75t_L g515 ( .A(n_516), .B(n_519), .C(n_523), .D(n_525), .Y(n_515) );
BUFx3_ASAP7_75t_L g662 ( .A(n_517), .Y(n_662) );
BUFx3_ASAP7_75t_L g659 ( .A(n_518), .Y(n_659) );
BUFx4f_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx6f_ASAP7_75t_L g775 ( .A(n_521), .Y(n_775) );
BUFx2_ASAP7_75t_SL g772 ( .A(n_526), .Y(n_772) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g635 ( .A(n_530), .Y(n_635) );
XNOR2x1_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
XNOR2xp5_ASAP7_75t_L g636 ( .A(n_531), .B(n_532), .Y(n_636) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_548), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_541), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_545), .Y(n_541) );
NOR3xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_555), .C(n_562), .Y(n_548) );
OAI22xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_559), .B2(n_560), .Y(n_555) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVxp67_ASAP7_75t_L g680 ( .A(n_560), .Y(n_680) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OAI21xp5_ASAP7_75t_SL g562 ( .A1(n_563), .A2(n_564), .B(n_566), .Y(n_562) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx4_ASAP7_75t_L g874 ( .A(n_567), .Y(n_874) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g588 ( .A(n_570), .Y(n_588) );
OAI21x1_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_572), .B(n_584), .Y(n_570) );
NAND3xp33_ASAP7_75t_SL g584 ( .A(n_571), .B(n_585), .C(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_579), .Y(n_573) );
INVx1_ASAP7_75t_L g586 ( .A(n_574), .Y(n_586) );
NAND4xp25_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .C(n_577), .D(n_578), .Y(n_574) );
INVxp67_ASAP7_75t_L g585 ( .A(n_579), .Y(n_585) );
NAND4xp25_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .C(n_582), .D(n_583), .Y(n_579) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B1(n_670), .B2(n_783), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI22x1_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_638), .B1(n_639), .B2(n_669), .Y(n_593) );
INVx2_ASAP7_75t_L g669 ( .A(n_594), .Y(n_669) );
AO22x2_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_635), .B1(n_636), .B2(n_637), .Y(n_594) );
INVx2_ASAP7_75t_L g637 ( .A(n_595), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_596), .B(n_607), .Y(n_634) );
AND4x1_ASAP7_75t_L g596 ( .A(n_597), .B(n_600), .C(n_602), .D(n_604), .Y(n_596) );
BUFx3_ASAP7_75t_L g664 ( .A(n_605), .Y(n_664) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_633), .Y(n_606) );
NOR3xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_616), .C(n_624), .Y(n_607) );
OAI22xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B1(n_612), .B2(n_613), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_610), .A2(n_615), .B1(n_734), .B2(n_735), .Y(n_733) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx3_ASAP7_75t_L g909 ( .A(n_615), .Y(n_909) );
INVx2_ASAP7_75t_L g1280 ( .A(n_615), .Y(n_1280) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B1(n_621), .B2(n_622), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_618), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_729) );
INVx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g894 ( .A(n_620), .Y(n_894) );
INVx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx3_ASAP7_75t_L g752 ( .A(n_623), .Y(n_752) );
OAI21xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B(n_629), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_628), .Y(n_646) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_632), .B(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_632), .B(n_822), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g1276 ( .A(n_632), .B(n_1277), .Y(n_1276) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_633), .A2(n_1058), .B1(n_1060), .B2(n_1061), .Y(n_1057) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2x1_ASAP7_75t_L g640 ( .A(n_641), .B(n_656), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_649), .C(n_653), .Y(n_641) );
INVx2_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g758 ( .A(n_646), .Y(n_758) );
INVx2_ASAP7_75t_L g872 ( .A(n_646), .Y(n_872) );
BUFx3_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND4xp25_ASAP7_75t_SL g656 ( .A(n_657), .B(n_660), .C(n_663), .D(n_665), .Y(n_656) );
BUFx2_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g783 ( .A(n_670), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_746), .B1(n_781), .B2(n_782), .Y(n_670) );
INVx1_ASAP7_75t_L g781 ( .A(n_671), .Y(n_781) );
AO22x2_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_721), .B1(n_744), .B2(n_745), .Y(n_671) );
INVx1_ASAP7_75t_L g745 ( .A(n_672), .Y(n_745) );
XNOR2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_691), .Y(n_672) );
XNOR2x1_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
NOR2x1_ASAP7_75t_L g675 ( .A(n_676), .B(n_682), .Y(n_675) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .C(n_681), .Y(n_676) );
NAND4xp25_ASAP7_75t_SL g682 ( .A(n_683), .B(n_684), .C(n_685), .D(n_688), .Y(n_682) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_712), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_702), .C(n_708), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_700), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g895 ( .A(n_698), .B(n_896), .Y(n_895) );
NOR2xp33_ASAP7_75t_L g978 ( .A(n_698), .B(n_979), .Y(n_978) );
INVx3_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_706), .B2(n_707), .Y(n_702) );
INVx1_ASAP7_75t_L g754 ( .A(n_704), .Y(n_754) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OAI21xp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_710), .B(n_711), .Y(n_708) );
NOR2xp33_ASAP7_75t_SL g712 ( .A(n_713), .B(n_716), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
BUFx6f_ASAP7_75t_L g765 ( .A(n_718), .Y(n_765) );
INVx1_ASAP7_75t_L g744 ( .A(n_721), .Y(n_744) );
AND2x4_ASAP7_75t_L g722 ( .A(n_723), .B(n_728), .Y(n_722) );
AND4x1_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .C(n_726), .D(n_727), .Y(n_723) );
NOR3xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_733), .C(n_736), .Y(n_728) );
OAI21xp33_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .B(n_740), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx4_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g923 ( .A(n_742), .B(n_924), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g1253 ( .A(n_742), .B(n_1254), .Y(n_1253) );
INVx4_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx3_ASAP7_75t_L g761 ( .A(n_743), .Y(n_761) );
BUFx3_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g782 ( .A(n_747), .Y(n_782) );
OR2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_762), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_749), .B(n_762), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_755), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_751), .B(n_753), .Y(n_750) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g800 ( .A(n_761), .B(n_801), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g949 ( .A(n_761), .B(n_950), .Y(n_949) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_761), .B(n_964), .Y(n_963) );
NAND2x1p5_ASAP7_75t_L g762 ( .A(n_763), .B(n_773), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_769), .Y(n_763) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g795 ( .A(n_771), .Y(n_795) );
INVx2_ASAP7_75t_L g943 ( .A(n_771), .Y(n_943) );
AND2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_778), .Y(n_773) );
BUFx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
XNOR2x1_ASAP7_75t_L g784 ( .A(n_785), .B(n_882), .Y(n_784) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
XNOR2x1_ASAP7_75t_SL g786 ( .A(n_787), .B(n_809), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
AND3x1_ASAP7_75t_L g792 ( .A(n_793), .B(n_798), .C(n_805), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_796), .Y(n_793) );
AND2x2_ASAP7_75t_L g798 ( .A(n_799), .B(n_802), .Y(n_798) );
AND2x2_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
XOR2x1_ASAP7_75t_L g809 ( .A(n_810), .B(n_853), .Y(n_809) );
XNOR2x1_ASAP7_75t_L g810 ( .A(n_811), .B(n_836), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
OAI21x1_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_815), .B(n_830), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_813), .B(n_824), .Y(n_833) );
CKINVDCx5p33_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
NOR2xp67_ASAP7_75t_L g815 ( .A(n_816), .B(n_825), .Y(n_815) );
NAND3xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_823), .C(n_824), .Y(n_816) );
INVx1_ASAP7_75t_L g834 ( .A(n_817), .Y(n_834) );
AND2x2_ASAP7_75t_L g817 ( .A(n_818), .B(n_820), .Y(n_817) );
INVxp67_ASAP7_75t_L g832 ( .A(n_823), .Y(n_832) );
INVx1_ASAP7_75t_L g835 ( .A(n_825), .Y(n_835) );
NAND4xp25_ASAP7_75t_L g825 ( .A(n_826), .B(n_827), .C(n_828), .D(n_829), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_835), .Y(n_830) );
NOR3xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .C(n_834), .Y(n_831) );
INVx2_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
XOR2x2_ASAP7_75t_L g837 ( .A(n_838), .B(n_852), .Y(n_837) );
NOR2x1_ASAP7_75t_L g838 ( .A(n_839), .B(n_844), .Y(n_838) );
NAND4xp25_ASAP7_75t_L g839 ( .A(n_840), .B(n_841), .C(n_842), .D(n_843), .Y(n_839) );
NAND4xp25_ASAP7_75t_L g844 ( .A(n_845), .B(n_846), .C(n_847), .D(n_850), .Y(n_844) );
INVx3_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NOR2x1_ASAP7_75t_L g854 ( .A(n_855), .B(n_870), .Y(n_854) );
NAND4xp25_ASAP7_75t_L g855 ( .A(n_856), .B(n_862), .C(n_865), .D(n_867), .Y(n_855) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
NAND3xp33_ASAP7_75t_L g870 ( .A(n_871), .B(n_877), .C(n_879), .Y(n_870) );
OAI21xp5_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_875), .B(n_876), .Y(n_873) );
INVx2_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
OA22x2_ASAP7_75t_L g882 ( .A1(n_883), .A2(n_931), .B1(n_932), .B2(n_996), .Y(n_882) );
INVx1_ASAP7_75t_L g996 ( .A(n_883), .Y(n_996) );
BUFx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
OA22x2_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_887), .B1(n_915), .B2(n_916), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
OAI21x1_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .B(n_912), .Y(n_887) );
NOR4xp75_ASAP7_75t_L g889 ( .A(n_890), .B(n_897), .C(n_901), .D(n_906), .Y(n_889) );
INVx3_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
NAND4xp75_ASAP7_75t_L g912 ( .A(n_891), .B(n_898), .C(n_902), .D(n_913), .Y(n_912) );
AND2x2_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .Y(n_891) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_899), .B(n_900), .Y(n_898) );
INVx2_ASAP7_75t_SL g901 ( .A(n_902), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
AND2x2_ASAP7_75t_L g913 ( .A(n_907), .B(n_914), .Y(n_913) );
AND2x2_ASAP7_75t_L g907 ( .A(n_908), .B(n_910), .Y(n_907) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
XNOR2x1_ASAP7_75t_L g951 ( .A(n_916), .B(n_952), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_918), .B(n_925), .Y(n_917) );
AND4x1_ASAP7_75t_L g918 ( .A(n_919), .B(n_920), .C(n_921), .D(n_922), .Y(n_918) );
NOR4xp25_ASAP7_75t_L g925 ( .A(n_926), .B(n_928), .C(n_929), .D(n_930), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx2_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
OAI22x1_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_969), .B1(n_992), .B2(n_995), .Y(n_932) );
INVx4_ASAP7_75t_L g995 ( .A(n_933), .Y(n_995) );
AO22x2_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_951), .B1(n_967), .B2(n_968), .Y(n_933) );
INVxp67_ASAP7_75t_SL g967 ( .A(n_934), .Y(n_967) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
XNOR2x1_ASAP7_75t_L g935 ( .A(n_936), .B(n_937), .Y(n_935) );
NOR2x1_ASAP7_75t_L g937 ( .A(n_938), .B(n_944), .Y(n_937) );
NAND4xp25_ASAP7_75t_L g938 ( .A(n_939), .B(n_940), .C(n_941), .D(n_942), .Y(n_938) );
NAND4xp25_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .C(n_947), .D(n_948), .Y(n_944) );
INVx2_ASAP7_75t_L g968 ( .A(n_951), .Y(n_968) );
XOR2x2_ASAP7_75t_L g952 ( .A(n_953), .B(n_966), .Y(n_952) );
NOR2x1_ASAP7_75t_L g953 ( .A(n_954), .B(n_959), .Y(n_953) );
NAND4xp25_ASAP7_75t_L g954 ( .A(n_955), .B(n_956), .C(n_957), .D(n_958), .Y(n_954) );
NAND4xp25_ASAP7_75t_L g959 ( .A(n_960), .B(n_961), .C(n_962), .D(n_965), .Y(n_959) );
INVxp67_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx2_ASAP7_75t_SL g971 ( .A(n_972), .Y(n_971) );
INVx2_ASAP7_75t_L g994 ( .A(n_972), .Y(n_994) );
XNOR2x1_ASAP7_75t_L g972 ( .A(n_973), .B(n_974), .Y(n_972) );
NOR4xp75_ASAP7_75t_L g974 ( .A(n_975), .B(n_980), .C(n_985), .D(n_988), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_976), .B(n_977), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_981), .B(n_983), .Y(n_980) );
NAND2xp5_ASAP7_75t_SL g985 ( .A(n_986), .B(n_987), .Y(n_985) );
NAND2xp5_ASAP7_75t_SL g988 ( .A(n_989), .B(n_990), .Y(n_988) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
BUFx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
OAI221xp5_ASAP7_75t_L g997 ( .A1(n_998), .A2(n_1238), .B1(n_1239), .B2(n_1262), .C(n_1266), .Y(n_997) );
AOI211xp5_ASAP7_75t_L g998 ( .A1(n_999), .A2(n_1137), .B(n_1142), .C(n_1210), .Y(n_998) );
NAND4xp25_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1082), .C(n_1105), .D(n_1126), .Y(n_999) );
AOI211xp5_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1024), .B(n_1044), .C(n_1069), .Y(n_1000) );
AOI21xp33_ASAP7_75t_L g1179 ( .A1(n_1001), .A2(n_1180), .B(n_1181), .Y(n_1179) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
NOR2xp33_ASAP7_75t_L g1101 ( .A(n_1002), .B(n_1081), .Y(n_1101) );
OR2x2_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1016), .Y(n_1002) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1003), .Y(n_1064) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1003), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1011), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1008), .Y(n_1005) );
AND2x4_ASAP7_75t_L g1012 ( .A(n_1006), .B(n_1013), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_1006), .B(n_1008), .Y(n_1022) );
AND2x4_ASAP7_75t_L g1059 ( .A(n_1006), .B(n_1008), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_1008), .B(n_1010), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_1008), .B(n_1010), .Y(n_1023) );
AND2x4_ASAP7_75t_L g1028 ( .A(n_1008), .B(n_1010), .Y(n_1028) );
AND2x4_ASAP7_75t_L g1015 ( .A(n_1010), .B(n_1013), .Y(n_1015) );
AND2x4_ASAP7_75t_L g1020 ( .A(n_1010), .B(n_1013), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_1010), .B(n_1013), .Y(n_1055) );
INVx3_ASAP7_75t_L g1053 ( .A(n_1012), .Y(n_1053) );
CKINVDCx5p33_ASAP7_75t_R g1293 ( .A(n_1013), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1016), .B(n_1063), .Y(n_1062) );
OR2x2_ASAP7_75t_L g1065 ( .A(n_1016), .B(n_1051), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1016), .B(n_1081), .Y(n_1080) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1016), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1016), .B(n_1064), .Y(n_1104) );
OR2x2_ASAP7_75t_L g1109 ( .A(n_1016), .B(n_1081), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1016), .B(n_1051), .Y(n_1122) );
OR2x2_ASAP7_75t_L g1135 ( .A(n_1016), .B(n_1064), .Y(n_1135) );
HB1xp67_ASAP7_75t_L g1157 ( .A(n_1016), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_1017), .B(n_1021), .Y(n_1016) );
NOR2x1_ASAP7_75t_R g1024 ( .A(n_1025), .B(n_1030), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1025), .B(n_1034), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_1025), .B(n_1068), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1025), .B(n_1075), .Y(n_1099) );
NOR2xp33_ASAP7_75t_L g1114 ( .A(n_1025), .B(n_1115), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1025), .B(n_1037), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1025), .B(n_1113), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1025), .B(n_1033), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1025), .B(n_1180), .Y(n_1215) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_SL g1078 ( .A(n_1026), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1026), .B(n_1113), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1026), .B(n_1148), .Y(n_1147) );
OR2x2_ASAP7_75t_L g1162 ( .A(n_1026), .B(n_1087), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1026), .B(n_1034), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1026), .B(n_1180), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1029), .Y(n_1026) );
INVx2_ASAP7_75t_L g1061 ( .A(n_1028), .Y(n_1061) );
NAND2xp5_ASAP7_75t_SL g1030 ( .A(n_1031), .B(n_1040), .Y(n_1030) );
INVx3_ASAP7_75t_SL g1031 ( .A(n_1032), .Y(n_1031) );
NOR2x1_ASAP7_75t_L g1180 ( .A(n_1032), .B(n_1040), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1037), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1033), .B(n_1037), .Y(n_1075) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1034), .B(n_1037), .Y(n_1068) );
OR2x2_ASAP7_75t_L g1087 ( .A(n_1034), .B(n_1037), .Y(n_1087) );
AOI221xp5_ASAP7_75t_L g1200 ( .A1(n_1034), .A2(n_1049), .B1(n_1130), .B2(n_1201), .C(n_1203), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .Y(n_1034) );
O2A1O1Ixp33_ASAP7_75t_L g1069 ( .A1(n_1037), .A2(n_1070), .B(n_1073), .C(n_1079), .Y(n_1069) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1037), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1037), .B(n_1077), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1039), .Y(n_1037) );
NAND2xp5_ASAP7_75t_SL g1045 ( .A(n_1040), .B(n_1046), .Y(n_1045) );
NOR2xp33_ASAP7_75t_L g1071 ( .A(n_1040), .B(n_1072), .Y(n_1071) );
INVx2_ASAP7_75t_L g1084 ( .A(n_1040), .Y(n_1084) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1040), .Y(n_1118) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1040), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1040), .B(n_1075), .Y(n_1148) );
BUFx6f_ASAP7_75t_L g1160 ( .A(n_1040), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1040), .B(n_1184), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1040), .B(n_1050), .Y(n_1195) );
INVx4_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
OR2x2_ASAP7_75t_L g1076 ( .A(n_1041), .B(n_1077), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1041), .B(n_1081), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1041), .B(n_1051), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1043), .Y(n_1041) );
OAI22xp5_ASAP7_75t_L g1044 ( .A1(n_1045), .A2(n_1048), .B1(n_1065), .B2(n_1066), .Y(n_1044) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1062), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_1049), .B(n_1093), .Y(n_1092) );
INVx2_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1050), .B(n_1107), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1223 ( .A(n_1050), .B(n_1083), .Y(n_1223) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1051), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1051), .B(n_1104), .Y(n_1103) );
OR2x2_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1057), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_1053), .A2(n_1054), .B1(n_1055), .B2(n_1056), .Y(n_1052) );
OAI221xp5_ASAP7_75t_L g1138 ( .A1(n_1053), .A2(n_1055), .B1(n_1139), .B2(n_1140), .C(n_1141), .Y(n_1138) );
BUFx2_ASAP7_75t_L g1238 ( .A(n_1055), .Y(n_1238) );
INVx3_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
AOI221xp5_ASAP7_75t_L g1165 ( .A1(n_1062), .A2(n_1166), .B1(n_1168), .B2(n_1171), .C(n_1178), .Y(n_1165) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1063), .Y(n_1093) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
NOR2xp33_ASAP7_75t_L g1117 ( .A(n_1065), .B(n_1118), .Y(n_1117) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1065), .Y(n_1170) );
NOR2xp33_ASAP7_75t_L g1186 ( .A(n_1065), .B(n_1072), .Y(n_1186) );
OAI22xp5_ASAP7_75t_L g1228 ( .A1(n_1065), .A2(n_1229), .B1(n_1230), .B2(n_1232), .Y(n_1228) );
OAI221xp5_ASAP7_75t_L g1178 ( .A1(n_1066), .A2(n_1137), .B1(n_1179), .B2(n_1185), .C(n_1187), .Y(n_1178) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1067), .B(n_1080), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1068), .B(n_1090), .Y(n_1089) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_1068), .B(n_1103), .Y(n_1102) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1068), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1068), .B(n_1077), .Y(n_1125) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx2_ASAP7_75t_L g1107 ( .A(n_1072), .Y(n_1107) );
BUFx3_ASAP7_75t_L g1169 ( .A(n_1072), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1072), .B(n_1081), .Y(n_1198) );
OR2x2_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1076), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1075), .B(n_1077), .Y(n_1130) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1076), .Y(n_1090) );
AND2x4_ASAP7_75t_L g1085 ( .A(n_1077), .B(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
INVx2_ASAP7_75t_L g1128 ( .A(n_1081), .Y(n_1128) );
AOI21xp33_ASAP7_75t_SL g1214 ( .A1(n_1081), .A2(n_1215), .B(n_1216), .Y(n_1214) );
O2A1O1Ixp33_ASAP7_75t_L g1082 ( .A1(n_1083), .A2(n_1088), .B(n_1091), .C(n_1094), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1085), .Y(n_1083) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1084), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1084), .B(n_1112), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_1084), .B(n_1099), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1084), .B(n_1177), .Y(n_1176) );
NOR2xp33_ASAP7_75t_L g1236 ( .A(n_1084), .B(n_1087), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_1085), .B(n_1096), .Y(n_1095) );
INVx2_ASAP7_75t_SL g1174 ( .A(n_1085), .Y(n_1174) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_1087), .B(n_1116), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_1088), .A2(n_1104), .B1(n_1191), .B2(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
NOR2xp33_ASAP7_75t_L g1206 ( .A(n_1093), .B(n_1154), .Y(n_1206) );
OAI221xp5_ASAP7_75t_L g1094 ( .A1(n_1095), .A2(n_1097), .B1(n_1098), .B2(n_1100), .C(n_1102), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_1096), .B(n_1125), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1097), .B(n_1202), .Y(n_1201) );
CKINVDCx14_ASAP7_75t_R g1227 ( .A(n_1097), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1097), .B(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1103), .Y(n_1237) );
AOI211xp5_ASAP7_75t_L g1126 ( .A1(n_1104), .A2(n_1127), .B(n_1131), .C(n_1134), .Y(n_1126) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1104), .Y(n_1182) );
AOI221xp5_ASAP7_75t_L g1105 ( .A1(n_1106), .A2(n_1110), .B1(n_1114), .B2(n_1117), .C(n_1119), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1108), .Y(n_1106) );
NOR2xp33_ASAP7_75t_L g1196 ( .A(n_1107), .B(n_1137), .Y(n_1196) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1107), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1107), .B(n_1138), .Y(n_1217) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
NOR2xp33_ASAP7_75t_L g1221 ( .A(n_1109), .B(n_1118), .Y(n_1221) );
INVxp67_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1113), .B(n_1160), .Y(n_1167) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1117), .Y(n_1207) );
AOI21xp5_ASAP7_75t_L g1119 ( .A1(n_1120), .A2(n_1123), .B(n_1124), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1122), .Y(n_1120) );
NAND2xp67_ASAP7_75t_L g1129 ( .A(n_1121), .B(n_1130), .Y(n_1129) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1122), .Y(n_1161) );
AOI221xp5_ASAP7_75t_SL g1197 ( .A1(n_1122), .A2(n_1146), .B1(n_1176), .B2(n_1198), .C(n_1199), .Y(n_1197) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1123), .Y(n_1209) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
NOR2xp33_ASAP7_75t_L g1229 ( .A(n_1125), .B(n_1177), .Y(n_1229) );
NOR2xp67_ASAP7_75t_SL g1127 ( .A(n_1128), .B(n_1129), .Y(n_1127) );
INVx2_ASAP7_75t_L g1132 ( .A(n_1128), .Y(n_1132) );
NOR2xp33_ASAP7_75t_L g1173 ( .A(n_1128), .B(n_1174), .Y(n_1173) );
NAND2xp5_ASAP7_75t_L g1175 ( .A(n_1128), .B(n_1176), .Y(n_1175) );
AOI221xp5_ASAP7_75t_L g1218 ( .A1(n_1128), .A2(n_1194), .B1(n_1219), .B2(n_1221), .C(n_1222), .Y(n_1218) );
NOR2xp33_ASAP7_75t_L g1225 ( .A(n_1129), .B(n_1132), .Y(n_1225) );
NOR2xp33_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1133), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1132), .B(n_1213), .Y(n_1212) );
AOI21xp33_ASAP7_75t_L g1234 ( .A1(n_1133), .A2(n_1235), .B(n_1237), .Y(n_1234) );
NOR2xp33_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1136), .Y(n_1134) );
OAI211xp5_ASAP7_75t_L g1166 ( .A1(n_1137), .A2(n_1147), .B(n_1162), .C(n_1167), .Y(n_1166) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1137), .Y(n_1231) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
HB1xp67_ASAP7_75t_L g1144 ( .A(n_1138), .Y(n_1144) );
OAI211xp5_ASAP7_75t_L g1142 ( .A1(n_1143), .A2(n_1145), .B(n_1165), .C(n_1197), .Y(n_1142) );
INVx2_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
O2A1O1Ixp33_ASAP7_75t_L g1145 ( .A1(n_1146), .A2(n_1149), .B(n_1155), .C(n_1158), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
NAND3xp33_ASAP7_75t_L g1171 ( .A(n_1147), .B(n_1172), .C(n_1175), .Y(n_1171) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1148), .Y(n_1220) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1153), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
NOR2xp33_ASAP7_75t_L g1188 ( .A(n_1152), .B(n_1189), .Y(n_1188) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
A2O1A1Ixp33_ASAP7_75t_L g1158 ( .A1(n_1159), .A2(n_1161), .B(n_1162), .C(n_1163), .Y(n_1158) );
AOI221xp5_ASAP7_75t_L g1224 ( .A1(n_1159), .A2(n_1225), .B1(n_1226), .B2(n_1228), .C(n_1234), .Y(n_1224) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1162), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1162), .B(n_1220), .Y(n_1219) );
CKINVDCx5p33_ASAP7_75t_R g1163 ( .A(n_1164), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1170), .Y(n_1168) );
OAI321xp33_ASAP7_75t_L g1210 ( .A1(n_1170), .A2(n_1211), .A3(n_1214), .B1(n_1217), .B2(n_1218), .C(n_1224), .Y(n_1210) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
NOR2xp33_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1183), .Y(n_1181) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
OAI21xp33_ASAP7_75t_L g1187 ( .A1(n_1188), .A2(n_1191), .B(n_1196), .Y(n_1187) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1190), .Y(n_1189) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1195), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1196), .Y(n_1204) );
OAI221xp5_ASAP7_75t_L g1199 ( .A1(n_1200), .A2(n_1204), .B1(n_1205), .B2(n_1207), .C(n_1208), .Y(n_1199) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1203), .Y(n_1213) );
INVxp67_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
INVxp67_ASAP7_75t_SL g1211 ( .A(n_1212), .Y(n_1211) );
INVxp67_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
CKINVDCx14_ASAP7_75t_R g1226 ( .A(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
BUFx3_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
BUFx3_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
NAND4xp25_ASAP7_75t_L g1259 ( .A(n_1244), .B(n_1245), .C(n_1248), .D(n_1256), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1247), .B(n_1257), .Y(n_1261) );
NAND3xp33_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1256), .C(n_1257), .Y(n_1249) );
INVxp67_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1260 ( .A(n_1251), .B(n_1261), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1252), .B(n_1255), .Y(n_1251) );
NOR2x1_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1260), .Y(n_1258) );
CKINVDCx16_ASAP7_75t_R g1262 ( .A(n_1263), .Y(n_1262) );
INVxp33_ASAP7_75t_SL g1267 ( .A(n_1268), .Y(n_1267) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
INVxp33_ASAP7_75t_SL g1270 ( .A(n_1271), .Y(n_1270) );
OR2x2_ASAP7_75t_L g1271 ( .A(n_1272), .B(n_1281), .Y(n_1271) );
NAND3xp33_ASAP7_75t_L g1272 ( .A(n_1273), .B(n_1278), .C(n_1279), .Y(n_1272) );
NAND4xp25_ASAP7_75t_SL g1281 ( .A(n_1282), .B(n_1283), .C(n_1284), .D(n_1286), .Y(n_1281) );
HB1xp67_ASAP7_75t_SL g1288 ( .A(n_1289), .Y(n_1288) );
BUFx2_ASAP7_75t_SL g1289 ( .A(n_1290), .Y(n_1289) );
BUFx2_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
endmodule