module fake_jpeg_18449_n_74 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_64;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_71;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_67;
wire n_56;
wire n_43;
wire n_37;
wire n_29;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_10),
.A2(n_11),
.B(n_5),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_7),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_2),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_44),
.B(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_24),
.A2(n_37),
.B(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_20),
.B(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_22),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_30),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_31),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_25),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_54),
.A2(n_47),
.B1(n_53),
.B2(n_51),
.Y(n_59)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_61),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_60),
.B1(n_59),
.B2(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_49),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_56),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_64),
.B(n_55),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_48),
.B(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

OAI311xp33_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_62),
.A3(n_70),
.B1(n_40),
.C1(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_50),
.Y(n_74)
);


endmodule