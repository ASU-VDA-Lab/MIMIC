module fake_jpeg_3049_n_580 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_580);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_580;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_17),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_61),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_62),
.B(n_69),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_63),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_64),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_67),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_25),
.B(n_0),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_70),
.Y(n_193)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_71),
.Y(n_162)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g154 ( 
.A(n_73),
.Y(n_154)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_76),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_80),
.B(n_88),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_82),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_83),
.Y(n_173)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_86),
.Y(n_180)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_87),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_58),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_89),
.Y(n_176)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_91),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_21),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_92),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_21),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_95),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_94),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_21),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_18),
.B(n_1),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_97),
.B(n_100),
.Y(n_158)
);

INVx11_ASAP7_75t_SL g98 ( 
.A(n_43),
.Y(n_98)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_27),
.B(n_1),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_24),
.B(n_1),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_103),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_24),
.B(n_17),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_27),
.B(n_2),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_104),
.B(n_110),
.Y(n_165)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_28),
.B(n_2),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_107),
.B(n_115),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_56),
.Y(n_109)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_109),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_29),
.B(n_2),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_111),
.B(n_119),
.Y(n_178)
);

BUFx16f_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

INVx6_ASAP7_75t_SL g114 ( 
.A(n_26),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_28),
.B(n_38),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_22),
.Y(n_117)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_42),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_118),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_22),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_120),
.B(n_122),
.Y(n_189)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_26),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_31),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_31),
.B(n_3),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_123),
.B(n_3),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_34),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_124),
.Y(n_159)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_34),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_125),
.B(n_5),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_32),
.B(n_14),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_44),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_47),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_128),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_60),
.B1(n_55),
.B2(n_50),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_140),
.A2(n_149),
.B1(n_187),
.B2(n_194),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_142),
.B(n_181),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_84),
.B(n_60),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_148),
.B(n_174),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_73),
.A2(n_35),
.B1(n_55),
.B2(n_46),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_152),
.A2(n_184),
.B1(n_188),
.B2(n_195),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_66),
.A2(n_44),
.B1(n_74),
.B2(n_102),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_156),
.A2(n_161),
.B1(n_163),
.B2(n_168),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_77),
.A2(n_38),
.B1(n_54),
.B2(n_32),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_117),
.A2(n_39),
.B1(n_54),
.B2(n_41),
.Y(n_163)
);

NAND2x1_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_59),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_166),
.B(n_205),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_67),
.A2(n_45),
.B1(n_39),
.B2(n_48),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_78),
.B(n_59),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_75),
.A2(n_48),
.B1(n_45),
.B2(n_41),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_175),
.A2(n_179),
.B1(n_198),
.B2(n_68),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_92),
.A2(n_33),
.B1(n_46),
.B2(n_35),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_124),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_73),
.A2(n_50),
.B1(n_33),
.B2(n_47),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_81),
.A2(n_59),
.B1(n_57),
.B2(n_47),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_186),
.A2(n_199),
.B1(n_108),
.B2(n_51),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_122),
.A2(n_59),
.B1(n_57),
.B2(n_47),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_190),
.B(n_197),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_98),
.A2(n_59),
.B1(n_57),
.B2(n_47),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_112),
.B(n_4),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_116),
.A2(n_57),
.B1(n_26),
.B2(n_42),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_83),
.A2(n_57),
.B1(n_26),
.B2(n_42),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_79),
.B(n_4),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_5),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_85),
.A2(n_51),
.B1(n_6),
.B2(n_8),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_201),
.A2(n_202),
.B1(n_118),
.B2(n_64),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_71),
.A2(n_51),
.B1(n_6),
.B2(n_8),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_112),
.B(n_5),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_5),
.Y(n_214)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_207),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_154),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_210),
.B(n_212),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_148),
.A2(n_109),
.B(n_70),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_211),
.A2(n_232),
.B(n_227),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_214),
.B(n_254),
.Y(n_288)
);

OR2x4_ASAP7_75t_L g215 ( 
.A(n_128),
.B(n_96),
.Y(n_215)
);

O2A1O1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_215),
.A2(n_232),
.B(n_153),
.C(n_137),
.Y(n_300)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_167),
.Y(n_216)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_217),
.Y(n_278)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_218),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_82),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_219),
.B(n_225),
.Y(n_287)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_220),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_L g221 ( 
.A1(n_159),
.A2(n_113),
.B1(n_94),
.B2(n_99),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_221),
.A2(n_242),
.B1(n_271),
.B2(n_173),
.Y(n_316)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_223),
.Y(n_294)
);

OAI22x1_ASAP7_75t_L g224 ( 
.A1(n_154),
.A2(n_89),
.B1(n_64),
.B2(n_76),
.Y(n_224)
);

OA21x2_ASAP7_75t_L g284 ( 
.A1(n_224),
.A2(n_176),
.B(n_182),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_128),
.B(n_61),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_141),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_226),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_170),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_228),
.Y(n_306)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_229),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_131),
.B(n_86),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_230),
.B(n_239),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_142),
.B(n_106),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_231),
.B(n_238),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_166),
.A2(n_121),
.B(n_87),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_132),
.Y(n_233)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_233),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_135),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_234),
.B(n_237),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_133),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_235),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_236),
.A2(n_257),
.B1(n_266),
.B2(n_268),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_189),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_127),
.B(n_165),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_178),
.B(n_89),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_240),
.B(n_267),
.Y(n_301)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_132),
.Y(n_241)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_241),
.Y(n_322)
);

OAI22xp33_ASAP7_75t_L g242 ( 
.A1(n_159),
.A2(n_181),
.B1(n_140),
.B2(n_169),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_243),
.A2(n_253),
.B1(n_260),
.B2(n_246),
.Y(n_324)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_244),
.Y(n_308)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_174),
.B(n_8),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_SL g319 ( 
.A(n_246),
.B(n_264),
.Y(n_319)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_160),
.Y(n_247)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_247),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_158),
.B(n_10),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_248),
.B(n_249),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_144),
.B(n_10),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_174),
.B(n_11),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_261),
.Y(n_291)
);

AOI21xp33_ASAP7_75t_L g251 ( 
.A1(n_150),
.A2(n_96),
.B(n_63),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_251),
.B(n_252),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_138),
.B(n_12),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_168),
.A2(n_179),
.B1(n_130),
.B2(n_139),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_147),
.B(n_12),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_191),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_256),
.B(n_262),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_151),
.A2(n_65),
.B1(n_12),
.B2(n_14),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_147),
.Y(n_258)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_258),
.Y(n_314)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_129),
.Y(n_259)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_259),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_130),
.A2(n_129),
.B1(n_139),
.B2(n_194),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_143),
.B(n_166),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_171),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_138),
.B(n_136),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_263),
.B(n_269),
.Y(n_304)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_149),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_141),
.Y(n_265)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_265),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_151),
.A2(n_170),
.B1(n_177),
.B2(n_155),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_149),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_177),
.A2(n_155),
.B1(n_183),
.B2(n_146),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_191),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_160),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_270),
.B(n_273),
.Y(n_328)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_204),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_276),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_136),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_146),
.A2(n_143),
.B1(n_196),
.B2(n_134),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_274),
.A2(n_172),
.B1(n_180),
.B2(n_164),
.Y(n_292)
);

INVx6_ASAP7_75t_SL g276 ( 
.A(n_171),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_187),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_169),
.Y(n_310)
);

AO22x1_ASAP7_75t_SL g283 ( 
.A1(n_211),
.A2(n_215),
.B1(n_275),
.B2(n_227),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_283),
.B(n_296),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_284),
.Y(n_374)
);

OAI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_243),
.A2(n_193),
.B1(n_162),
.B2(n_196),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_286),
.A2(n_324),
.B1(n_276),
.B2(n_317),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_182),
.C(n_172),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_289),
.B(n_312),
.C(n_323),
.Y(n_360)
);

OAI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_292),
.A2(n_316),
.B1(n_321),
.B2(n_330),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_227),
.A2(n_180),
.B1(n_164),
.B2(n_183),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_261),
.A2(n_162),
.B1(n_193),
.B2(n_176),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_298),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_300),
.Y(n_373)
);

NAND2xp33_ASAP7_75t_SL g368 ( 
.A(n_305),
.B(n_315),
.Y(n_368)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_310),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_231),
.A2(n_134),
.B1(n_145),
.B2(n_173),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_311),
.A2(n_326),
.B1(n_284),
.B2(n_301),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_222),
.B(n_145),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_225),
.B(n_137),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_315),
.Y(n_363)
);

O2A1O1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_209),
.A2(n_153),
.B(n_206),
.C(n_250),
.Y(n_317)
);

O2A1O1Ixp33_ASAP7_75t_L g355 ( 
.A1(n_317),
.A2(n_270),
.B(n_229),
.C(n_226),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_242),
.A2(n_206),
.B1(n_271),
.B2(n_208),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_318),
.A2(n_258),
.B1(n_259),
.B2(n_218),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_246),
.A2(n_255),
.B1(n_219),
.B2(n_224),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_238),
.B(n_249),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_213),
.A2(n_212),
.B1(n_221),
.B2(n_248),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_235),
.A2(n_256),
.B1(n_269),
.B2(n_247),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_264),
.A2(n_267),
.B1(n_233),
.B2(n_217),
.Y(n_331)
);

INVx8_ASAP7_75t_L g358 ( 
.A(n_331),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_313),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_334),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_335),
.A2(n_341),
.B1(n_372),
.B2(n_284),
.Y(n_384)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_322),
.Y(n_337)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_337),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_297),
.B(n_220),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_338),
.B(n_342),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_340),
.A2(n_301),
.B1(n_330),
.B2(n_292),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_305),
.A2(n_234),
.B1(n_223),
.B2(n_265),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_297),
.B(n_241),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_322),
.Y(n_343)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_343),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_309),
.B(n_233),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_344),
.B(n_345),
.Y(n_380)
);

A2O1A1Ixp33_ASAP7_75t_L g345 ( 
.A1(n_283),
.A2(n_207),
.B(n_216),
.C(n_277),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_312),
.B(n_245),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_346),
.B(n_348),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_300),
.A2(n_283),
.B(n_333),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_347),
.A2(n_354),
.B(n_306),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_287),
.B(n_272),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_328),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_349),
.B(n_356),
.Y(n_398)
);

A2O1A1Ixp33_ASAP7_75t_L g350 ( 
.A1(n_287),
.A2(n_289),
.B(n_281),
.C(n_319),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_350),
.B(n_359),
.Y(n_407)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_278),
.Y(n_351)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_351),
.Y(n_388)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_278),
.Y(n_352)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_352),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_303),
.A2(n_244),
.B(n_229),
.Y(n_354)
);

OA21x2_ASAP7_75t_L g399 ( 
.A1(n_355),
.A2(n_329),
.B(n_332),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_309),
.B(n_229),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_325),
.B(n_293),
.Y(n_357)
);

BUFx24_ASAP7_75t_SL g409 ( 
.A(n_357),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_291),
.B(n_304),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_302),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_361),
.Y(n_381)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_280),
.Y(n_362)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_362),
.Y(n_396)
);

INVx8_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_364),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_291),
.B(n_323),
.C(n_315),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_375),
.C(n_326),
.Y(n_377)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g382 ( 
.A(n_367),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_368),
.B(n_299),
.Y(n_383)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_308),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_302),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_370),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_327),
.B(n_280),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_371),
.B(n_294),
.Y(n_395)
);

MAJx2_ASAP7_75t_L g375 ( 
.A(n_327),
.B(n_321),
.C(n_296),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_299),
.Y(n_376)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_376),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_408),
.C(n_339),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_372),
.A2(n_318),
.B1(n_301),
.B2(n_316),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_378),
.A2(n_389),
.B1(n_390),
.B2(n_392),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_379),
.B(n_384),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_383),
.A2(n_400),
.B(n_411),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_347),
.A2(n_295),
.B1(n_288),
.B2(n_311),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_373),
.A2(n_310),
.B1(n_302),
.B2(n_314),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_373),
.A2(n_310),
.B1(n_320),
.B2(n_279),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_395),
.B(n_412),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_399),
.B(n_374),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_339),
.A2(n_279),
.B1(n_332),
.B2(n_294),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_401),
.A2(n_335),
.B1(n_341),
.B2(n_336),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_353),
.A2(n_285),
.B1(n_306),
.B2(n_290),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_402),
.A2(n_374),
.B1(n_370),
.B2(n_363),
.Y(n_417)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_337),
.Y(n_404)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_404),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_360),
.B(n_282),
.C(n_290),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_348),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_410),
.B(n_371),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_361),
.B(n_282),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_360),
.B(n_307),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_343),
.Y(n_413)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_413),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_412),
.B(n_350),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_421),
.C(n_426),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_381),
.B(n_349),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_415),
.B(n_423),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_406),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_416),
.B(n_419),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_417),
.A2(n_443),
.B1(n_444),
.B2(n_336),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_400),
.A2(n_366),
.B(n_339),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_418),
.A2(n_438),
.B(n_436),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_405),
.B(n_398),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_424),
.B(n_427),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_409),
.B(n_342),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_425),
.B(n_440),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_365),
.C(n_346),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_411),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_377),
.B(n_359),
.C(n_338),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_428),
.B(n_442),
.C(n_395),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_386),
.B(n_345),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_429),
.B(n_432),
.Y(n_462)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_403),
.Y(n_430)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_430),
.Y(n_458)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_403),
.Y(n_431)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_431),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_387),
.B(n_376),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_411),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_434),
.Y(n_449)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_385),
.Y(n_435)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_435),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_399),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_437),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_380),
.A2(n_366),
.B(n_354),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_399),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_439),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_391),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_407),
.B(n_375),
.C(n_368),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_394),
.B(n_369),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_447),
.A2(n_438),
.B(n_424),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_436),
.A2(n_383),
.B(n_407),
.Y(n_452)
);

OAI31xp33_ASAP7_75t_L g487 ( 
.A1(n_452),
.A2(n_470),
.A3(n_433),
.B(n_441),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_453),
.B(n_456),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_441),
.A2(n_384),
.B1(n_386),
.B2(n_402),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_454),
.A2(n_441),
.B1(n_378),
.B2(n_433),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_426),
.B(n_394),
.Y(n_456)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_457),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_415),
.A2(n_358),
.B1(n_413),
.B2(n_396),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_459),
.A2(n_437),
.B1(n_439),
.B2(n_443),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_421),
.B(n_383),
.C(n_389),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_467),
.C(n_450),
.Y(n_476)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_420),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_464),
.Y(n_486)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_420),
.Y(n_466)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_466),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_414),
.B(n_390),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_432),
.Y(n_468)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_468),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_418),
.A2(n_358),
.B(n_401),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_444),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_471),
.Y(n_493)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_422),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_473),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_423),
.Y(n_473)
);

OAI21xp33_ASAP7_75t_L g504 ( 
.A1(n_474),
.A2(n_449),
.B(n_455),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_476),
.B(n_465),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_453),
.B(n_445),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_478),
.B(n_467),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_428),
.C(n_445),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_479),
.B(n_488),
.C(n_478),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_448),
.B(n_425),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_480),
.B(n_487),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_469),
.B(n_456),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_483),
.B(n_485),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_484),
.B(n_454),
.Y(n_501)
);

BUFx24_ASAP7_75t_SL g485 ( 
.A(n_473),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_442),
.C(n_434),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_489),
.A2(n_494),
.B1(n_461),
.B2(n_471),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_446),
.B(n_416),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_490),
.B(n_498),
.Y(n_509)
);

FAx1_ASAP7_75t_SL g491 ( 
.A(n_452),
.B(n_429),
.CI(n_427),
.CON(n_491),
.SN(n_491)
);

OA21x2_ASAP7_75t_SL g513 ( 
.A1(n_491),
.A2(n_472),
.B(n_465),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_446),
.B(n_468),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_492),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_449),
.A2(n_455),
.B1(n_461),
.B2(n_451),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_462),
.A2(n_417),
.B1(n_435),
.B2(n_431),
.Y(n_495)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_495),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_451),
.B(n_422),
.Y(n_497)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_497),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_462),
.B(n_385),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_507),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_SL g520 ( 
.A1(n_501),
.A2(n_496),
.B1(n_494),
.B2(n_482),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_504),
.A2(n_513),
.B(n_491),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_506),
.A2(n_515),
.B1(n_518),
.B2(n_477),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_481),
.B(n_447),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_497),
.Y(n_508)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_508),
.Y(n_532)
);

NAND3xp33_ASAP7_75t_L g527 ( 
.A(n_510),
.B(n_479),
.C(n_486),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_475),
.B(n_470),
.Y(n_511)
);

INVxp33_ASAP7_75t_L g523 ( 
.A(n_511),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_516),
.C(n_517),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_475),
.A2(n_463),
.B1(n_458),
.B2(n_466),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_481),
.B(n_476),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_488),
.B(n_463),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_489),
.A2(n_458),
.B1(n_464),
.B2(n_392),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_505),
.A2(n_492),
.B(n_493),
.Y(n_519)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_519),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_520),
.A2(n_521),
.B1(n_382),
.B2(n_396),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_512),
.A2(n_496),
.B1(n_482),
.B2(n_474),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_509),
.A2(n_486),
.B(n_477),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_522),
.B(n_531),
.Y(n_535)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_503),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_525),
.B(n_527),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_526),
.B(n_529),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_517),
.A2(n_507),
.B(n_499),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_530),
.B(n_531),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_506),
.A2(n_487),
.B1(n_491),
.B2(n_430),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_504),
.A2(n_355),
.B(n_440),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_533),
.B(n_534),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_511),
.A2(n_404),
.B(n_388),
.Y(n_534)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_535),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_528),
.B(n_514),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_536),
.B(n_532),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_528),
.B(n_516),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_538),
.A2(n_540),
.B(n_367),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_523),
.B(n_510),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_524),
.B(n_502),
.C(n_500),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_SL g555 ( 
.A(n_543),
.B(n_544),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_524),
.B(n_501),
.C(n_515),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_526),
.B(n_518),
.C(n_382),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_545),
.B(n_548),
.C(n_544),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_547),
.A2(n_533),
.B1(n_542),
.B2(n_534),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_523),
.B(n_382),
.C(n_397),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_539),
.B(n_530),
.Y(n_549)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_549),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_546),
.Y(n_550)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_550),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_552),
.B(n_553),
.Y(n_567)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_548),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_554),
.B(n_559),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g556 ( 
.A1(n_537),
.A2(n_541),
.B(n_521),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g562 ( 
.A1(n_556),
.A2(n_537),
.B(n_542),
.Y(n_562)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_547),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_557),
.B(n_558),
.Y(n_560)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_562),
.Y(n_568)
);

AOI21x1_ASAP7_75t_L g564 ( 
.A1(n_549),
.A2(n_551),
.B(n_550),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_564),
.A2(n_555),
.B(n_388),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_552),
.B(n_545),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_565),
.B(n_543),
.Y(n_569)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_569),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_570),
.B(n_571),
.C(n_351),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_567),
.B(n_397),
.C(n_391),
.Y(n_571)
);

OAI322xp33_ASAP7_75t_L g572 ( 
.A1(n_563),
.A2(n_566),
.A3(n_560),
.B1(n_561),
.B2(n_393),
.C1(n_352),
.C2(n_362),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_572),
.A2(n_393),
.B(n_560),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_573),
.A2(n_334),
.B(n_329),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_574),
.A2(n_568),
.B1(n_571),
.B2(n_364),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_576),
.B(n_577),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_578),
.A2(n_575),
.B(n_334),
.Y(n_579)
);

XNOR2x2_ASAP7_75t_SL g580 ( 
.A(n_579),
.B(n_307),
.Y(n_580)
);


endmodule