module fake_jpeg_5171_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx4f_ASAP7_75t_SL g13 ( 
.A(n_7),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_6),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_34),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_14),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_35),
.A2(n_14),
.B1(n_13),
.B2(n_26),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_46),
.B1(n_47),
.B2(n_34),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_15),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_13),
.B(n_20),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_32),
.B(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_49),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_26),
.B1(n_25),
.B2(n_17),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_33),
.B1(n_20),
.B2(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_33),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_57),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_30),
.B1(n_32),
.B2(n_31),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_44),
.B1(n_43),
.B2(n_36),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_20),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_55),
.A2(n_59),
.B1(n_47),
.B2(n_49),
.Y(n_63)
);

AOI32xp33_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_28),
.A3(n_20),
.B1(n_33),
.B2(n_34),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_41),
.C(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_15),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_18),
.B1(n_24),
.B2(n_21),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_38),
.B1(n_18),
.B2(n_22),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_39),
.B1(n_25),
.B2(n_17),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_41),
.B1(n_36),
.B2(n_38),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_73),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_70),
.A2(n_62),
.B1(n_51),
.B2(n_56),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_38),
.C(n_19),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_51),
.C(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_18),
.B1(n_22),
.B2(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_62),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_86),
.C(n_21),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_80),
.B1(n_79),
.B2(n_81),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_62),
.C(n_55),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_80),
.C(n_87),
.Y(n_90)
);

AO32x1_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_62),
.A3(n_50),
.B1(n_53),
.B2(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_1),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_89),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_24),
.C(n_18),
.Y(n_86)
);

OAI21x1_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_24),
.B(n_22),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_24),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_86),
.A2(n_76),
.B(n_68),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_5),
.B(n_8),
.Y(n_110)
);

AOI221xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_64),
.B1(n_69),
.B2(n_63),
.C(n_74),
.Y(n_93)
);

NOR3xp33_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_2),
.C(n_3),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_98),
.C(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_75),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_70),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_99),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_12),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_95),
.B1(n_90),
.B2(n_92),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_81),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_104),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_106),
.C(n_110),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_11),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_11),
.C(n_3),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_2),
.B(n_3),
.C(n_5),
.D(n_6),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_108),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_98),
.A2(n_5),
.B(n_7),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_96),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_112),
.A2(n_105),
.B(n_108),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_9),
.B(n_10),
.Y(n_124)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_124),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_103),
.B1(n_106),
.B2(n_107),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_120),
.A2(n_122),
.B1(n_111),
.B2(n_118),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_113),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_127),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_121),
.B(n_118),
.Y(n_128)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_128),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_111),
.Y(n_129)
);

OAI311xp33_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_9),
.A3(n_10),
.B1(n_128),
.C1(n_126),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_10),
.B(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_9),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_134),
.Y(n_135)
);


endmodule