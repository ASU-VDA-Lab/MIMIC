module fake_jpeg_28445_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx5_ASAP7_75t_SL g45 ( 
.A(n_31),
.Y(n_45)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_38),
.Y(n_41)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_28),
.A2(n_16),
.B1(n_14),
.B2(n_12),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_51),
.B1(n_44),
.B2(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_26),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_50),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_25),
.C(n_14),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_30),
.A2(n_23),
.B1(n_22),
.B2(n_17),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_58),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_12),
.B1(n_16),
.B2(n_27),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_52),
.B1(n_49),
.B2(n_45),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_63),
.Y(n_84)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_13),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_61),
.B(n_66),
.Y(n_89)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_26),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_70),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_69),
.Y(n_91)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_72),
.Y(n_78)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_75),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_40),
.B1(n_27),
.B2(n_23),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_45),
.B1(n_20),
.B2(n_2),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_20),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_0),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_82),
.B(n_6),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_2),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_45),
.B1(n_20),
.B2(n_7),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_4),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_74),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_100),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_99),
.B(n_103),
.Y(n_108)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_102),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_62),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_104),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_9),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_9),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_106),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_90),
.B(n_85),
.Y(n_111)
);

NAND2x1_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_101),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_114),
.C(n_78),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_78),
.Y(n_114)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_110),
.B1(n_107),
.B2(n_121),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_111),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_90),
.C(n_94),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_120),
.C(n_114),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_94),
.C(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_124),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_86),
.Y(n_129)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_127),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_95),
.B1(n_106),
.B2(n_83),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_131),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_129),
.Y(n_135)
);

NAND4xp25_ASAP7_75t_SL g133 ( 
.A(n_128),
.B(n_91),
.C(n_77),
.D(n_11),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_10),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_136),
.B(n_134),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_130),
.B(n_132),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_10),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_69),
.Y(n_140)
);


endmodule