module fake_jpeg_28520_n_421 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_421);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_421;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_51),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_97),
.Y(n_104)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

BUFx12f_ASAP7_75t_SL g70 ( 
.A(n_31),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_87),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_20),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_20),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_76),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_20),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_84),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

BUFx4f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_79),
.Y(n_145)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_82),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_16),
.Y(n_84)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

BUFx16f_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_16),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_90),
.Y(n_133)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_92),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_96),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_23),
.B(n_1),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_95),
.Y(n_144)
);

BUFx24_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_28),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_32),
.B1(n_33),
.B2(n_47),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_101),
.A2(n_107),
.B1(n_114),
.B2(n_128),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_32),
.B1(n_28),
.B2(n_41),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_32),
.B1(n_33),
.B2(n_47),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_95),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_31),
.C(n_38),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_124),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_31),
.C(n_38),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_68),
.A2(n_41),
.B1(n_44),
.B2(n_38),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_53),
.A2(n_41),
.B1(n_44),
.B2(n_18),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_134),
.A2(n_146),
.B1(n_147),
.B2(n_150),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_55),
.A2(n_44),
.B1(n_43),
.B2(n_46),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_149),
.B(n_151),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_56),
.A2(n_15),
.B1(n_22),
.B2(n_18),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_66),
.A2(n_15),
.B1(n_22),
.B2(n_43),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_62),
.B(n_45),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_78),
.A2(n_45),
.B1(n_42),
.B2(n_39),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_86),
.B(n_42),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_83),
.B(n_39),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_46),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_93),
.A2(n_46),
.B1(n_92),
.B2(n_82),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_153),
.A2(n_46),
.B1(n_95),
.B2(n_71),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_162),
.Y(n_204)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_157),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_100),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_160),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_140),
.A2(n_57),
.B1(n_85),
.B2(n_67),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_161),
.A2(n_106),
.B1(n_108),
.B2(n_132),
.Y(n_201)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_163),
.Y(n_223)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_164),
.Y(n_197)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_23),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_169),
.Y(n_214)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_23),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_105),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_175),
.A2(n_178),
.B1(n_180),
.B2(n_182),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_46),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_179),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_137),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_104),
.B(n_71),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_187),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_137),
.Y(n_182)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_111),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_185),
.B1(n_190),
.B2(n_136),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_184),
.A2(n_191),
.B(n_192),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_188),
.B(n_189),
.Y(n_229)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_102),
.B(n_88),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_110),
.B(n_148),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_148),
.C(n_108),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_124),
.B(n_121),
.Y(n_194)
);

OAI32xp33_ASAP7_75t_L g219 ( 
.A1(n_194),
.A2(n_130),
.A3(n_138),
.B1(n_126),
.B2(n_145),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_200),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_162),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_159),
.A2(n_127),
.B1(n_136),
.B2(n_113),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_203),
.A2(n_208),
.B1(n_213),
.B2(n_217),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_195),
.A2(n_138),
.B1(n_106),
.B2(n_113),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_206),
.A2(n_215),
.B1(n_221),
.B2(n_165),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_186),
.A2(n_130),
.B1(n_142),
.B2(n_129),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_159),
.A2(n_181),
.B1(n_156),
.B2(n_186),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_138),
.B1(n_142),
.B2(n_122),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_177),
.A2(n_129),
.B1(n_122),
.B2(n_115),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_219),
.B(n_183),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_162),
.A2(n_126),
.B1(n_145),
.B2(n_132),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_170),
.A2(n_135),
.B1(n_118),
.B2(n_111),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_225),
.A2(n_227),
.B1(n_190),
.B2(n_185),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_160),
.A2(n_137),
.B(n_135),
.C(n_118),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_226),
.B(n_154),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_169),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_231),
.A2(n_197),
.B1(n_207),
.B2(n_180),
.Y(n_284)
);

NAND2xp33_ASAP7_75t_SL g232 ( 
.A(n_229),
.B(n_187),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_251),
.C(n_220),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_155),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_246),
.Y(n_268)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_222),
.Y(n_235)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_202),
.Y(n_237)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_238),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_196),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_239),
.B(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_244),
.Y(n_260)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_249),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_179),
.C(n_168),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_213),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_256),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_219),
.A2(n_189),
.B1(n_175),
.B2(n_171),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_250),
.B1(n_203),
.B2(n_231),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_228),
.Y(n_251)
);

CKINVDCx6p67_ASAP7_75t_R g252 ( 
.A(n_226),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_252),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_163),
.C(n_157),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_257),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_212),
.A2(n_214),
.B(n_209),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_199),
.B(n_224),
.Y(n_282)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_167),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_205),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_240),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_259),
.A2(n_214),
.B(n_209),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_261),
.A2(n_280),
.B1(n_164),
.B2(n_222),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_263),
.B(n_282),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_242),
.A2(n_206),
.B1(n_201),
.B2(n_221),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_264),
.A2(n_271),
.B1(n_276),
.B2(n_278),
.Y(n_297)
);

AO22x1_ASAP7_75t_L g265 ( 
.A1(n_252),
.A2(n_247),
.B1(n_242),
.B2(n_231),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_283),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_267),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_252),
.A2(n_244),
.B1(n_255),
.B2(n_234),
.Y(n_271)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_252),
.A2(n_217),
.B1(n_230),
.B2(n_210),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_234),
.A2(n_230),
.B1(n_196),
.B2(n_198),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_250),
.A2(n_227),
.B1(n_211),
.B2(n_220),
.Y(n_280)
);

OA21x2_ASAP7_75t_L g281 ( 
.A1(n_241),
.A2(n_211),
.B(n_197),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_281),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_199),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_254),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_224),
.Y(n_286)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_286),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_260),
.B(n_246),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_287),
.B(n_288),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_285),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_295),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_275),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_292),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_260),
.B(n_233),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_299),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_272),
.A2(n_249),
.B(n_253),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_238),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_298),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_265),
.A2(n_253),
.B1(n_258),
.B2(n_256),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_285),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_305),
.Y(n_323)
);

OAI21xp33_ASAP7_75t_L g301 ( 
.A1(n_279),
.A2(n_245),
.B(n_154),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_284),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_228),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_302),
.B(n_307),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_272),
.B(n_235),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_304),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_223),
.Y(n_306)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_306),
.Y(n_320)
);

XOR2x1_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_223),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_276),
.A2(n_192),
.B1(n_2),
.B2(n_4),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_308),
.A2(n_273),
.B1(n_270),
.B2(n_269),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_261),
.A2(n_192),
.B1(n_2),
.B2(n_4),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_308),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_277),
.C(n_268),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_312),
.C(n_328),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_277),
.C(n_278),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_313),
.B(n_294),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_314),
.Y(n_335)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_321),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_297),
.A2(n_274),
.B1(n_280),
.B2(n_266),
.Y(n_325)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_325),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_283),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_305),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_309),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_287),
.B(n_266),
.C(n_264),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_293),
.C(n_303),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_329),
.B(n_330),
.C(n_296),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_270),
.C(n_269),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_300),
.Y(n_331)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_331),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_332),
.A2(n_281),
.B1(n_262),
.B2(n_5),
.Y(n_351)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_333),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_292),
.Y(n_337)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_337),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_341),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_294),
.Y(n_342)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_342),
.Y(n_358)
);

AND3x1_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_307),
.C(n_290),
.Y(n_343)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_343),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_330),
.B(n_324),
.Y(n_344)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_344),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_319),
.B(n_296),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_345),
.B(n_348),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_290),
.Y(n_346)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_346),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_311),
.B(n_295),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_312),
.C(n_322),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_273),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_349),
.B(n_350),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_329),
.B(n_262),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_351),
.A2(n_327),
.B1(n_320),
.B2(n_315),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_316),
.Y(n_352)
);

INVx13_ASAP7_75t_L g363 ( 
.A(n_352),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_346),
.A2(n_318),
.B(n_317),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_347),
.Y(n_374)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_356),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_334),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_338),
.A2(n_317),
.B1(n_320),
.B2(n_323),
.Y(n_364)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_364),
.Y(n_372)
);

BUFx24_ASAP7_75t_SL g366 ( 
.A(n_344),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_366),
.B(n_342),
.Y(n_378)
);

OA21x2_ASAP7_75t_L g367 ( 
.A1(n_343),
.A2(n_323),
.B(n_310),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_367),
.B(n_337),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_365),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_369),
.B(n_373),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_359),
.B(n_334),
.C(n_348),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_375),
.C(n_381),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_374),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_341),
.Y(n_375)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_376),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_338),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_377),
.B(n_378),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_335),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_379),
.A2(n_380),
.B(n_353),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_354),
.B(n_339),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_322),
.C(n_326),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_371),
.A2(n_361),
.B(n_365),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_382),
.A2(n_367),
.B(n_357),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_370),
.A2(n_361),
.B(n_362),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_383),
.A2(n_389),
.B(n_374),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_362),
.C(n_355),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_386),
.B(n_375),
.Y(n_401)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_388),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_371),
.A2(n_368),
.B(n_358),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_372),
.A2(n_357),
.B1(n_358),
.B2(n_335),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_390),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_385),
.B(n_386),
.C(n_384),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_395),
.Y(n_405)
);

AO21x1_ASAP7_75t_L g406 ( 
.A1(n_394),
.A2(n_397),
.B(n_401),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_392),
.B(n_363),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_364),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_389),
.B(n_339),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_398),
.B(n_336),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_399),
.B(n_313),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_396),
.A2(n_391),
.B(n_385),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_402),
.B(n_332),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_403),
.B(n_408),
.Y(n_412)
);

AOI21xp33_ASAP7_75t_L g404 ( 
.A1(n_398),
.A2(n_387),
.B(n_336),
.Y(n_404)
);

BUFx24_ASAP7_75t_SL g411 ( 
.A(n_404),
.Y(n_411)
);

AOI31xp33_ASAP7_75t_L g407 ( 
.A1(n_400),
.A2(n_382),
.A3(n_367),
.B(n_381),
.Y(n_407)
);

A2O1A1Ixp33_ASAP7_75t_L g410 ( 
.A1(n_407),
.A2(n_333),
.B(n_351),
.C(n_281),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_405),
.B(n_397),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_409),
.B(n_410),
.C(n_413),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_412),
.A2(n_406),
.B(n_281),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_414),
.A2(n_415),
.B(n_9),
.Y(n_417)
);

AOI321xp33_ASAP7_75t_L g415 ( 
.A1(n_411),
.A2(n_1),
.A3(n_4),
.B1(n_5),
.B2(n_7),
.C(n_8),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g419 ( 
.A1(n_417),
.A2(n_418),
.B(n_9),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_416),
.B(n_9),
.C(n_12),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_419),
.B(n_9),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_420),
.B(n_12),
.C(n_352),
.Y(n_421)
);


endmodule