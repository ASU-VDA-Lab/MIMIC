module real_jpeg_6888_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_1),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_1),
.Y(n_108)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_1),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_2),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_2),
.A2(n_42),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_2),
.A2(n_42),
.B1(n_112),
.B2(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_2),
.A2(n_42),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_2),
.B(n_147),
.C(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_2),
.B(n_246),
.Y(n_245)
);

O2A1O1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_2),
.A2(n_253),
.B(n_255),
.C(n_256),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_2),
.B(n_266),
.C(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_2),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_2),
.B(n_212),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_2),
.B(n_21),
.Y(n_292)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_4),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_4),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_4),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_5),
.Y(n_367)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_6),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_7),
.A2(n_46),
.B1(n_50),
.B2(n_53),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_7),
.A2(n_38),
.B1(n_53),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_7),
.A2(n_53),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_7),
.A2(n_53),
.B1(n_71),
.B2(n_185),
.Y(n_184)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_9),
.Y(n_125)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_9),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_9),
.Y(n_231)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_10),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_11),
.A2(n_80),
.B1(n_84),
.B2(n_87),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_11),
.A2(n_87),
.B1(n_111),
.B2(n_114),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_11),
.A2(n_87),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_11),
.A2(n_87),
.B1(n_160),
.B2(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_12),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_362),
.B(n_364),
.Y(n_13)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_135),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_133),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_128),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_17),
.B(n_128),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_116),
.C(n_127),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_18),
.A2(n_19),
.B1(n_358),
.B2(n_359),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_44),
.C(n_88),
.Y(n_19)
);

XNOR2x1_ASAP7_75t_L g142 ( 
.A(n_20),
.B(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_20),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_20),
.B(n_200),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_20),
.A2(n_177),
.B1(n_178),
.B2(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_20),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_20),
.A2(n_219),
.B1(n_249),
.B2(n_259),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_20),
.B(n_169),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_20),
.A2(n_219),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_20),
.A2(n_177),
.B(n_215),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_20),
.A2(n_219),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_20),
.A2(n_219),
.B1(n_349),
.B2(n_350),
.Y(n_348)
);

OA21x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_31),
.B(n_40),
.Y(n_20)
);

NOR2x1_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_21),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_27),
.Y(n_146)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_31),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_32)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_33),
.Y(n_130)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_42),
.A2(n_68),
.B(n_71),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_44),
.A2(n_88),
.B1(n_89),
.B2(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_44),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_54),
.B1(n_67),
.B2(n_79),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_45),
.A2(n_54),
.B1(n_67),
.B2(n_144),
.Y(n_340)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AO21x1_ASAP7_75t_L g127 ( 
.A1(n_54),
.A2(n_67),
.B(n_79),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AO21x2_ASAP7_75t_SL g143 ( 
.A1(n_55),
.A2(n_67),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_67),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_56)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_57),
.Y(n_254)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_61),
.Y(n_147)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_67),
.Y(n_246)
);

OA22x2_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_70),
.B1(n_73),
.B2(n_76),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_86),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_88),
.A2(n_89),
.B1(n_340),
.B2(n_341),
.Y(n_339)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_89),
.B(n_219),
.C(n_340),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_99),
.B(n_110),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_90),
.B(n_99),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_90),
.A2(n_99),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_90),
.Y(n_210)
);

NAND2x1_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_99),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_98),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_94),
.Y(n_267)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_99),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_105),
.B2(n_109),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_100),
.B(n_276),
.Y(n_275)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_102),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_102),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_110),
.Y(n_211)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g268 ( 
.A(n_113),
.Y(n_268)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_116),
.B(n_127),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_126),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_119),
.B1(n_126),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_356),
.B(n_361),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_334),
.B(n_353),
.Y(n_136)
);

OAI211xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_239),
.B(n_328),
.C(n_333),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_221),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g328 ( 
.A1(n_139),
.A2(n_221),
.B(n_329),
.C(n_332),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_203),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_140),
.B(n_203),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_176),
.C(n_188),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_141),
.B(n_176),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_148),
.B1(n_174),
.B2(n_175),
.Y(n_141)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_142),
.B(n_189),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_142),
.A2(n_174),
.B1(n_228),
.B2(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_143),
.B(n_209),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_143),
.A2(n_202),
.B(n_219),
.C(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_143),
.A2(n_169),
.B1(n_200),
.B2(n_225),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_143),
.A2(n_200),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_148),
.A2(n_199),
.B(n_201),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_169),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_149),
.A2(n_169),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_149),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_156),
.B1(n_162),
.B2(n_166),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_154),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_150),
.A2(n_156),
.B1(n_191),
.B2(n_197),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_152),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_155),
.Y(n_198)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_166),
.B(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_169),
.B(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_169),
.A2(n_225),
.B1(n_245),
.B2(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_169),
.A2(n_225),
.B1(n_263),
.B2(n_264),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_169),
.A2(n_225),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

O2A1O1Ixp33_ASAP7_75t_L g296 ( 
.A1(n_169),
.A2(n_200),
.B(n_251),
.C(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_169),
.B(n_200),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_169),
.A2(n_190),
.B1(n_225),
.B2(n_319),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_181),
.B2(n_187),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_181),
.Y(n_216)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_180),
.B(n_192),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_184),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_209)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_188),
.B(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_199),
.B(n_201),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_190),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_200),
.A2(n_208),
.B(n_213),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_200),
.B(n_236),
.C(n_291),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AND3x1_ASAP7_75t_L g321 ( 
.A(n_202),
.B(n_298),
.C(n_322),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_220),
.Y(n_203)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_214),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_207),
.B(n_214),
.C(n_220),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

FAx1_ASAP7_75t_L g336 ( 
.A(n_213),
.B(n_337),
.CI(n_342),
.CON(n_336),
.SN(n_336)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_219),
.B(n_348),
.C(n_352),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_237),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_222),
.B(n_237),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.C(n_227),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_223),
.B(n_224),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_245),
.C(n_247),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_225),
.B(n_288),
.C(n_295),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_227),
.B(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_228),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_236),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_229),
.A2(n_230),
.B1(n_236),
.B2(n_247),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_236),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_236),
.A2(n_247),
.B1(n_252),
.B2(n_258),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_236),
.B(n_283),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_236),
.A2(n_247),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_236),
.B(n_252),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_310),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_300),
.B(n_309),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_286),
.B(n_299),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_260),
.B(n_285),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_244),
.B(n_248),
.Y(n_285)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_247),
.B(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_247),
.B(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_259),
.Y(n_248)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_272),
.B(n_284),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_269),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_269),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_282),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_280),
.Y(n_273)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_296),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_296),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_293),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_302),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_306),
.C(n_307),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_323),
.Y(n_310)
);

NOR2x1_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_313),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_316),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_320),
.B2(n_321),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_320),
.C(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_323),
.A2(n_330),
.B(n_331),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_326),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_326),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_344),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_343),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_336),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_343),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_345),
.Y(n_355)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_340),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_344),
.A2(n_354),
.B(n_355),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_352),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_360),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_357),
.B(n_360),
.Y(n_361)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx6_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx13_ASAP7_75t_L g366 ( 
.A(n_363),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);


endmodule