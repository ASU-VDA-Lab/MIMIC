module real_jpeg_67_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_288;
wire n_166;
wire n_176;
wire n_300;
wire n_221;
wire n_215;
wire n_249;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_293;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_70;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_41;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_297;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_209;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_244;
wire n_213;
wire n_133;
wire n_216;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_1),
.A2(n_44),
.B1(n_45),
.B2(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_1),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_1),
.A2(n_62),
.B1(n_63),
.B2(n_85),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_1),
.A2(n_39),
.B1(n_40),
.B2(n_85),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_1),
.A2(n_29),
.B1(n_34),
.B2(n_85),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_53),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_2),
.A2(n_53),
.B1(n_62),
.B2(n_63),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_2),
.A2(n_29),
.B1(n_34),
.B2(n_53),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_3),
.A2(n_62),
.B1(n_63),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_29),
.B1(n_34),
.B2(n_72),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_72),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_5),
.B(n_150),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_5),
.B(n_63),
.C(n_81),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_5),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_5),
.B(n_80),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_5),
.B(n_29),
.C(n_65),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_185),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_5),
.B(n_31),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_5),
.B(n_98),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_185),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_6),
.Y(n_81)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_8),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_8),
.A2(n_35),
.B1(n_62),
.B2(n_63),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_11),
.A2(n_62),
.B1(n_63),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_70),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_11),
.A2(n_29),
.B1(n_34),
.B2(n_70),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_13),
.A2(n_39),
.B1(n_40),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_13),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_104),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_104),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_13),
.A2(n_29),
.B1(n_34),
.B2(n_104),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_14),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_14),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_14),
.A2(n_42),
.B1(n_62),
.B2(n_63),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_14),
.A2(n_29),
.B1(n_34),
.B2(n_42),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_15),
.A2(n_39),
.B1(n_40),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_15),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_149),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_15),
.A2(n_62),
.B1(n_63),
.B2(n_149),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_15),
.A2(n_29),
.B1(n_34),
.B2(n_149),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_125),
.B1(n_299),
.B2(n_300),
.Y(n_18)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_19),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_108),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_21),
.B(n_108),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_74),
.C(n_89),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_22),
.A2(n_23),
.B1(n_74),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_57),
.B2(n_73),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_36),
.B1(n_37),
.B2(n_56),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_26),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_26),
.A2(n_37),
.B(n_73),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_26),
.A2(n_56),
.B1(n_58),
.B2(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_31),
.B(n_32),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_27),
.A2(n_31),
.B1(n_94),
.B2(n_142),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_27),
.A2(n_185),
.B(n_212),
.Y(n_232)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_28),
.A2(n_30),
.B1(n_33),
.B2(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_28),
.A2(n_30),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_28),
.B(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_28),
.A2(n_30),
.B1(n_165),
.B2(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_28),
.A2(n_210),
.B(n_211),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_28),
.A2(n_30),
.B1(n_210),
.B2(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_29),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_29),
.A2(n_34),
.B1(n_65),
.B2(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_29),
.B(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_30),
.A2(n_164),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_30),
.B(n_179),
.Y(n_212)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_31),
.A2(n_178),
.B(n_235),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B(n_50),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_38),
.A2(n_43),
.B1(n_105),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_40),
.B1(n_47),
.B2(n_48),
.Y(n_55)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_40),
.A2(n_105),
.B(n_185),
.C(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_40),
.B(n_185),
.Y(n_186)
);

AOI32xp33_ASAP7_75t_L g197 ( 
.A1(n_40),
.A2(n_45),
.A3(n_47),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_43),
.B(n_52),
.Y(n_107)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_43),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_43),
.A2(n_50),
.B(n_271),
.Y(n_270)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_44),
.A2(n_45),
.B1(n_81),
.B2(n_82),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_44),
.B(n_175),
.Y(n_174)
);

NAND2xp33_ASAP7_75t_SL g199 ( 
.A(n_44),
.B(n_48),
.Y(n_199)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_54),
.A2(n_103),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_58),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_67),
.B1(n_71),
.B2(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_59),
.A2(n_170),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_59),
.A2(n_67),
.B1(n_168),
.B2(n_218),
.Y(n_252)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_69),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_60),
.A2(n_98),
.B(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_60),
.A2(n_97),
.B1(n_98),
.B2(n_140),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_60),
.A2(n_167),
.B(n_169),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_60),
.B(n_171),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_67),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_63),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_63),
.B(n_224),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_67),
.A2(n_191),
.B(n_192),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_67),
.A2(n_192),
.B(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_77),
.B(n_88),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_77),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_78),
.A2(n_84),
.B1(n_86),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_86),
.B1(n_87),
.B2(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_78),
.A2(n_86),
.B1(n_158),
.B2(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_78),
.A2(n_250),
.B(n_251),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_78),
.A2(n_189),
.B(n_251),
.Y(n_269)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_79),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_80),
.B(n_146),
.Y(n_251)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_86),
.A2(n_100),
.B(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_86),
.A2(n_145),
.B(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_99),
.C(n_101),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_91),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_92),
.A2(n_95),
.B1(n_96),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_92),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_98),
.B(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_99),
.B(n_101),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_105),
.B(n_106),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_107),
.B(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_122),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_114),
.B2(n_121),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_125),
.Y(n_300)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_151),
.B(n_298),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_127),
.B(n_130),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.C(n_136),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_131),
.B(n_134),
.Y(n_296)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_136),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_143),
.C(n_147),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_137),
.A2(n_138),
.B1(n_286),
.B2(n_288),
.Y(n_285)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_139),
.B(n_141),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_140),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_142),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_143),
.A2(n_144),
.B1(n_147),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_147),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_148),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_293),
.B(n_297),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_262),
.B(n_290),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_204),
.B(n_261),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_180),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_155),
.B(n_180),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_166),
.C(n_172),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_156),
.B(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_160),
.C(n_163),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_166),
.B(n_172),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_176),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_194),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_181),
.B(n_195),
.C(n_203),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_187),
.B2(n_193),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_182),
.B(n_188),
.C(n_190),
.Y(n_275)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_203),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_196),
.B(n_201),
.Y(n_266)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_256),
.B(n_260),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_245),
.B(n_255),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_227),
.B(n_244),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_221),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_221),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_213),
.B1(n_219),
.B2(n_220),
.Y(n_208)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_216),
.C(n_219),
.Y(n_246)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_238),
.B(n_243),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_233),
.B(n_237),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_236),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_235),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_241),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_247),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_253),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_252),
.C(n_253),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_259),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_277),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_276),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_276),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_273),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_274),
.C(n_275),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_268),
.C(n_272),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_272),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_270),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_289),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_289),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_283),
.C(n_285),
.Y(n_294)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_295),
.Y(n_297)
);


endmodule