module real_jpeg_26423_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_0),
.B(n_25),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_0),
.B(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_0),
.B(n_60),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_0),
.B(n_39),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_0),
.B(n_43),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_0),
.B(n_27),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_0),
.B(n_16),
.Y(n_171)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_2),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_2),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_2),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_2),
.B(n_27),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_2),
.B(n_43),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_2),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_3),
.B(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_3),
.B(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_4),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_4),
.B(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_4),
.B(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_4),
.B(n_27),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_4),
.B(n_142),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_6),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_8),
.Y(n_105)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_27),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_12),
.B(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_12),
.B(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_13),
.B(n_30),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_13),
.B(n_60),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_13),
.B(n_25),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_13),
.B(n_39),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_13),
.B(n_27),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_15),
.B(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_15),
.B(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_15),
.B(n_25),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_15),
.B(n_39),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_15),
.B(n_43),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_15),
.B(n_27),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_15),
.B(n_181),
.Y(n_180)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_16),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_124),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_109),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_72),
.B2(n_108),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_45),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_31),
.C(n_37),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_23),
.B(n_122),
.Y(n_121)
);

BUFx24_ASAP7_75t_SL g199 ( 
.A(n_23),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_26),
.CI(n_29),
.CON(n_23),
.SN(n_23)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_24),
.B(n_26),
.C(n_29),
.Y(n_98)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_31),
.A2(n_32),
.B1(n_37),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_37),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.C(n_42),
.Y(n_37)
);

FAx1_ASAP7_75t_SL g114 ( 
.A(n_38),
.B(n_41),
.CI(n_42),
.CON(n_114),
.SN(n_114)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_43),
.Y(n_177)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_55),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_53),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_64),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_63),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_59),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_70),
.C(n_71),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_66),
.B(n_177),
.Y(n_176)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_71),
.Y(n_75)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_96),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.C(n_83),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_76),
.B1(n_77),
.B2(n_112),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_74),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B(n_82),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_81),
.Y(n_82)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_92),
.C(n_94),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_84),
.A2(n_85),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_92),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_100),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_104),
.CI(n_107),
.CON(n_100),
.SN(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.C(n_120),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_110),
.B(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_113),
.A2(n_120),
.B1(n_121),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_113),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.C(n_119),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_114),
.B(n_189),
.Y(n_188)
);

BUFx24_ASAP7_75t_SL g202 ( 
.A(n_114),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_115),
.B(n_119),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.C(n_118),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_195),
.C(n_196),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_186),
.C(n_187),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_148),
.C(n_160),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_138),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_136),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_129),
.B(n_136),
.C(n_138),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_134),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_131),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_145),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_139),
.B(n_146),
.C(n_147),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_159),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_153),
.B1(n_159),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_164)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_182),
.C(n_183),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_169),
.C(n_174),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_167),
.C(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.C(n_178),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_191),
.C(n_194),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);


endmodule