module real_jpeg_22660_n_12 (n_5, n_4, n_8, n_0, n_318, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_318;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_0),
.A2(n_20),
.B1(n_21),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_0),
.A2(n_32),
.B1(n_44),
.B2(n_45),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_0),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_112)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_3),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_3),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_3),
.B(n_168),
.Y(n_167)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_3),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_3),
.B(n_157),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_5),
.A2(n_20),
.B1(n_21),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_5),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_118),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_118),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_118),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_6),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_6),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_6),
.A2(n_22),
.B1(n_44),
.B2(n_45),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_6),
.A2(n_22),
.B1(n_38),
.B2(n_39),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_8),
.A2(n_38),
.B1(n_39),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_50),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_8),
.A2(n_20),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_8),
.B(n_20),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_8),
.B(n_70),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_50),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g172 ( 
.A1(n_8),
.A2(n_10),
.B(n_44),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_8),
.B(n_53),
.Y(n_194)
);

O2A1O1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_8),
.A2(n_24),
.B(n_55),
.C(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_9),
.A2(n_20),
.B(n_23),
.C(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_20),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_38),
.B(n_42),
.C(n_43),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_10),
.B(n_38),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_10),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_11),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_96),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_94),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_81),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_15),
.B(n_81),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_68),
.C(n_76),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_16),
.A2(n_17),
.B1(n_68),
.B2(n_304),
.Y(n_310)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_33),
.B1(n_34),
.B2(n_67),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_18),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_23),
.B(n_27),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_23),
.B(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_23),
.A2(n_29),
.B(n_74),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_24),
.A2(n_54),
.B(n_55),
.C(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_24),
.B(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_24),
.B(n_26),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_25),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_28),
.B(n_116),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_29),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_30),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_51),
.B1(n_65),
.B2(n_66),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_35),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_35),
.B(n_66),
.C(n_67),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_35),
.A2(n_65),
.B1(n_119),
.B2(n_120),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_35),
.A2(n_65),
.B1(n_77),
.B2(n_307),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_47),
.B(n_48),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_36),
.A2(n_111),
.B(n_250),
.Y(n_276)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_37),
.B(n_49),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_37),
.B(n_176),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_37),
.B(n_112),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_39),
.B1(n_55),
.B2(n_57),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_38),
.A2(n_50),
.B(n_57),
.Y(n_208)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_39),
.A2(n_46),
.B(n_50),
.C(n_172),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_43),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_43),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_43),
.B(n_49),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_44),
.B(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_45),
.B(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_47),
.B(n_50),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_47),
.A2(n_213),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_50),
.B(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_59),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_52),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_53),
.B(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_54),
.B(n_64),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_61),
.B(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_54),
.A2(n_59),
.B(n_79),
.Y(n_287)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_58),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_58),
.B(n_60),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_59),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_78),
.B(n_80),
.Y(n_77)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_61),
.B(n_132),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_68),
.C(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_115),
.C(n_119),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_68),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_68),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_69),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_69),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_70),
.B(n_270),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_74),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_76),
.B(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_77),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_80),
.B(n_131),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_80),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_88),
.B2(n_90),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B(n_87),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_85),
.B(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_88),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_88),
.A2(n_90),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_90),
.B(n_252),
.C(n_255),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI321xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_301),
.A3(n_311),
.B1(n_314),
.B2(n_315),
.C(n_318),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_280),
.B(n_300),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_259),
.B(n_279),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_159),
.B(n_242),
.C(n_258),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_146),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_101),
.B(n_146),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_123),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_114),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_103),
.B(n_114),
.C(n_123),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_110),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_104),
.B(n_110),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_107),
.B(n_108),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_105),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_105),
.A2(n_158),
.B(n_186),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_107),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_108),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_111),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_113),
.B(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_117),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_121),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_134),
.B1(n_135),
.B2(n_145),
.Y(n_123)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_133),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_125),
.B(n_133),
.C(n_134),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_127),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_136),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_138),
.B(n_199),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_139),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_168),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_150),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_147),
.B(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.C(n_154),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_152),
.B(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_153),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_167),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_241),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_235),
.B(n_240),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_220),
.B(n_234),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_201),
.B(n_219),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_189),
.B(n_200),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_177),
.B(n_188),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_169),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_171),
.B(n_173),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_182),
.B(n_187),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_180),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_191),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_198),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_196),
.C(n_198),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_203),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_210),
.B1(n_211),
.B2(n_218),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_204),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_209),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_205),
.A2(n_206),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_205),
.A2(n_206),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_205),
.A2(n_293),
.B(n_295),
.Y(n_308)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_207),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_206),
.B(n_276),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_214),
.B1(n_215),
.B2(n_217),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_212),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_213),
.B(n_230),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_217),
.C(n_218),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_216),
.B(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_221),
.B(n_222),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_227),
.B2(n_228),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_229),
.C(n_233),
.Y(n_236)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_229),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_231),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_236),
.B(n_237),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_243),
.B(n_244),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_256),
.B2(n_257),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_251),
.C(n_257),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_249),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_256),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_260),
.B(n_261),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_278),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_274),
.B2(n_275),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_275),
.C(n_278),
.Y(n_281)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_267),
.C(n_273),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_271),
.B2(n_273),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_271),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_276),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_281),
.B(n_282),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_298),
.B2(n_299),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_289),
.B1(n_296),
.B2(n_297),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_285),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_297),
.C(n_299),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B(n_288),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_287),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_303),
.C(n_308),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g313 ( 
.A(n_288),
.B(n_303),
.CI(n_308),
.CON(n_313),
.SN(n_313)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_289),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_290),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_291),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_298),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_309),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_309),
.Y(n_315)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_312),
.B(n_313),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_313),
.Y(n_316)
);


endmodule