module real_jpeg_19929_n_11 (n_5, n_4, n_8, n_0, n_256, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_256;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_247;
wire n_146;
wire n_249;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_240;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_244;
wire n_213;
wire n_179;
wire n_128;
wire n_167;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_0),
.A2(n_2),
.B1(n_16),
.B2(n_17),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_0),
.A2(n_6),
.B1(n_16),
.B2(n_23),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_0),
.A2(n_5),
.B1(n_16),
.B2(n_46),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_0),
.A2(n_4),
.B1(n_16),
.B2(n_40),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_1),
.A2(n_2),
.B1(n_17),
.B2(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_1),
.A2(n_6),
.B1(n_23),
.B2(n_25),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_1),
.A2(n_4),
.B1(n_25),
.B2(n_40),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_1),
.A2(n_5),
.B1(n_25),
.B2(n_46),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

A2O1A1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_2),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_20),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_2),
.A2(n_10),
.B1(n_17),
.B2(n_33),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_2),
.A2(n_20),
.B(n_33),
.C(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_3),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_4),
.A2(n_7),
.B1(n_38),
.B2(n_40),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_4),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_4),
.A2(n_9),
.B1(n_40),
.B2(n_47),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_4),
.A2(n_10),
.B1(n_33),
.B2(n_40),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_4),
.A2(n_33),
.B(n_47),
.C(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_5),
.A2(n_9),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_5),
.B(n_79),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_5),
.A2(n_10),
.B1(n_33),
.B2(n_46),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_5),
.A2(n_9),
.B(n_10),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_6),
.A2(n_8),
.B1(n_20),
.B2(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_7),
.B1(n_23),
.B2(n_38),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_6),
.A2(n_10),
.B1(n_23),
.B2(n_33),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_SL g91 ( 
.A1(n_6),
.A2(n_10),
.B(n_92),
.Y(n_91)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_7),
.A2(n_10),
.B(n_23),
.C(n_137),
.Y(n_136)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_10),
.B(n_26),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_10),
.B(n_39),
.Y(n_119)
);

AO21x1_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_249),
.B(n_252),
.Y(n_11)
);

OAI21xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_56),
.B(n_248),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_27),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_14),
.B(n_27),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_14),
.B(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_14),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_18),
.B1(n_24),
.B2(n_26),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_15),
.A2(n_18),
.B1(n_26),
.B2(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_19),
.B(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_24),
.B(n_31),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_51),
.C(n_52),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_28),
.A2(n_29),
.B1(n_244),
.B2(n_246),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.C(n_42),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_30),
.B(n_70),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_30),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_30),
.A2(n_68),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_30),
.A2(n_70),
.B(n_88),
.C(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_30),
.A2(n_68),
.B1(n_188),
.B2(n_189),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_30),
.A2(n_68),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_30),
.A2(n_189),
.B(n_208),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_30),
.A2(n_68),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_30),
.A2(n_68),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_33),
.B(n_45),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_33),
.B(n_82),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_33),
.A2(n_38),
.B(n_40),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_34),
.A2(n_42),
.B1(n_218),
.B2(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_34),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_39),
.B2(n_41),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_35),
.A2(n_36),
.B1(n_39),
.B2(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_42),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_42),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_50),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_44),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_45),
.B(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_45),
.A2(n_48),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OA22x2_ASAP7_75t_SL g204 ( 
.A1(n_45),
.A2(n_48),
.B1(n_50),
.B2(n_193),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_46),
.B(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_51),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_241),
.B(n_247),
.Y(n_56)
);

OAI321xp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_213),
.A3(n_233),
.B1(n_239),
.B2(n_240),
.C(n_256),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_198),
.B(n_212),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_180),
.B(n_197),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_107),
.B(n_162),
.C(n_179),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_96),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_62),
.B(n_96),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_85),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_75),
.B2(n_76),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_64),
.B(n_76),
.C(n_85),
.Y(n_163)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI211xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_68),
.B(n_69),
.C(n_74),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_73),
.B1(n_77),
.B2(n_84),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_66),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_66),
.A2(n_73),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_66),
.A2(n_73),
.B1(n_114),
.B2(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_66),
.B(n_93),
.C(n_118),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_66),
.A2(n_73),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_66),
.B(n_145),
.C(n_151),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_66),
.A2(n_73),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_66),
.B(n_77),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_66),
.B(n_169),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_67),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_68),
.B(n_71),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_68),
.B(n_218),
.C(n_220),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_68),
.B(n_227),
.C(n_232),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_69),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_70),
.A2(n_73),
.B(n_139),
.C(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_70),
.A2(n_71),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_70),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_70),
.B(n_204),
.Y(n_205)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_93),
.C(n_105),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_72),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_73),
.B(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_74),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_79),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_78),
.A2(n_82),
.B1(n_83),
.B2(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_95),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_86),
.A2(n_87),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_86),
.A2(n_87),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_103),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_103),
.B1(n_117),
.B2(n_120),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_93),
.A2(n_103),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_93),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_148)
);

NAND2x1_ASAP7_75t_SL g152 ( 
.A(n_93),
.B(n_136),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_94),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.C(n_104),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_97),
.A2(n_98),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_99),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_100),
.B1(n_135),
.B2(n_139),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_101),
.A2(n_102),
.B1(n_104),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_104),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_161),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_154),
.B(n_160),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_141),
.B(n_153),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_132),
.B(n_140),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_121),
.B(n_131),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_116),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_114),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_117),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_128),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_134),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_135),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_136),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_142),
.B(n_144),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_155),
.B(n_156),
.Y(n_160)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_164),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_176),
.B2(n_178),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_171),
.B1(n_174),
.B2(n_175),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_167),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_175),
.C(n_178),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_171),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_172),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_172),
.A2(n_177),
.B(n_196),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_176),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_SL g210 ( 
.A1(n_177),
.A2(n_185),
.B(n_196),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_181),
.B(n_182),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_183),
.B(n_199),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_187),
.CI(n_195),
.CON(n_183),
.SN(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_185),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_191),
.B2(n_194),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_191),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_191),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_210),
.B2(n_211),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_206),
.B2(n_207),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_207),
.C(n_211),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_205),
.A2(n_215),
.B1(n_222),
.B2(n_237),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_210),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_225),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_225),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_222),
.C(n_223),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_215),
.Y(n_237)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_223),
.A2(n_224),
.B1(n_236),
.B2(n_238),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_232),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_234),
.B(n_235),
.Y(n_239)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_236),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_244),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);


endmodule