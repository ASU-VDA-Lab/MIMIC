module fake_jpeg_109_n_222 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_222);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_23),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_52),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_2),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_3),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_3),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_38),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_14),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_14),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_84),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_22),
.B(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_80),
.B(n_57),
.Y(n_93)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_60),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_51),
.C(n_49),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_0),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_58),
.B1(n_57),
.B2(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_86),
.A2(n_84),
.B1(n_78),
.B2(n_63),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_87),
.Y(n_100)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_83),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_96),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_64),
.B1(n_74),
.B2(n_69),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_84),
.B1(n_79),
.B2(n_81),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_70),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

BUFx4f_ASAP7_75t_SL g108 ( 
.A(n_99),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_64),
.B1(n_74),
.B2(n_81),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_107),
.B1(n_113),
.B2(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_54),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_85),
.C(n_68),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_118),
.Y(n_119)
);

NAND2x1p5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_80),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_78),
.B1(n_69),
.B2(n_72),
.Y(n_114)
);

BUFx2_ASAP7_75t_SL g115 ( 
.A(n_89),
.Y(n_115)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_70),
.B1(n_53),
.B2(n_67),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_116),
.A2(n_66),
.B(n_55),
.Y(n_124)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_68),
.B1(n_59),
.B2(n_62),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_120),
.A2(n_124),
.B(n_1),
.Y(n_146)
);

OAI32xp33_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_72),
.A3(n_62),
.B1(n_65),
.B2(n_75),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_2),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_59),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_130),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_136),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_99),
.B1(n_89),
.B2(n_75),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_129),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_116),
.A2(n_99),
.B1(n_89),
.B2(n_65),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_117),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_61),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_132),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_71),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_76),
.B1(n_89),
.B2(n_99),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_101),
.B(n_0),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_77),
.B(n_47),
.C(n_44),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_139),
.A2(n_108),
.B(n_35),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_146),
.C(n_147),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_123),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_150),
.Y(n_180)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_144),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_137),
.A2(n_111),
.B1(n_77),
.B2(n_4),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_148),
.B1(n_9),
.B2(n_10),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_138),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_5),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_151),
.B(n_158),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_43),
.C(n_42),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_156),
.C(n_161),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_133),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_160),
.C(n_162),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_6),
.C(n_7),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_154),
.A2(n_135),
.B(n_10),
.Y(n_167)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_39),
.C(n_37),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

CKINVDCx12_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_7),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_36),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_8),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_33),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_168),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_122),
.B(n_129),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_159),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_170),
.Y(n_185)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_9),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_176),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

A2O1A1O1Ixp25_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_28),
.B(n_27),
.C(n_26),
.D(n_25),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_146),
.C(n_161),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_165),
.C(n_168),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_140),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_178)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_11),
.B1(n_12),
.B2(n_16),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_179),
.A2(n_184),
.B1(n_150),
.B2(n_156),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_16),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_154),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_194),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_177),
.B(n_160),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_178),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_191),
.B(n_184),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_144),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_166),
.B(n_182),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_204),
.C(n_205),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_185),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_201),
.Y(n_210)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_180),
.B1(n_172),
.B2(n_164),
.Y(n_202)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_202),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_SL g211 ( 
.A(n_203),
.B(n_195),
.C(n_183),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_169),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_202),
.B(n_187),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_211),
.B(n_176),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_190),
.C(n_188),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_179),
.C(n_175),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_197),
.B(n_205),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_215),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_189),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_214),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_210),
.Y(n_218)
);

AOI221xp5_ASAP7_75t_L g219 ( 
.A1(n_218),
.A2(n_216),
.B1(n_208),
.B2(n_171),
.C(n_24),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_219),
.A2(n_18),
.B(n_19),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_20),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_21),
.C(n_200),
.Y(n_222)
);


endmodule