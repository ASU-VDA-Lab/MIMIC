module real_aes_17599_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g119 ( .A(n_0), .B(n_120), .Y(n_119) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_1), .A2(n_3), .B1(n_188), .B2(n_513), .Y(n_512) );
OAI22x1_ASAP7_75t_R g124 ( .A1(n_2), .A2(n_46), .B1(n_125), .B2(n_126), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_2), .Y(n_125) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_4), .A2(n_44), .B1(n_145), .B2(n_168), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_5), .A2(n_27), .B1(n_168), .B2(n_244), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_6), .A2(n_16), .B1(n_187), .B2(n_223), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_7), .A2(n_62), .B1(n_205), .B2(n_246), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_8), .A2(n_17), .B1(n_144), .B2(n_145), .Y(n_529) );
INVx1_ASAP7_75t_L g120 ( .A(n_9), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_10), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_11), .Y(n_143) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_12), .A2(n_19), .B1(n_204), .B2(n_207), .Y(n_203) );
OR2x2_ASAP7_75t_L g110 ( .A(n_13), .B(n_40), .Y(n_110) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_14), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_15), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_18), .A2(n_26), .B1(n_842), .B2(n_846), .Y(n_841) );
INVx2_ASAP7_75t_L g831 ( .A(n_20), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g839 ( .A(n_21), .Y(n_839) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_22), .A2(n_101), .B1(n_187), .B2(n_188), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_23), .A2(n_41), .B1(n_153), .B2(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_24), .B(n_148), .Y(n_147) );
OAI21x1_ASAP7_75t_L g139 ( .A1(n_25), .A2(n_58), .B(n_140), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_26), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_26), .A2(n_79), .B1(n_492), .B2(n_819), .Y(n_818) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_28), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_29), .B(n_150), .Y(n_499) );
INVx4_ASAP7_75t_R g541 ( .A(n_30), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_31), .A2(n_49), .B1(n_173), .B2(n_174), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_32), .A2(n_55), .B1(n_174), .B2(n_187), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_33), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_34), .B(n_153), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_35), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_36), .B(n_168), .Y(n_506) );
INVx1_ASAP7_75t_L g515 ( .A(n_37), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_SL g581 ( .A1(n_38), .A2(n_145), .B(n_149), .C(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_39), .A2(n_56), .B1(n_145), .B2(n_174), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_42), .A2(n_89), .B1(n_145), .B2(n_243), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_43), .A2(n_48), .B1(n_144), .B2(n_145), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_45), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_46), .Y(n_126) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_47), .A2(n_61), .B1(n_187), .B2(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g503 ( .A(n_50), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_51), .B(n_145), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_52), .Y(n_562) );
INVx2_ASAP7_75t_L g118 ( .A(n_53), .Y(n_118) );
BUFx3_ASAP7_75t_L g109 ( .A(n_54), .Y(n_109) );
INVx1_ASAP7_75t_L g826 ( .A(n_54), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_57), .A2(n_90), .B1(n_145), .B2(n_174), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_59), .Y(n_542) );
AOI22x1_ASAP7_75t_SL g803 ( .A1(n_60), .A2(n_69), .B1(n_804), .B2(n_805), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_60), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_63), .A2(n_77), .B1(n_173), .B2(n_191), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_64), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_65), .A2(n_80), .B1(n_144), .B2(n_145), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_66), .A2(n_99), .B1(n_187), .B2(n_207), .Y(n_233) );
INVx1_ASAP7_75t_L g140 ( .A(n_67), .Y(n_140) );
AND2x4_ASAP7_75t_L g159 ( .A(n_68), .B(n_160), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_69), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_70), .A2(n_830), .B1(n_831), .B2(n_832), .Y(n_829) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_70), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_71), .A2(n_92), .B1(n_173), .B2(n_174), .Y(n_511) );
AO22x1_ASAP7_75t_L g520 ( .A1(n_72), .A2(n_78), .B1(n_220), .B2(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g160 ( .A(n_73), .Y(n_160) );
AND2x2_ASAP7_75t_L g584 ( .A(n_74), .B(n_162), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_75), .B(n_246), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_76), .Y(n_577) );
CKINVDCx16_ASAP7_75t_R g819 ( .A(n_79), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_81), .B(n_168), .Y(n_563) );
INVx2_ASAP7_75t_L g150 ( .A(n_82), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_83), .B(n_162), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_84), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_85), .A2(n_100), .B1(n_174), .B2(n_246), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_86), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_87), .B(n_195), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g177 ( .A(n_88), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_91), .B(n_162), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_93), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_94), .B(n_162), .Y(n_559) );
INVx1_ASAP7_75t_L g114 ( .A(n_95), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_95), .B(n_825), .Y(n_824) );
NAND2xp33_ASAP7_75t_L g155 ( .A(n_96), .B(n_148), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g536 ( .A1(n_97), .A2(n_210), .B(n_246), .C(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g543 ( .A(n_98), .B(n_544), .Y(n_543) );
NAND2xp33_ASAP7_75t_L g567 ( .A(n_102), .B(n_154), .Y(n_567) );
AOI21xp33_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_121), .B(n_808), .Y(n_103) );
INVx4_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx4f_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_111), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g112 ( .A(n_108), .B(n_113), .Y(n_112) );
NOR2x1_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g827 ( .A(n_110), .Y(n_827) );
OR2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_115), .Y(n_111) );
AND2x2_ASAP7_75t_L g842 ( .A(n_112), .B(n_843), .Y(n_842) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_113), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g802 ( .A(n_113), .Y(n_802) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_115), .B(n_844), .Y(n_843) );
NAND2xp5_ASAP7_75t_SL g115 ( .A(n_116), .B(n_119), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_117), .B(n_814), .Y(n_813) );
INVx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g847 ( .A(n_118), .B(n_848), .Y(n_847) );
INVx2_ASAP7_75t_SL g815 ( .A(n_119), .Y(n_815) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_803), .B1(n_806), .B2(n_807), .Y(n_122) );
INVx2_ASAP7_75t_L g806 ( .A(n_123), .Y(n_806) );
XNOR2x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_127), .Y(n_123) );
AOI22x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_474), .B1(n_476), .B2(n_800), .Y(n_127) );
XNOR2x1_ASAP7_75t_SL g828 ( .A(n_128), .B(n_829), .Y(n_828) );
NAND2x1p5_ASAP7_75t_L g128 ( .A(n_129), .B(n_418), .Y(n_128) );
NOR3x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_336), .C(n_373), .Y(n_129) );
NAND4xp75_ASAP7_75t_L g130 ( .A(n_131), .B(n_256), .C(n_290), .D(n_320), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OAI32xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_178), .A3(n_228), .B1(n_237), .B2(n_251), .Y(n_132) );
OR2x2_ASAP7_75t_L g237 ( .A(n_133), .B(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_134), .A2(n_448), .B(n_450), .Y(n_447) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_163), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_135), .B(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g319 ( .A(n_135), .B(n_265), .Y(n_319) );
AND2x2_ASAP7_75t_L g414 ( .A(n_135), .B(n_230), .Y(n_414) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx2_ASAP7_75t_L g263 ( .A(n_136), .Y(n_263) );
OAI21x1_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_141), .B(n_161), .Y(n_136) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_137), .A2(n_141), .B(n_161), .Y(n_296) );
INVx2_ASAP7_75t_SL g137 ( .A(n_138), .Y(n_137) );
INVx4_ASAP7_75t_L g162 ( .A(n_138), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_138), .B(n_177), .Y(n_176) );
BUFx3_ASAP7_75t_L g225 ( .A(n_138), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_138), .B(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_138), .B(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g507 ( .A(n_138), .B(n_490), .Y(n_507) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g195 ( .A(n_139), .Y(n_195) );
OAI21x1_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_151), .B(n_157), .Y(n_141) );
O2A1O1Ixp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_147), .C(n_149), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_L g561 ( .A1(n_144), .A2(n_562), .B(n_563), .C(n_564), .Y(n_561) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g191 ( .A(n_145), .Y(n_191) );
INVx1_ASAP7_75t_L g207 ( .A(n_145), .Y(n_207) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_146), .Y(n_148) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_146), .Y(n_168) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
INVx1_ASAP7_75t_L g189 ( .A(n_146), .Y(n_189) );
INVx1_ASAP7_75t_L g206 ( .A(n_146), .Y(n_206) );
INVx1_ASAP7_75t_L g221 ( .A(n_146), .Y(n_221) );
INVx1_ASAP7_75t_L g224 ( .A(n_146), .Y(n_224) );
INVx2_ASAP7_75t_L g244 ( .A(n_146), .Y(n_244) );
INVx1_ASAP7_75t_L g246 ( .A(n_146), .Y(n_246) );
INVx3_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
INVxp67_ASAP7_75t_SL g521 ( .A(n_148), .Y(n_521) );
INVx6_ASAP7_75t_L g156 ( .A(n_149), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_149), .A2(n_520), .B(n_522), .C(n_525), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_149), .A2(n_567), .B(n_568), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_149), .B(n_520), .Y(n_593) );
BUFx8_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g171 ( .A(n_150), .Y(n_171) );
INVx1_ASAP7_75t_L g210 ( .A(n_150), .Y(n_210) );
INVx1_ASAP7_75t_L g502 ( .A(n_150), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_155), .B(n_156), .Y(n_151) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g173 ( .A(n_154), .Y(n_173) );
OAI22xp33_ASAP7_75t_L g540 ( .A1(n_154), .A2(n_224), .B1(n_541), .B2(n_542), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g166 ( .A1(n_156), .A2(n_167), .B1(n_169), .B2(n_172), .Y(n_166) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_156), .A2(n_169), .B1(n_186), .B2(n_190), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_156), .A2(n_203), .B1(n_208), .B2(n_209), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_156), .A2(n_169), .B1(n_219), .B2(n_222), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_156), .A2(n_209), .B1(n_233), .B2(n_234), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_156), .A2(n_242), .B1(n_245), .B2(n_247), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_156), .A2(n_169), .B1(n_281), .B2(n_282), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_156), .A2(n_487), .B1(n_488), .B2(n_489), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_156), .A2(n_247), .B1(n_511), .B2(n_512), .Y(n_510) );
OAI22x1_ASAP7_75t_L g528 ( .A1(n_156), .A2(n_247), .B1(n_529), .B2(n_530), .Y(n_528) );
INVx2_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_SL g248 ( .A(n_158), .Y(n_248) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx10_ASAP7_75t_L g165 ( .A(n_159), .Y(n_165) );
BUFx10_ASAP7_75t_L g490 ( .A(n_159), .Y(n_490) );
INVx1_ASAP7_75t_L g526 ( .A(n_159), .Y(n_526) );
INVx2_ASAP7_75t_L g175 ( .A(n_162), .Y(n_175) );
NOR2x1_ASAP7_75t_L g569 ( .A(n_162), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g287 ( .A(n_163), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_163), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_164), .Y(n_274) );
INVx1_ASAP7_75t_L g318 ( .A(n_164), .Y(n_318) );
AND2x2_ASAP7_75t_L g362 ( .A(n_164), .B(n_296), .Y(n_362) );
OR2x2_ASAP7_75t_L g416 ( .A(n_164), .B(n_240), .Y(n_416) );
AO31x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .A3(n_175), .B(n_176), .Y(n_164) );
INVx2_ASAP7_75t_L g184 ( .A(n_165), .Y(n_184) );
AO31x2_ASAP7_75t_L g201 ( .A1(n_165), .A2(n_202), .A3(n_211), .B(n_213), .Y(n_201) );
AO31x2_ASAP7_75t_L g217 ( .A1(n_165), .A2(n_218), .A3(n_225), .B(n_226), .Y(n_217) );
AO31x2_ASAP7_75t_L g527 ( .A1(n_165), .A2(n_198), .A3(n_528), .B(n_531), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_168), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g489 ( .A(n_170), .Y(n_489) );
BUFx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g565 ( .A(n_171), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_174), .B(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g513 ( .A(n_174), .Y(n_513) );
AO31x2_ASAP7_75t_L g485 ( .A1(n_175), .A2(n_486), .A3(n_490), .B(n_491), .Y(n_485) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_179), .A2(n_342), .B1(n_434), .B2(n_436), .Y(n_433) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_199), .Y(n_179) );
INVx4_ASAP7_75t_L g259 ( .A(n_180), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_180), .A2(n_239), .B1(n_271), .B2(n_273), .Y(n_270) );
OR2x2_ASAP7_75t_L g276 ( .A(n_180), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g395 ( .A(n_180), .B(n_294), .Y(n_395) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g315 ( .A(n_181), .B(n_200), .Y(n_315) );
AND2x2_ASAP7_75t_L g406 ( .A(n_181), .B(n_278), .Y(n_406) );
AND2x2_ASAP7_75t_L g461 ( .A(n_181), .B(n_217), .Y(n_461) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g255 ( .A(n_182), .Y(n_255) );
AND2x4_ASAP7_75t_L g382 ( .A(n_182), .B(n_278), .Y(n_382) );
AO31x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_185), .A3(n_192), .B(n_196), .Y(n_182) );
AO31x2_ASAP7_75t_L g231 ( .A1(n_183), .A2(n_211), .A3(n_232), .B(n_235), .Y(n_231) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_184), .A2(n_536), .B(n_539), .Y(n_535) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_189), .B(n_579), .Y(n_578) );
AO31x2_ASAP7_75t_L g279 ( .A1(n_192), .A2(n_248), .A3(n_280), .B(n_283), .Y(n_279) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_192), .A2(n_535), .B(n_543), .Y(n_534) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_SL g213 ( .A(n_194), .B(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_194), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g198 ( .A(n_195), .Y(n_198) );
INVx2_ASAP7_75t_L g212 ( .A(n_195), .Y(n_212) );
OAI21xp33_ASAP7_75t_L g525 ( .A1(n_195), .A2(n_524), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_198), .B(n_284), .Y(n_283) );
NAND2x1_ASAP7_75t_L g258 ( .A(n_199), .B(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_199), .B(n_366), .Y(n_365) );
AND2x4_ASAP7_75t_L g199 ( .A(n_200), .B(n_215), .Y(n_199) );
INVx2_ASAP7_75t_L g253 ( .A(n_200), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_200), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g301 ( .A(n_200), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_200), .B(n_303), .Y(n_328) );
AND2x2_ASAP7_75t_L g331 ( .A(n_200), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g391 ( .A(n_200), .Y(n_391) );
INVx4_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_201), .B(n_216), .Y(n_269) );
BUFx2_ASAP7_75t_L g307 ( .A(n_201), .Y(n_307) );
AND2x2_ASAP7_75t_L g356 ( .A(n_201), .B(n_217), .Y(n_356) );
AND2x2_ASAP7_75t_L g398 ( .A(n_201), .B(n_279), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_201), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_206), .B(n_538), .Y(n_537) );
INVx1_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g247 ( .A(n_210), .Y(n_247) );
AO31x2_ASAP7_75t_L g509 ( .A1(n_211), .A2(n_248), .A3(n_510), .B(n_514), .Y(n_509) );
AOI21x1_ASAP7_75t_L g573 ( .A1(n_211), .A2(n_574), .B(n_584), .Y(n_573) );
BUFx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_212), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_212), .B(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_212), .B(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g544 ( .A(n_212), .Y(n_544) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_217), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g309 ( .A(n_217), .B(n_279), .Y(n_309) );
INVx1_ASAP7_75t_L g332 ( .A(n_217), .Y(n_332) );
INVx2_ASAP7_75t_L g352 ( .A(n_217), .Y(n_352) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_217), .Y(n_397) );
OAI21xp33_ASAP7_75t_SL g498 ( .A1(n_220), .A2(n_499), .B(n_500), .Y(n_498) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AO31x2_ASAP7_75t_L g240 ( .A1(n_225), .A2(n_241), .A3(n_248), .B(n_249), .Y(n_240) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g316 ( .A(n_229), .B(n_317), .Y(n_316) );
NOR2x1p5_ASAP7_75t_L g422 ( .A(n_229), .B(n_416), .Y(n_422) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x4_ASAP7_75t_L g239 ( .A(n_230), .B(n_240), .Y(n_239) );
INVx3_ASAP7_75t_L g272 ( .A(n_230), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_230), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_230), .B(n_348), .Y(n_347) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g264 ( .A(n_231), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g322 ( .A(n_231), .B(n_240), .Y(n_322) );
BUFx2_ASAP7_75t_L g435 ( .A(n_231), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_237), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g473 ( .A(n_237), .Y(n_473) );
INVx2_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g409 ( .A(n_239), .Y(n_409) );
AND2x4_ASAP7_75t_L g432 ( .A(n_239), .B(n_362), .Y(n_432) );
AND2x2_ASAP7_75t_L g456 ( .A(n_239), .B(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g265 ( .A(n_240), .Y(n_265) );
BUFx2_ASAP7_75t_L g289 ( .A(n_240), .Y(n_289) );
INVx1_ASAP7_75t_L g345 ( .A(n_240), .Y(n_345) );
OR2x2_ASAP7_75t_L g467 ( .A(n_240), .B(n_324), .Y(n_467) );
INVx2_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_244), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_247), .B(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
INVx2_ASAP7_75t_L g313 ( .A(n_253), .Y(n_313) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_254), .Y(n_330) );
INVx1_ASAP7_75t_L g334 ( .A(n_254), .Y(n_334) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g275 ( .A(n_255), .Y(n_275) );
OR2x2_ASAP7_75t_L g312 ( .A(n_255), .B(n_304), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_260), .B(n_266), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_261), .A2(n_355), .B1(n_357), .B2(n_360), .Y(n_354) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
OR2x2_ASAP7_75t_L g400 ( .A(n_263), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g408 ( .A(n_263), .Y(n_408) );
AND2x2_ASAP7_75t_L g421 ( .A(n_263), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g383 ( .A(n_264), .B(n_362), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_270), .B1(n_276), .B2(n_285), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g335 ( .A(n_269), .Y(n_335) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x4_ASAP7_75t_L g293 ( .A(n_272), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g361 ( .A(n_272), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g370 ( .A(n_272), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_272), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_273), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AND2x2_ASAP7_75t_L g358 ( .A(n_275), .B(n_359), .Y(n_358) );
INVx3_ASAP7_75t_L g372 ( .A(n_275), .Y(n_372) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g304 ( .A(n_279), .Y(n_304) );
AND2x4_ASAP7_75t_L g351 ( .A(n_279), .B(n_352), .Y(n_351) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_279), .Y(n_367) );
INVx1_ASAP7_75t_L g431 ( .A(n_279), .Y(n_431) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
AND2x4_ASAP7_75t_L g323 ( .A(n_287), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g340 ( .A(n_287), .Y(n_340) );
INVx1_ASAP7_75t_L g298 ( .A(n_289), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_299), .B1(n_310), .B2(n_316), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2x1p5_ASAP7_75t_L g292 ( .A(n_293), .B(n_297), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVxp67_ASAP7_75t_SL g348 ( .A(n_295), .Y(n_348) );
INVx1_ASAP7_75t_L g324 ( .A(n_296), .Y(n_324) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_300), .B(n_305), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_301), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g453 ( .A(n_302), .Y(n_453) );
INVx1_ASAP7_75t_L g472 ( .A(n_302), .Y(n_472) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2x1_ASAP7_75t_L g449 ( .A(n_306), .B(n_372), .Y(n_449) );
AND2x4_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g465 ( .A(n_307), .Y(n_465) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
INVx2_ASAP7_75t_L g403 ( .A(n_311), .Y(n_403) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx2_ASAP7_75t_L g392 ( .A(n_312), .Y(n_392) );
AND2x4_ASAP7_75t_L g394 ( .A(n_313), .B(n_351), .Y(n_394) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_317), .A2(n_463), .B1(n_466), .B2(n_468), .Y(n_462) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_L g387 ( .A(n_318), .Y(n_387) );
INVx1_ASAP7_75t_L g341 ( .A(n_319), .Y(n_341) );
AND2x4_ASAP7_75t_L g434 ( .A(n_319), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g442 ( .A(n_319), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_325), .Y(n_320) );
AND2x4_ASAP7_75t_SL g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_SL g385 ( .A(n_322), .Y(n_385) );
INVx2_ASAP7_75t_L g401 ( .A(n_322), .Y(n_401) );
INVx1_ASAP7_75t_L g428 ( .A(n_323), .Y(n_428) );
AND2x2_ASAP7_75t_L g459 ( .A(n_323), .B(n_370), .Y(n_459) );
NAND3xp33_ASAP7_75t_L g325 ( .A(n_326), .B(n_329), .C(n_333), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_330), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g371 ( .A(n_331), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_331), .B(n_406), .Y(n_439) );
INVx1_ASAP7_75t_L g359 ( .A(n_332), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_334), .B(n_398), .Y(n_424) );
INVx1_ASAP7_75t_L g379 ( .A(n_335), .Y(n_379) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_353), .C(n_363), .Y(n_336) );
OAI21xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_342), .B(n_349), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g457 ( .A(n_340), .Y(n_457) );
AND2x4_ASAP7_75t_L g342 ( .A(n_343), .B(n_346), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI32xp33_ASAP7_75t_L g393 ( .A1(n_344), .A2(n_394), .A3(n_395), .B1(n_396), .B2(n_399), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_344), .B(n_428), .Y(n_427) );
BUFx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g377 ( .A(n_351), .Y(n_377) );
NAND2x1p5_ASAP7_75t_L g412 ( .A(n_351), .B(n_372), .Y(n_412) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_356), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g417 ( .A(n_356), .B(n_366), .Y(n_417) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g445 ( .A(n_359), .Y(n_445) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
AOI22xp33_ASAP7_75t_SL g363 ( .A1(n_361), .A2(n_364), .B1(n_368), .B2(n_371), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_362), .B(n_370), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_364), .A2(n_422), .B1(n_459), .B2(n_460), .Y(n_458) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g460 ( .A(n_366), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_368), .A2(n_411), .B1(n_413), .B2(n_417), .Y(n_410) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g452 ( .A(n_372), .Y(n_452) );
NAND4xp25_ASAP7_75t_L g373 ( .A(n_374), .B(n_393), .C(n_402), .D(n_410), .Y(n_373) );
O2A1O1Ixp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_380), .B(n_383), .C(n_384), .Y(n_374) );
NOR2x1_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_L g438 ( .A(n_382), .B(n_397), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_382), .B(n_465), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B(n_388), .Y(n_384) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_389), .A2(n_427), .B1(n_429), .B2(n_432), .Y(n_426) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_394), .A2(n_399), .B(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI21xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B(n_407), .Y(n_402) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_R g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_417), .A2(n_434), .B1(n_471), .B2(n_473), .Y(n_470) );
NOR3x1_ASAP7_75t_L g418 ( .A(n_419), .B(n_440), .C(n_454), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_433), .Y(n_419) );
AOI21xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B(n_425), .Y(n_420) );
INVx1_ASAP7_75t_L g446 ( .A(n_421), .Y(n_446) );
INVx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g469 ( .A(n_431), .Y(n_469) );
INVx1_ASAP7_75t_L g443 ( .A(n_435), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
OAI221xp5_ASAP7_75t_L g440 ( .A1(n_437), .A2(n_441), .B1(n_444), .B2(n_446), .C(n_447), .Y(n_440) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
NAND4xp25_ASAP7_75t_SL g454 ( .A(n_455), .B(n_458), .C(n_462), .D(n_470), .Y(n_454) );
AND2x2_ASAP7_75t_L g468 ( .A(n_461), .B(n_469), .Y(n_468) );
INVxp67_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
INVxp67_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_478), .B(n_677), .Y(n_477) );
NOR2x1_ASAP7_75t_L g478 ( .A(n_479), .B(n_625), .Y(n_478) );
OAI211xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_516), .B(n_545), .C(n_610), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g760 ( .A1(n_482), .A2(n_546), .B(n_761), .Y(n_760) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_493), .Y(n_482) );
INVx2_ASAP7_75t_L g606 ( .A(n_483), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_483), .B(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g717 ( .A(n_484), .B(n_495), .Y(n_717) );
BUFx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_SL g585 ( .A(n_485), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_485), .B(n_509), .Y(n_622) );
AND2x2_ASAP7_75t_L g655 ( .A(n_485), .B(n_572), .Y(n_655) );
OR2x2_ASAP7_75t_L g660 ( .A(n_485), .B(n_509), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_489), .A2(n_505), .B(n_506), .Y(n_504) );
OAI21x1_ASAP7_75t_L g522 ( .A1(n_489), .A2(n_523), .B(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g570 ( .A(n_490), .Y(n_570) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g799 ( .A(n_494), .Y(n_799) );
OR2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_508), .Y(n_494) );
AND2x2_ASAP7_75t_L g600 ( .A(n_495), .B(n_509), .Y(n_600) );
INVx3_ASAP7_75t_L g608 ( .A(n_495), .Y(n_608) );
NAND2x1p5_ASAP7_75t_SL g640 ( .A(n_495), .B(n_624), .Y(n_640) );
INVx1_ASAP7_75t_L g658 ( .A(n_495), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_495), .B(n_603), .Y(n_683) );
BUFx2_ASAP7_75t_L g769 ( .A(n_495), .Y(n_769) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_504), .B(n_507), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
BUFx4f_ASAP7_75t_L g580 ( .A(n_502), .Y(n_580) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g553 ( .A(n_509), .Y(n_553) );
INVx1_ASAP7_75t_L g609 ( .A(n_509), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_509), .B(n_585), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_509), .B(n_572), .Y(n_718) );
OR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_533), .Y(n_516) );
INVx1_ASAP7_75t_L g776 ( .A(n_517), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_527), .Y(n_517) );
OR2x2_ASAP7_75t_L g548 ( .A(n_518), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g613 ( .A(n_518), .Y(n_613) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g592 ( .A(n_522), .Y(n_592) );
INVx1_ASAP7_75t_L g594 ( .A(n_525), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_526), .A2(n_575), .B(n_581), .Y(n_574) );
INVx2_ASAP7_75t_L g549 ( .A(n_527), .Y(n_549) );
OR2x2_ASAP7_75t_L g614 ( .A(n_527), .B(n_534), .Y(n_614) );
AND2x2_ASAP7_75t_L g619 ( .A(n_527), .B(n_534), .Y(n_619) );
INVx2_ASAP7_75t_L g664 ( .A(n_527), .Y(n_664) );
AND2x2_ASAP7_75t_L g705 ( .A(n_527), .B(n_558), .Y(n_705) );
AND2x2_ASAP7_75t_L g739 ( .A(n_527), .B(n_636), .Y(n_739) );
INVx1_ASAP7_75t_L g550 ( .A(n_533), .Y(n_550) );
INVx1_ASAP7_75t_L g669 ( .A(n_533), .Y(n_669) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g589 ( .A(n_534), .B(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g630 ( .A(n_534), .B(n_591), .Y(n_630) );
INVx2_ASAP7_75t_L g636 ( .A(n_534), .Y(n_636) );
AND2x2_ASAP7_75t_L g691 ( .A(n_534), .B(n_558), .Y(n_691) );
AND2x2_ASAP7_75t_L g748 ( .A(n_534), .B(n_557), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_551), .B1(n_586), .B2(n_597), .Y(n_545) );
INVx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
NAND3xp33_ASAP7_75t_SL g726 ( .A(n_548), .B(n_727), .C(n_729), .Y(n_726) );
INVx1_ASAP7_75t_L g645 ( .A(n_549), .Y(n_645) );
AND2x2_ASAP7_75t_L g695 ( .A(n_549), .B(n_557), .Y(n_695) );
INVx1_ASAP7_75t_L g795 ( .A(n_550), .Y(n_795) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_554), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_552), .B(n_750), .Y(n_786) );
BUFx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g641 ( .A(n_553), .Y(n_641) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_571), .Y(n_555) );
INVx1_ASAP7_75t_L g629 ( .A(n_556), .Y(n_629) );
BUFx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g709 ( .A(n_557), .B(n_590), .Y(n_709) );
AND2x2_ASAP7_75t_L g728 ( .A(n_557), .B(n_635), .Y(n_728) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g596 ( .A(n_558), .Y(n_596) );
BUFx3_ASAP7_75t_L g634 ( .A(n_558), .Y(n_634) );
AND2x2_ASAP7_75t_L g663 ( .A(n_558), .B(n_664), .Y(n_663) );
NAND2x1p5_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
OAI21x1_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_566), .B(n_569), .Y(n_560) );
INVx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g756 ( .A(n_571), .Y(n_756) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_585), .Y(n_571) );
INVx2_ASAP7_75t_L g624 ( .A(n_572), .Y(n_624) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g603 ( .A(n_573), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_578), .B(n_580), .Y(n_575) );
INVx1_ASAP7_75t_L g604 ( .A(n_585), .Y(n_604) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x6_ASAP7_75t_L g587 ( .A(n_588), .B(n_595), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g643 ( .A(n_589), .B(n_644), .Y(n_643) );
BUFx2_ASAP7_75t_L g773 ( .A(n_589), .Y(n_773) );
INVx1_ASAP7_75t_L g618 ( .A(n_590), .Y(n_618) );
AND2x2_ASAP7_75t_L g698 ( .A(n_590), .B(n_636), .Y(n_698) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g635 ( .A(n_591), .B(n_636), .Y(n_635) );
AOI21x1_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B(n_594), .Y(n_591) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NOR2x1_ASAP7_75t_L g647 ( .A(n_596), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g731 ( .A(n_596), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_605), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_598), .A2(n_639), .B1(n_642), .B2(n_646), .Y(n_638) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_599), .A2(n_619), .B1(n_651), .B2(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
BUFx2_ASAP7_75t_SL g637 ( .A(n_600), .Y(n_637) );
AND2x4_ASAP7_75t_L g755 ( .A(n_600), .B(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g764 ( .A(n_600), .Y(n_764) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g676 ( .A(n_602), .Y(n_676) );
OR2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_603), .B(n_608), .Y(n_734) );
INVxp67_ASAP7_75t_L g763 ( .A(n_603), .Y(n_763) );
AND2x2_ASAP7_75t_L g768 ( .A(n_603), .B(n_634), .Y(n_768) );
OR2x2_ASAP7_75t_L g750 ( .A(n_604), .B(n_624), .Y(n_750) );
INVx1_ASAP7_75t_L g631 ( .A(n_605), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_606), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g670 ( .A(n_607), .B(n_655), .Y(n_670) );
AND2x4_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_608), .B(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g654 ( .A(n_608), .Y(n_654) );
OR2x2_ASAP7_75t_L g749 ( .A(n_608), .B(n_750), .Y(n_749) );
OAI21xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_615), .B(n_620), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g673 ( .A(n_612), .Y(n_673) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g667 ( .A(n_613), .B(n_664), .Y(n_667) );
INVx2_ASAP7_75t_L g791 ( .A(n_613), .Y(n_791) );
INVx2_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
AND2x2_ASAP7_75t_L g720 ( .A(n_617), .B(n_663), .Y(n_720) );
AND2x2_ASAP7_75t_L g745 ( .A(n_617), .B(n_691), .Y(n_745) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g648 ( .A(n_618), .Y(n_648) );
AND2x2_ASAP7_75t_L g675 ( .A(n_619), .B(n_629), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_619), .B(n_674), .Y(n_687) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g772 ( .A(n_622), .Y(n_772) );
OR2x2_ASAP7_75t_L g788 ( .A(n_622), .B(n_683), .Y(n_788) );
INVx1_ASAP7_75t_L g712 ( .A(n_624), .Y(n_712) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_649), .C(n_671), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_631), .B1(n_632), .B2(n_637), .C(n_638), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
AND2x2_ASAP7_75t_L g651 ( .A(n_630), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_630), .B(n_695), .Y(n_779) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
BUFx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx3_ASAP7_75t_L g674 ( .A(n_634), .Y(n_674) );
AND3x1_ASAP7_75t_L g770 ( .A(n_634), .B(n_771), .C(n_772), .Y(n_770) );
AND2x2_ASAP7_75t_L g757 ( .A(n_635), .B(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g767 ( .A(n_635), .Y(n_767) );
INVxp67_ASAP7_75t_L g781 ( .A(n_637), .Y(n_781) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
OR2x2_ASAP7_75t_L g736 ( .A(n_640), .B(n_660), .Y(n_736) );
INVx2_ASAP7_75t_L g771 ( .A(n_640), .Y(n_771) );
INVx1_ASAP7_75t_L g689 ( .A(n_641), .Y(n_689) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g690 ( .A1(n_643), .A2(n_691), .B(n_692), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_644), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g652 ( .A(n_645), .Y(n_652) );
OR2x2_ASAP7_75t_L g746 ( .A(n_645), .B(n_747), .Y(n_746) );
INVxp67_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g706 ( .A(n_648), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_648), .B(n_705), .Y(n_785) );
AND3x1_ASAP7_75t_L g649 ( .A(n_650), .B(n_656), .C(n_661), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
AND2x2_ASAP7_75t_L g700 ( .A(n_652), .B(n_691), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_653), .A2(n_720), .B1(n_721), .B2(n_723), .Y(n_719) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
OAI321xp33_ASAP7_75t_L g742 ( .A1(n_654), .A2(n_743), .A3(n_744), .B1(n_746), .B2(n_749), .C(n_751), .Y(n_742) );
AND2x2_ASAP7_75t_L g794 ( .A(n_654), .B(n_659), .Y(n_794) );
AND2x2_ASAP7_75t_L g692 ( .A(n_655), .B(n_658), .Y(n_692) );
INVx2_ASAP7_75t_L g701 ( .A(n_657), .Y(n_701) );
AND2x2_ASAP7_75t_L g710 ( .A(n_657), .B(n_711), .Y(n_710) );
AND2x4_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g722 ( .A(n_660), .B(n_712), .Y(n_722) );
INVx2_ASAP7_75t_L g754 ( .A(n_660), .Y(n_754) );
OAI21xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_665), .B(n_670), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g758 ( .A(n_664), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_666), .B(n_668), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2x1p5_ASAP7_75t_L g684 ( .A(n_667), .B(n_674), .Y(n_684) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OAI21xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_675), .B(n_676), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_674), .B(n_698), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_674), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g775 ( .A(n_674), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g743 ( .A(n_676), .Y(n_743) );
NOR2xp67_ASAP7_75t_L g677 ( .A(n_678), .B(n_740), .Y(n_677) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_702), .C(n_725), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_693), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_684), .B1(n_685), .B2(n_688), .C(n_690), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
OR2x2_ASAP7_75t_L g733 ( .A(n_682), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI21xp33_ASAP7_75t_SL g693 ( .A1(n_694), .A2(n_699), .B(n_701), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g730 ( .A(n_698), .B(n_731), .Y(n_730) );
OAI21xp33_ASAP7_75t_SL g713 ( .A1(n_699), .A2(n_714), .B(n_719), .Y(n_713) );
INVx2_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_707), .B(n_710), .C(n_713), .Y(n_702) );
INVx2_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_704), .B(n_779), .Y(n_778) );
NAND2x1_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_712), .B(n_754), .Y(n_753) );
INVxp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g774 ( .A(n_715), .B(n_775), .Y(n_774) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_732), .B1(n_735), .B2(n_737), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
HB1xp67_ASAP7_75t_L g797 ( .A(n_734), .Y(n_797) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_777), .C(n_792), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_759), .Y(n_741) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
OAI21xp33_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_755), .B(n_757), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_765), .C(n_774), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
OR2x2_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
AOI32xp33_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_768), .A3(n_769), .B1(n_770), .B2(n_773), .Y(n_765) );
INVx3_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
AND2x2_ASAP7_75t_L g793 ( .A(n_768), .B(n_794), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_780), .B(n_782), .Y(n_777) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AOI22x1_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_786), .B1(n_787), .B2(n_789), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AOI21xp33_ASAP7_75t_L g796 ( .A1(n_785), .A2(n_797), .B(n_798), .Y(n_796) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_795), .B(n_796), .Y(n_792) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx8_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
BUFx12f_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_SL g807 ( .A(n_803), .Y(n_807) );
OAI21xp33_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_816), .B(n_841), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
INVx4_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
BUFx3_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
OR2x4_ASAP7_75t_L g846 ( .A(n_814), .B(n_847), .Y(n_846) );
BUFx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_820), .B(n_833), .Y(n_817) );
OAI31xp33_ASAP7_75t_SL g833 ( .A1(n_818), .A2(n_828), .A3(n_834), .B(n_837), .Y(n_833) );
AND2x2_ASAP7_75t_L g820 ( .A(n_821), .B(n_828), .Y(n_820) );
BUFx12f_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx4_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx5_ASAP7_75t_L g836 ( .A(n_823), .Y(n_836) );
INVx5_ASAP7_75t_L g840 ( .A(n_823), .Y(n_840) );
CKINVDCx8_ASAP7_75t_R g845 ( .A(n_823), .Y(n_845) );
INVx3_ASAP7_75t_L g848 ( .A(n_823), .Y(n_848) );
AND2x6_ASAP7_75t_SL g823 ( .A(n_824), .B(n_827), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
BUFx3_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVxp67_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
INVx3_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
endmodule