module fake_jpeg_10708_n_134 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_134);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx2_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_57),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_40),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_64),
.Y(n_68)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_0),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_44),
.Y(n_74)
);

FAx1_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_47),
.CI(n_48),
.CON(n_75),
.SN(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_64),
.B(n_58),
.C(n_56),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_48),
.B1(n_53),
.B2(n_49),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_76),
.A2(n_78),
.B1(n_77),
.B2(n_56),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_48),
.B1(n_51),
.B2(n_50),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_82),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_81),
.B(n_1),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_63),
.B(n_55),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_61),
.B1(n_42),
.B2(n_52),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_90),
.B1(n_3),
.B2(n_4),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_78),
.B(n_46),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_88),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_1),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_21),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_20),
.B(n_39),
.C(n_36),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

BUFx4f_ASAP7_75t_SL g95 ( 
.A(n_93),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_99),
.B1(n_104),
.B2(n_100),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_85),
.B(n_2),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_101),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_97),
.B(n_106),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_23),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_17),
.B(n_34),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_14),
.B(n_32),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_4),
.B(n_5),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_5),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_108),
.B(n_9),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_93),
.B1(n_82),
.B2(n_8),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_R g110 ( 
.A1(n_103),
.A2(n_24),
.B(n_33),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_112),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_107),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_104),
.A2(n_25),
.B1(n_30),
.B2(n_10),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_114),
.C(n_116),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_6),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_9),
.Y(n_116)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

AOI321xp33_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_119),
.A3(n_115),
.B1(n_110),
.B2(n_118),
.C(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_125),
.B(n_126),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_113),
.B(n_100),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_95),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_119),
.C(n_120),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_95),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_128),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_121),
.B(n_26),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_12),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_121),
.C(n_28),
.Y(n_134)
);


endmodule