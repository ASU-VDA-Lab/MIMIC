module fake_jpeg_22809_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_46),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_25),
.Y(n_64)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_61),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_9),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_58),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_8),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_8),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_7),
.Y(n_99)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_63),
.A2(n_45),
.B1(n_22),
.B2(n_33),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_64),
.B(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_0),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_73),
.Y(n_84)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_78),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_32),
.B1(n_29),
.B2(n_40),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_75),
.A2(n_88),
.B1(n_98),
.B2(n_16),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_50),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_83),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_82),
.Y(n_128)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_41),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_35),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_39),
.B1(n_46),
.B2(n_45),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_107),
.B1(n_71),
.B2(n_61),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_33),
.B1(n_22),
.B2(n_24),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_90),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_92),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_55),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_56),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_100),
.B(n_106),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_SL g101 ( 
.A1(n_58),
.A2(n_47),
.B(n_37),
.C(n_27),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_110),
.B1(n_111),
.B2(n_68),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_0),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_59),
.A2(n_38),
.B1(n_37),
.B2(n_35),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_109),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_59),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_67),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_0),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_15),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_113),
.A2(n_133),
.B1(n_135),
.B2(n_93),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_31),
.B(n_16),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_118),
.A2(n_123),
.B(n_31),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_120),
.B(n_105),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_35),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_125),
.Y(n_150)
);

NAND2xp33_ASAP7_75t_SL g123 ( 
.A(n_107),
.B(n_1),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_28),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_28),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_127),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_28),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_27),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_129),
.B(n_138),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_142),
.B1(n_84),
.B2(n_103),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_34),
.Y(n_139)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_139),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_98),
.A2(n_52),
.B1(n_18),
.B2(n_17),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_94),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_145),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_87),
.B1(n_52),
.B2(n_101),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_146),
.A2(n_151),
.B1(n_161),
.B2(n_172),
.Y(n_197)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_152),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_87),
.B1(n_111),
.B2(n_104),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_155),
.Y(n_183)
);

AO22x1_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_87),
.B1(n_107),
.B2(n_93),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_154),
.A2(n_169),
.B(n_170),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_76),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_158),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_157),
.B(n_163),
.Y(n_190)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_167),
.B1(n_175),
.B2(n_140),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_83),
.B1(n_84),
.B2(n_107),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_76),
.Y(n_162)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_121),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_86),
.Y(n_164)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_171),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_77),
.Y(n_166)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_135),
.A2(n_100),
.B1(n_95),
.B2(n_99),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_120),
.A2(n_89),
.B1(n_79),
.B2(n_74),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_174),
.A2(n_142),
.B(n_133),
.Y(n_200)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_150),
.B(n_138),
.CI(n_129),
.CON(n_182),
.SN(n_182)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_205),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_168),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_187),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_167),
.A2(n_123),
.B1(n_139),
.B2(n_127),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_186),
.A2(n_203),
.B1(n_153),
.B2(n_152),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_119),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_118),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_201),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_119),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_189),
.B(n_191),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_119),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_131),
.B(n_132),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_194),
.A2(n_200),
.B(n_202),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_195),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_143),
.B(n_133),
.Y(n_198)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_204),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_128),
.C(n_132),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_149),
.A2(n_140),
.B(n_96),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_160),
.A2(n_82),
.B1(n_34),
.B2(n_30),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_154),
.A2(n_34),
.B(n_23),
.C(n_4),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_128),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_206),
.Y(n_211)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_3),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_2),
.Y(n_209)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

OA22x2_ASAP7_75t_L g213 ( 
.A1(n_205),
.A2(n_154),
.B1(n_146),
.B2(n_169),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_213),
.A2(n_194),
.B1(n_201),
.B2(n_203),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_171),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_217),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_204),
.A2(n_147),
.B1(n_144),
.B2(n_156),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_218),
.B1(n_230),
.B2(n_234),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_163),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_186),
.B(n_23),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_188),
.Y(n_251)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_226),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_159),
.B(n_3),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_224),
.A2(n_209),
.B(n_178),
.Y(n_255)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_183),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_229),
.Y(n_244)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_181),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_208),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_232),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_179),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_197),
.A2(n_4),
.B1(n_7),
.B2(n_10),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_197),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_237),
.A2(n_190),
.B1(n_184),
.B2(n_177),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_192),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_247),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_246),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_185),
.C(n_191),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_256),
.C(n_258),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_227),
.A2(n_200),
.B(n_198),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_221),
.B(n_182),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_257),
.Y(n_267)
);

NOR2x1_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_178),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_254),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_250),
.Y(n_274)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_213),
.Y(n_277)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_206),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_254),
.A2(n_255),
.B(n_184),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_182),
.C(n_199),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_224),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_212),
.B(n_176),
.C(n_177),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_190),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_211),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_260),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_239),
.A2(n_222),
.B1(n_210),
.B2(n_227),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_271),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_249),
.Y(n_262)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_264),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_268),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_252),
.A2(n_218),
.B1(n_213),
.B2(n_219),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_270),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_217),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_237),
.B1(n_236),
.B2(n_230),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_277),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_213),
.B1(n_215),
.B2(n_179),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_273),
.B(n_275),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_279),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_244),
.Y(n_275)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_242),
.B(n_193),
.C(n_11),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_247),
.C(n_251),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_258),
.C(n_238),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_292),
.C(n_295),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g283 ( 
.A(n_262),
.B(n_256),
.CI(n_255),
.CON(n_283),
.SN(n_283)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_279),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_284),
.A2(n_292),
.B(n_293),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_250),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_266),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_254),
.C(n_241),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_241),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_241),
.C(n_243),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_270),
.C(n_265),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_298),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_R g298 ( 
.A(n_283),
.B(n_269),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_290),
.Y(n_299)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_300),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_193),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_304),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_303),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_267),
.B(n_264),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_263),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_305),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_282),
.A2(n_261),
.B1(n_273),
.B2(n_272),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_307),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_280),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_308),
.B(n_309),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_10),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_294),
.C(n_295),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_312),
.C(n_294),
.Y(n_320)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_321),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_320),
.B(n_322),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_311),
.C(n_310),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_310),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_315),
.B(n_299),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_306),
.C(n_303),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_284),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_316),
.B(n_289),
.C(n_307),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_326),
.A2(n_323),
.B(n_313),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_331),
.C(n_328),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_289),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_327),
.Y(n_333)
);

OAI321xp33_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C(n_303),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_336),
.Y(n_337)
);


endmodule