module fake_jpeg_4051_n_39 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_39);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_6),
.B(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_17),
.B(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_15),
.B(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_0),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_32),
.B(n_33),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_27),
.B1(n_22),
.B2(n_31),
.Y(n_36)
);

NOR3xp33_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_35),
.C(n_1),
.Y(n_37)
);

AOI322xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_26),
.A3(n_24),
.B1(n_0),
.B2(n_12),
.C1(n_16),
.C2(n_18),
.Y(n_38)
);

OAI221xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_2),
.B1(n_4),
.B2(n_19),
.C(n_27),
.Y(n_39)
);


endmodule