module fake_jpeg_3642_n_450 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_450);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_450;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_SL g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_20),
.B(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_54),
.B(n_76),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_56),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_57),
.Y(n_160)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_58),
.Y(n_114)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_61),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_63),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_64),
.Y(n_169)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_27),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_73),
.Y(n_128)
);

BUFx4f_ASAP7_75t_SL g68 ( 
.A(n_27),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_68),
.Y(n_117)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

BUFx16f_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

BUFx2_ASAP7_75t_R g72 ( 
.A(n_17),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g181 ( 
.A(n_72),
.B(n_103),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_74),
.Y(n_159)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_31),
.B(n_16),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_39),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_77),
.B(n_79),
.Y(n_145)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_39),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_28),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_81),
.B(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_83),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_20),
.B(n_26),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_88),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_33),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_26),
.B(n_15),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_37),
.B(n_15),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_91),
.B(n_94),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_37),
.B(n_12),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_96),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_38),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_97),
.B(n_99),
.Y(n_157)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_38),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_41),
.B(n_30),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_100),
.B(n_101),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_38),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_18),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_18),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_41),
.B(n_10),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_42),
.B(n_9),
.Y(n_111)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_112),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_70),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_121),
.B(n_125),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_70),
.A2(n_35),
.B1(n_42),
.B2(n_46),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_SL g191 ( 
.A1(n_122),
.A2(n_129),
.B(n_130),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_61),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_103),
.A2(n_35),
.B1(n_42),
.B2(n_46),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_58),
.A2(n_22),
.B1(n_21),
.B2(n_49),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_55),
.A2(n_44),
.B1(n_22),
.B2(n_49),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_134),
.A2(n_143),
.B1(n_144),
.B2(n_165),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_72),
.A2(n_22),
.B1(n_48),
.B2(n_49),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_141),
.A2(n_162),
.B1(n_63),
.B2(n_75),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_60),
.B(n_66),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g234 ( 
.A(n_142),
.B(n_161),
.C(n_177),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_71),
.A2(n_44),
.B1(n_48),
.B2(n_51),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_74),
.A2(n_90),
.B1(n_87),
.B2(n_93),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_62),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_153),
.B(n_5),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_95),
.B(n_44),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_108),
.A2(n_51),
.B1(n_50),
.B2(n_45),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_83),
.A2(n_50),
.B1(n_45),
.B2(n_43),
.Y(n_165)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_64),
.Y(n_168)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_96),
.A2(n_43),
.B1(n_34),
.B2(n_30),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_173),
.A2(n_180),
.B1(n_1),
.B2(n_3),
.Y(n_201)
);

INVx5_ASAP7_75t_SL g174 ( 
.A(n_68),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_89),
.B(n_34),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_107),
.B(n_29),
.C(n_24),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_1),
.C(n_3),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_102),
.A2(n_24),
.B1(n_29),
.B2(n_23),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_106),
.A2(n_23),
.B1(n_10),
.B2(n_4),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_1),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_68),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_185),
.B(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_113),
.Y(n_186)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_186),
.Y(n_269)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

O2A1O1Ixp33_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_92),
.B(n_85),
.C(n_112),
.Y(n_192)
);

OA21x2_ASAP7_75t_L g276 ( 
.A1(n_192),
.A2(n_182),
.B(n_169),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_120),
.A2(n_57),
.B1(n_56),
.B2(n_105),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_193),
.A2(n_201),
.B1(n_210),
.B2(n_231),
.Y(n_278)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_194),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_196),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_197),
.A2(n_232),
.B1(n_237),
.B2(n_239),
.Y(n_254)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_198),
.Y(n_264)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_199),
.Y(n_281)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_200),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_202),
.B(n_209),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_203),
.Y(n_282)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_204),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_128),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_205),
.B(n_208),
.Y(n_250)
);

OR2x2_ASAP7_75t_SL g206 ( 
.A(n_152),
.B(n_3),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g267 ( 
.A1(n_206),
.A2(n_225),
.B(n_226),
.Y(n_267)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_114),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_145),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_118),
.Y(n_209)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_211),
.Y(n_270)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_214),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_133),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_213),
.A2(n_220),
.B1(n_221),
.B2(n_224),
.Y(n_258)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_151),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_124),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_215),
.B(n_216),
.Y(n_268)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_158),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_131),
.B(n_4),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_217),
.B(n_218),
.Y(n_255)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_132),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_115),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_114),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_149),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_142),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_222),
.B(n_223),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_177),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_146),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_154),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_4),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_135),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_228),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_119),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_119),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_230),
.Y(n_257)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_137),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_233),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_152),
.B(n_6),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_159),
.Y(n_233)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_137),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_236),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_159),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_116),
.B(n_6),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_136),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_238),
.B(n_241),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_174),
.B(n_6),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g241 ( 
.A(n_117),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_178),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_242),
.A2(n_135),
.B1(n_167),
.B2(n_126),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_161),
.B1(n_138),
.B2(n_134),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_244),
.A2(n_277),
.B1(n_278),
.B2(n_275),
.Y(n_300)
);

OA22x2_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_162),
.B1(n_130),
.B2(n_141),
.Y(n_249)
);

AO21x2_ASAP7_75t_L g302 ( 
.A1(n_249),
.A2(n_187),
.B(n_241),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_139),
.C(n_166),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_251),
.B(n_279),
.C(n_274),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_201),
.A2(n_147),
.B1(n_148),
.B2(n_170),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_252),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_195),
.A2(n_147),
.B1(n_148),
.B2(n_170),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_197),
.A2(n_166),
.B1(n_133),
.B2(n_150),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_234),
.A2(n_150),
.B1(n_160),
.B2(n_172),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_263),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_190),
.A2(n_122),
.B(n_129),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_271),
.A2(n_274),
.B(n_275),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_192),
.A2(n_167),
.B(n_127),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_191),
.A2(n_178),
.B1(n_172),
.B2(n_160),
.Y(n_275)
);

O2A1O1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_276),
.A2(n_271),
.B(n_272),
.C(n_260),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_202),
.A2(n_169),
.B1(n_182),
.B2(n_7),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_235),
.A2(n_8),
.B1(n_212),
.B2(n_203),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_280),
.A2(n_285),
.B(n_263),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_210),
.A2(n_225),
.B(n_207),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_281),
.Y(n_287)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_287),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_220),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_288),
.B(n_294),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_289),
.B(n_254),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_244),
.A2(n_184),
.B1(n_198),
.B2(n_194),
.Y(n_290)
);

AOI22x1_ASAP7_75t_L g346 ( 
.A1(n_290),
.A2(n_302),
.B1(n_314),
.B2(n_320),
.Y(n_346)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_281),
.Y(n_291)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_291),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_184),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_292),
.B(n_300),
.Y(n_347)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_250),
.B(n_227),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_209),
.C(n_214),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_295),
.B(n_304),
.C(n_306),
.Y(n_335)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_296),
.Y(n_329)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_247),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_297),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_255),
.B(n_187),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_311),
.Y(n_325)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_247),
.Y(n_301)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_301),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_251),
.B(n_273),
.C(n_262),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_265),
.A2(n_213),
.B1(n_189),
.B2(n_221),
.Y(n_305)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_305),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_188),
.C(n_200),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_265),
.A2(n_211),
.B1(n_215),
.B2(n_241),
.Y(n_307)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_307),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_257),
.A2(n_215),
.B1(n_276),
.B2(n_267),
.Y(n_308)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_308),
.Y(n_340)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_309),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_248),
.B(n_257),
.C(n_249),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_315),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_256),
.B(n_269),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_264),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_316),
.Y(n_333)
);

AO22x1_ASAP7_75t_L g314 ( 
.A1(n_252),
.A2(n_259),
.B1(n_276),
.B2(n_261),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_248),
.B(n_249),
.C(n_256),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_284),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_249),
.A2(n_277),
.B1(n_243),
.B2(n_272),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_317),
.A2(n_319),
.B(n_280),
.Y(n_334)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_253),
.Y(n_342)
);

MAJx2_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_254),
.C(n_260),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_323),
.C(n_344),
.Y(n_356)
);

A2O1A1Ixp33_ASAP7_75t_L g326 ( 
.A1(n_310),
.A2(n_285),
.B(n_268),
.C(n_246),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_306),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_292),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_328),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_316),
.Y(n_330)
);

BUFx2_ASAP7_75t_SL g360 ( 
.A(n_330),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_291),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_331),
.Y(n_353)
);

NAND3xp33_ASAP7_75t_L g366 ( 
.A(n_334),
.B(n_336),
.C(n_339),
.Y(n_366)
);

AOI322xp5_ASAP7_75t_L g341 ( 
.A1(n_315),
.A2(n_282),
.A3(n_270),
.B1(n_266),
.B2(n_258),
.C1(n_253),
.C2(n_284),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_341),
.Y(n_365)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_342),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_304),
.B(n_266),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_340),
.B(n_317),
.Y(n_349)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_349),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_347),
.A2(n_302),
.B1(n_314),
.B2(n_303),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_350),
.A2(n_352),
.B1(n_355),
.B2(n_358),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_346),
.A2(n_302),
.B(n_312),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_351),
.A2(n_366),
.B(n_369),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_347),
.A2(n_302),
.B1(n_314),
.B2(n_303),
.Y(n_352)
);

AOI22x1_ASAP7_75t_SL g354 ( 
.A1(n_340),
.A2(n_320),
.B1(n_302),
.B2(n_312),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_354),
.A2(n_361),
.B(n_363),
.Y(n_386)
);

OA21x2_ASAP7_75t_L g355 ( 
.A1(n_346),
.A2(n_307),
.B(n_290),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_338),
.A2(n_339),
.B1(n_346),
.B2(n_325),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_357),
.A2(n_324),
.B1(n_327),
.B2(n_329),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_334),
.A2(n_299),
.B1(n_319),
.B2(n_318),
.Y(n_358)
);

XNOR2x1_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_295),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_363),
.C(n_367),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_344),
.B(n_245),
.C(n_299),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_338),
.A2(n_297),
.B1(n_301),
.B2(n_245),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_364),
.A2(n_332),
.B1(n_322),
.B2(n_337),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_343),
.C(n_323),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_333),
.B(n_330),
.Y(n_368)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_368),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_326),
.A2(n_335),
.B(n_329),
.Y(n_369)
);

BUFx24_ASAP7_75t_SL g370 ( 
.A(n_369),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_370),
.B(n_361),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_368),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_375),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_367),
.B(n_321),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_382),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_348),
.Y(n_375)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_362),
.Y(n_378)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_378),
.Y(n_393)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_362),
.Y(n_379)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_379),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_381),
.A2(n_350),
.B1(n_352),
.B2(n_351),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_356),
.B(n_345),
.C(n_324),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_345),
.C(n_327),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_386),
.Y(n_399)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_360),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_384),
.B(n_387),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_353),
.Y(n_391)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_337),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_359),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_390),
.B(n_401),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_391),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_382),
.B(n_348),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_389),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_378),
.B(n_353),
.Y(n_396)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_396),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_372),
.A2(n_349),
.B1(n_365),
.B2(n_366),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_398),
.B(n_400),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_372),
.A2(n_349),
.B1(n_354),
.B2(n_355),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_381),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_403),
.B(n_358),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_404),
.B(n_405),
.Y(n_424)
);

INVx11_ASAP7_75t_L g405 ( 
.A(n_402),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_396),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_413),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_380),
.C(n_383),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_409),
.B(n_380),
.C(n_392),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_393),
.B(n_377),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_376),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_414),
.B(n_394),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_415),
.A2(n_398),
.B1(n_385),
.B2(n_354),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_417),
.B(n_421),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_408),
.A2(n_373),
.B(n_386),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_418),
.A2(n_407),
.B(n_424),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_419),
.B(n_420),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_399),
.C(n_401),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_399),
.C(n_374),
.Y(n_421)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_413),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_422),
.B(n_406),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_423),
.B(n_412),
.Y(n_429)
);

OAI21xp33_ASAP7_75t_L g425 ( 
.A1(n_416),
.A2(n_407),
.B(n_414),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_425),
.B(n_400),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_426),
.A2(n_405),
.B1(n_355),
.B2(n_332),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_417),
.B(n_388),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_411),
.C(n_410),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_429),
.B(n_430),
.Y(n_434)
);

NOR2x1_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_411),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_431),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_428),
.B(n_412),
.C(n_410),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_433),
.B(n_437),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_436),
.B(n_432),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_425),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_440),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_434),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_441),
.A2(n_442),
.B(n_433),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_443),
.B(n_430),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_444),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_445),
.A2(n_446),
.B(n_439),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_447),
.B(n_435),
.C(n_438),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_397),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_449),
.A2(n_355),
.B1(n_322),
.B2(n_364),
.Y(n_450)
);


endmodule