module fake_jpeg_13538_n_491 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_491);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_491;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_479;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_12),
.B(n_13),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_12),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_27),
.B(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_59),
.B(n_72),
.Y(n_128)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_63),
.Y(n_167)
);

BUFx12f_ASAP7_75t_SL g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_64),
.B(n_89),
.Y(n_121)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_65),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_66),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_70),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_71),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_27),
.B(n_16),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_73),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_74),
.B(n_87),
.Y(n_125)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_75),
.Y(n_176)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_76),
.Y(n_153)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_77),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_79),
.Y(n_173)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_81),
.Y(n_194)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_82),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_83),
.Y(n_180)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_84),
.Y(n_175)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_85),
.Y(n_172)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_86),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_15),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_25),
.B(n_11),
.C(n_15),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_91),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_92),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_93),
.B(n_113),
.Y(n_178)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_94),
.B(n_95),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_96),
.B(n_98),
.Y(n_135)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_97),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_0),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_99),
.B(n_101),
.Y(n_147)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_100),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_21),
.B(n_9),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_41),
.B(n_0),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_103),
.Y(n_122)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_104),
.Y(n_166)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_35),
.B(n_0),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_107),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_109),
.Y(n_127)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_45),
.B(n_1),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_33),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_115),
.Y(n_144)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_114),
.B(n_118),
.Y(n_193)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_119),
.Y(n_155)
);

BUFx8_ASAP7_75t_L g118 ( 
.A(n_24),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_18),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_32),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_47),
.B1(n_48),
.B2(n_25),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_129),
.A2(n_145),
.B1(n_151),
.B2(n_170),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_60),
.A2(n_47),
.B1(n_49),
.B2(n_18),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_L g247 ( 
.A1(n_137),
.A2(n_162),
.B1(n_163),
.B2(n_188),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_59),
.B(n_45),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_138),
.B(n_146),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_63),
.A2(n_48),
.B1(n_49),
.B2(n_26),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_143),
.A2(n_149),
.B1(n_161),
.B2(n_142),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_55),
.B1(n_22),
.B2(n_36),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_72),
.B(n_36),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_61),
.A2(n_66),
.B1(n_71),
.B2(n_81),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_104),
.A2(n_29),
.B1(n_22),
.B2(n_44),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_102),
.A2(n_29),
.B(n_43),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_154),
.A2(n_185),
.B(n_131),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_99),
.B(n_44),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_156),
.B(n_159),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_43),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_32),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_160),
.B(n_165),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_L g161 ( 
.A1(n_70),
.A2(n_26),
.B1(n_19),
.B2(n_3),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_107),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_83),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_67),
.B(n_1),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_82),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_168),
.A2(n_156),
.B1(n_193),
.B2(n_146),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_67),
.A2(n_5),
.B1(n_8),
.B2(n_68),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_91),
.B(n_5),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_171),
.B(n_183),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_92),
.B(n_98),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_95),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_184),
.B(n_190),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_68),
.A2(n_78),
.B1(n_96),
.B2(n_108),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_117),
.B(n_78),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_186),
.B(n_171),
.C(n_193),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_118),
.A2(n_60),
.B1(n_63),
.B2(n_66),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_59),
.A2(n_72),
.B(n_101),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_74),
.B(n_106),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_125),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_182),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_195),
.B(n_198),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_193),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_196),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_182),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_171),
.A2(n_122),
.B1(n_168),
.B2(n_121),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_200),
.A2(n_201),
.B1(n_212),
.B2(n_243),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_144),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_202),
.B(n_205),
.Y(n_268)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_203),
.Y(n_302)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_204),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_132),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_206),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_127),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_207),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_164),
.Y(n_208)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_208),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_140),
.B(n_123),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_209),
.B(n_215),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_210),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_147),
.A2(n_128),
.B1(n_190),
.B2(n_138),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_213),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_128),
.A2(n_147),
.B1(n_143),
.B2(n_136),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_214),
.A2(n_242),
.B(n_245),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_154),
.B(n_155),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_158),
.Y(n_216)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_216),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_217),
.A2(n_230),
.B1(n_231),
.B2(n_247),
.Y(n_280)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_141),
.Y(n_218)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_218),
.Y(n_292)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_141),
.Y(n_219)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_186),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_220),
.B(n_237),
.Y(n_279)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_139),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_221),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_164),
.Y(n_223)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_223),
.Y(n_301)
);

OR2x2_ASAP7_75t_SL g224 ( 
.A(n_178),
.B(n_177),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_224),
.B(n_246),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_189),
.A2(n_132),
.B1(n_177),
.B2(n_175),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_225),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_142),
.B(n_189),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_227),
.B(n_229),
.Y(n_307)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_136),
.B(n_172),
.Y(n_228)
);

AND2x4_ASAP7_75t_SL g275 ( 
.A(n_228),
.B(n_238),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_172),
.B(n_133),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_149),
.A2(n_161),
.B1(n_169),
.B2(n_166),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_230),
.A2(n_231),
.B1(n_217),
.B2(n_255),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_166),
.A2(n_169),
.B1(n_167),
.B2(n_134),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_158),
.Y(n_232)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_232),
.Y(n_306)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_176),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_234),
.Y(n_272)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_235),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_175),
.A2(n_148),
.B1(n_173),
.B2(n_153),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_236),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_135),
.Y(n_237)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_173),
.B(n_148),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_153),
.A2(n_180),
.B1(n_130),
.B2(n_126),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_240),
.A2(n_254),
.B1(n_206),
.B2(n_208),
.Y(n_303)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_134),
.Y(n_241)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_178),
.B(n_131),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_185),
.A2(n_180),
.B1(n_167),
.B2(n_139),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_150),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_249),
.Y(n_284)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_187),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_SL g250 ( 
.A(n_150),
.B(n_184),
.C(n_152),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_250),
.B(n_257),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_174),
.A2(n_181),
.B1(n_192),
.B2(n_194),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_251),
.A2(n_247),
.B1(n_238),
.B2(n_221),
.Y(n_287)
);

AND2x2_ASAP7_75t_SL g252 ( 
.A(n_130),
.B(n_152),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_253),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_187),
.A2(n_174),
.B(n_194),
.C(n_192),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_181),
.A2(n_37),
.B1(n_88),
.B2(n_27),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_251),
.Y(n_283)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_182),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_256),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_144),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_258),
.B(n_207),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_262),
.A2(n_265),
.B1(n_280),
.B2(n_293),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_233),
.A2(n_204),
.B1(n_214),
.B2(n_220),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_228),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_276),
.B(n_252),
.Y(n_316)
);

AOI32xp33_ASAP7_75t_L g277 ( 
.A1(n_233),
.A2(n_226),
.A3(n_248),
.B1(n_200),
.B2(n_224),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_277),
.A2(n_291),
.B(n_250),
.Y(n_319)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_283),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_287),
.A2(n_297),
.B1(n_298),
.B2(n_246),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_248),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_299),
.Y(n_311)
);

AOI32xp33_ASAP7_75t_L g291 ( 
.A1(n_212),
.A2(n_222),
.A3(n_258),
.B1(n_202),
.B2(n_211),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_245),
.A2(n_199),
.B1(n_196),
.B2(n_201),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_294),
.B(n_305),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_242),
.A2(n_228),
.B1(n_238),
.B2(n_197),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_242),
.A2(n_197),
.B1(n_253),
.B2(n_235),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_195),
.B(n_198),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_303),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_216),
.B(n_232),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_281),
.A2(n_241),
.B1(n_208),
.B2(n_223),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_308),
.A2(n_321),
.B1(n_328),
.B2(n_332),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_265),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_310),
.B(n_312),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_267),
.B(n_304),
.C(n_277),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_304),
.A2(n_269),
.B(n_288),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_315),
.A2(n_322),
.B(n_327),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_316),
.B(n_324),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_268),
.B(n_234),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_317),
.B(n_326),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_299),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_331),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_SL g347 ( 
.A(n_319),
.B(n_274),
.C(n_292),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_286),
.A2(n_223),
.B1(n_239),
.B2(n_206),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_320),
.A2(n_323),
.B1(n_263),
.B2(n_300),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_281),
.A2(n_203),
.B1(n_213),
.B2(n_218),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_261),
.A2(n_252),
.B(n_256),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_267),
.B(n_219),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_325),
.B(n_330),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_270),
.B(n_210),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_293),
.A2(n_239),
.B1(n_249),
.B2(n_261),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_287),
.A2(n_298),
.B1(n_269),
.B2(n_279),
.Y(n_328)
);

BUFx12f_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_329),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_275),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_270),
.B(n_307),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_269),
.A2(n_262),
.B1(n_276),
.B2(n_297),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_291),
.B(n_266),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_333),
.B(n_342),
.Y(n_363)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_285),
.Y(n_334)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_334),
.Y(n_348)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_285),
.Y(n_335)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_335),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_284),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_338),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_283),
.A2(n_260),
.B1(n_275),
.B2(n_259),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_337),
.A2(n_341),
.B1(n_263),
.B2(n_295),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_275),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_273),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_278),
.Y(n_360)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_306),
.Y(n_340)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_340),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_271),
.A2(n_286),
.B1(n_275),
.B2(n_260),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_282),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_272),
.B(n_282),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_278),
.Y(n_364)
);

OA21x2_ASAP7_75t_L g344 ( 
.A1(n_314),
.A2(n_271),
.B(n_301),
.Y(n_344)
);

AO21x2_ASAP7_75t_L g386 ( 
.A1(n_344),
.A2(n_343),
.B(n_337),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_314),
.A2(n_307),
.B1(n_272),
.B2(n_301),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_345),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_341),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_309),
.B(n_292),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_351),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_342),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_364),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_310),
.B(n_295),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_354),
.Y(n_373)
);

HAxp5_ASAP7_75t_SL g355 ( 
.A(n_315),
.B(n_300),
.CON(n_355),
.SN(n_355)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_355),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_359),
.Y(n_378)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_360),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_365),
.A2(n_323),
.B(n_322),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_313),
.A2(n_289),
.B1(n_296),
.B2(n_302),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_327),
.A2(n_289),
.B1(n_302),
.B2(n_264),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_313),
.A2(n_289),
.B1(n_318),
.B2(n_311),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_325),
.A2(n_328),
.B1(n_332),
.B2(n_321),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_369),
.B(n_371),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_311),
.B(n_339),
.Y(n_371)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_360),
.Y(n_374)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_374),
.Y(n_398)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_364),
.Y(n_376)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_376),
.Y(n_400)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_348),
.Y(n_377)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_377),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_350),
.B(n_312),
.C(n_333),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_379),
.B(n_383),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_380),
.B(n_361),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_363),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_371),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_348),
.Y(n_384)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_384),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_386),
.A2(n_357),
.B1(n_369),
.B2(n_359),
.Y(n_404)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_358),
.Y(n_387)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_387),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_346),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_389),
.Y(n_412)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_356),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_356),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_390),
.B(n_393),
.Y(n_415)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_372),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_352),
.B(n_324),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_394),
.B(n_397),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_361),
.A2(n_319),
.B(n_330),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_396),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_308),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_375),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_408),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_404),
.A2(n_374),
.B1(n_381),
.B2(n_391),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_378),
.A2(n_345),
.B1(n_344),
.B2(n_362),
.Y(n_405)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_405),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_375),
.B(n_346),
.Y(n_406)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_406),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_407),
.A2(n_380),
.B(n_344),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_392),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_392),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_419),
.Y(n_436)
);

FAx1_ASAP7_75t_SL g411 ( 
.A(n_379),
.B(n_363),
.CI(n_368),
.CON(n_411),
.SN(n_411)
);

FAx1_ASAP7_75t_SL g435 ( 
.A(n_411),
.B(n_386),
.CI(n_349),
.CON(n_435),
.SN(n_435)
);

OAI21x1_ASAP7_75t_L g434 ( 
.A1(n_413),
.A2(n_353),
.B(n_373),
.Y(n_434)
);

NAND3xp33_ASAP7_75t_L g416 ( 
.A(n_395),
.B(n_353),
.C(n_370),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_416),
.B(n_418),
.Y(n_422)
);

NOR3xp33_ASAP7_75t_SL g418 ( 
.A(n_391),
.B(n_347),
.C(n_362),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_376),
.A2(n_344),
.B1(n_362),
.B2(n_367),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_396),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_430),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_424),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_403),
.B(n_397),
.C(n_382),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_427),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_399),
.B(n_406),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_412),
.Y(n_428)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_428),
.Y(n_440)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_429),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_408),
.A2(n_386),
.B1(n_385),
.B2(n_394),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_413),
.B(n_349),
.C(n_373),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_431),
.B(n_432),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_413),
.B(n_411),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_398),
.Y(n_433)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_433),
.Y(n_444)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_434),
.Y(n_451)
);

FAx1_ASAP7_75t_SL g442 ( 
.A(n_435),
.B(n_411),
.CI(n_386),
.CON(n_442),
.SN(n_442)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_417),
.B(n_385),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_437),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_420),
.A2(n_398),
.B1(n_417),
.B2(n_400),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_438),
.B(n_442),
.Y(n_459)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_421),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_436),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_429),
.A2(n_407),
.B(n_405),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_448),
.A2(n_424),
.B(n_407),
.Y(n_454)
);

OAI31xp33_ASAP7_75t_SL g450 ( 
.A1(n_435),
.A2(n_402),
.A3(n_409),
.B(n_386),
.Y(n_450)
);

OAI321xp33_ASAP7_75t_L g456 ( 
.A1(n_450),
.A2(n_421),
.A3(n_436),
.B1(n_425),
.B2(n_420),
.C(n_400),
.Y(n_456)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_440),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_452),
.B(n_453),
.Y(n_464)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_444),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_454),
.A2(n_441),
.B1(n_439),
.B2(n_450),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_443),
.B(n_426),
.C(n_437),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_455),
.B(n_457),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_456),
.A2(n_357),
.B1(n_410),
.B2(n_401),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_443),
.B(n_432),
.C(n_423),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_451),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_461),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_449),
.C(n_445),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_460),
.B(n_449),
.C(n_447),
.Y(n_463)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_439),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_462),
.A2(n_414),
.B1(n_387),
.B2(n_358),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_463),
.B(n_470),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_465),
.B(n_468),
.Y(n_472)
);

NOR2x1_ASAP7_75t_L g466 ( 
.A(n_460),
.B(n_422),
.Y(n_466)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_466),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_459),
.A2(n_430),
.B1(n_419),
.B2(n_441),
.Y(n_467)
);

AOI322xp5_ASAP7_75t_L g476 ( 
.A1(n_467),
.A2(n_462),
.A3(n_442),
.B1(n_435),
.B2(n_418),
.C1(n_370),
.C2(n_431),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_466),
.A2(n_457),
.B(n_455),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_476),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_463),
.A2(n_454),
.B(n_448),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_474),
.A2(n_470),
.B(n_442),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_427),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_478),
.B(n_472),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_471),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_480),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_477),
.B(n_468),
.C(n_467),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_481),
.B(n_482),
.C(n_483),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_479),
.B(n_472),
.C(n_465),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_486),
.A2(n_464),
.B(n_414),
.Y(n_487)
);

OAI211xp5_ASAP7_75t_L g489 ( 
.A1(n_487),
.A2(n_488),
.B(n_415),
.C(n_401),
.Y(n_489)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_485),
.Y(n_488)
);

MAJx2_ASAP7_75t_L g490 ( 
.A(n_489),
.B(n_484),
.C(n_410),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_490),
.B(n_384),
.Y(n_491)
);


endmodule