module fake_netlist_1_325_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_10), .Y(n_12) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
BUFx6f_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
INVxp67_ASAP7_75t_L g16 ( .A(n_5), .Y(n_16) );
INVx3_ASAP7_75t_L g17 ( .A(n_8), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_13), .B(n_1), .Y(n_18) );
CKINVDCx16_ASAP7_75t_R g19 ( .A(n_11), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_11), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_17), .B(n_1), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_15), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_21), .A2(n_15), .B1(n_16), .B2(n_14), .Y(n_24) );
AND2x4_ASAP7_75t_L g25 ( .A(n_21), .B(n_17), .Y(n_25) );
NAND3xp33_ASAP7_75t_L g26 ( .A(n_18), .B(n_14), .C(n_12), .Y(n_26) );
NAND3xp33_ASAP7_75t_L g27 ( .A(n_24), .B(n_19), .C(n_21), .Y(n_27) );
INVx2_ASAP7_75t_SL g28 ( .A(n_25), .Y(n_28) );
AOI221xp5_ASAP7_75t_L g29 ( .A1(n_23), .A2(n_20), .B1(n_14), .B2(n_17), .C(n_2), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_20), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_27), .B(n_25), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
OAI32xp33_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_17), .A3(n_26), .B1(n_29), .B2(n_2), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
OAI22xp5_ASAP7_75t_L g36 ( .A1(n_32), .A2(n_14), .B1(n_4), .B2(n_3), .Y(n_36) );
INVx2_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
NAND4xp75_ASAP7_75t_L g38 ( .A(n_36), .B(n_3), .C(n_14), .D(n_7), .Y(n_38) );
AOI21xp33_ASAP7_75t_L g39 ( .A1(n_37), .A2(n_34), .B(n_6), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_38), .Y(n_40) );
NAND3xp33_ASAP7_75t_L g41 ( .A(n_40), .B(n_9), .C(n_39), .Y(n_41) );
endmodule