module fake_jpeg_18485_n_45 (n_3, n_2, n_1, n_0, n_4, n_5, n_45);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_45;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx5_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_16),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_14),
.B(n_15),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_7),
.B(n_0),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_18),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_7),
.B(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_11),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_10),
.C(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_23),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_15),
.A2(n_4),
.B1(n_5),
.B2(n_2),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_25),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_16),
.B1(n_13),
.B2(n_4),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_12),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_22),
.C(n_25),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_26),
.C(n_30),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_38),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

A2O1A1O1Ixp25_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_1),
.B(n_2),
.C(n_37),
.D(n_36),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_43),
.B(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_1),
.Y(n_45)
);


endmodule