module real_jpeg_21814_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_333, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_332, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_333;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_332;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_0),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_0),
.A2(n_27),
.B1(n_31),
.B2(n_101),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_0),
.A2(n_50),
.B1(n_51),
.B2(n_101),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_101),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_1),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_1),
.B(n_22),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g156 ( 
.A1(n_1),
.A2(n_16),
.B(n_50),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_106),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_1),
.A2(n_84),
.B1(n_87),
.B2(n_165),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_1),
.B(n_61),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g194 ( 
.A1(n_1),
.A2(n_25),
.B(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_2),
.A2(n_27),
.B1(n_31),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_35),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_2),
.A2(n_35),
.B1(n_50),
.B2(n_51),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_2),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_3),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_103),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_103),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_3),
.A2(n_27),
.B1(n_31),
.B2(n_103),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_4),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_91),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_91),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_4),
.A2(n_27),
.B1(n_31),
.B2(n_91),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_5),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_97),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_97),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_5),
.A2(n_27),
.B1(n_31),
.B2(n_97),
.Y(n_257)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_7),
.A2(n_27),
.B1(n_31),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_7),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_108),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_108),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_7),
.A2(n_50),
.B1(n_51),
.B2(n_108),
.Y(n_165)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_8),
.A2(n_148),
.B1(n_149),
.B2(n_151),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_9),
.A2(n_27),
.B1(n_31),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_9),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_9),
.A2(n_50),
.B1(n_51),
.B2(n_69),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_69),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_69),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_10),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_10),
.A2(n_30),
.B1(n_46),
.B2(n_47),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_10),
.A2(n_30),
.B1(n_50),
.B2(n_51),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_12),
.A2(n_27),
.B1(n_31),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_66),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_66),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_66),
.Y(n_261)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_59)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_14),
.A2(n_25),
.A3(n_47),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_15),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_16),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_16),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_16),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

BUFx3_ASAP7_75t_SL g47 ( 
.A(n_17),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_38),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_26),
.B(n_29),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_23),
.B(n_27),
.C(n_28),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_26),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_22),
.A2(n_26),
.B1(n_34),
.B2(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_22),
.A2(n_26),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_22),
.A2(n_26),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_27),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_23),
.B(n_25),
.Y(n_120)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_24),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_24),
.B(n_57),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_24),
.A2(n_28),
.B1(n_105),
.B2(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_24),
.B(n_106),
.Y(n_191)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

HAxp5_ASAP7_75t_SL g105 ( 
.A(n_27),
.B(n_106),
.CON(n_105),
.SN(n_105)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_33),
.B(n_40),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_74),
.B(n_330),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_70),
.C(n_72),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_41),
.A2(n_42),
.B1(n_326),
.B2(n_328),
.Y(n_325)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_53),
.C(n_62),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_43),
.A2(n_297),
.B1(n_298),
.B2(n_300),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_43),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_43),
.A2(n_53),
.B1(n_300),
.B2(n_313),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_49),
.B(n_52),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_44),
.A2(n_49),
.B1(n_90),
.B2(n_92),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_44),
.A2(n_49),
.B1(n_90),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_44),
.A2(n_49),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_44),
.A2(n_49),
.B1(n_160),
.B2(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_44),
.A2(n_49),
.B1(n_180),
.B2(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_44),
.A2(n_49),
.B1(n_96),
.B2(n_198),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_44),
.A2(n_49),
.B1(n_92),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_44),
.A2(n_49),
.B1(n_234),
.B2(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_44),
.A2(n_49),
.B1(n_52),
.B2(n_267),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_46),
.B(n_57),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_47),
.A2(n_48),
.B(n_106),
.C(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_49),
.B(n_106),
.Y(n_163)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_50),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_51),
.B(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_53),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_54),
.A2(n_55),
.B1(n_61),
.B2(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_60),
.B(n_61),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_55),
.A2(n_61),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_55),
.A2(n_61),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_56),
.A2(n_59),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_56),
.A2(n_59),
.B1(n_102),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_56),
.A2(n_59),
.B1(n_132),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_56),
.A2(n_59),
.B1(n_116),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_56),
.A2(n_59),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_62),
.A2(n_63),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_64),
.A2(n_67),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_64),
.A2(n_67),
.B1(n_114),
.B2(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_64),
.A2(n_67),
.B1(n_241),
.B2(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_327),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_72),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_323),
.B(n_329),
.Y(n_74)
);

OAI321xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_292),
.A3(n_315),
.B1(n_321),
.B2(n_322),
.C(n_332),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_271),
.B(n_291),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_247),
.B(n_270),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_140),
.B(n_223),
.C(n_246),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_123),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_80),
.B(n_123),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_109),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_93),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_82),
.B(n_93),
.C(n_109),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_89),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_83),
.B(n_89),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_84),
.A2(n_122),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_84),
.A2(n_87),
.B1(n_150),
.B2(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_84),
.A2(n_87),
.B1(n_152),
.B2(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_84),
.A2(n_85),
.B1(n_137),
.B2(n_182),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_84),
.A2(n_87),
.B1(n_88),
.B2(n_232),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_84),
.A2(n_138),
.B(n_232),
.Y(n_265)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.C(n_104),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_106),
.B(n_138),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_107),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_118),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_117),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_111),
.B(n_117),
.C(n_118),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_115),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_121),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.C(n_128),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_124),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.C(n_135),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_130),
.B(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_134),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_222),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_217),
.B(n_221),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_203),
.B(n_216),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_184),
.B(n_202),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_172),
.B(n_183),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_161),
.B(n_171),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_153),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_153),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_157),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_166),
.B(n_170),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_164),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_174),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_181),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_179),
.C(n_181),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_186),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_192),
.B1(n_200),
.B2(n_201),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_187),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_189),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_191),
.Y(n_195)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_196),
.B1(n_197),
.B2(n_199),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_193),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_199),
.C(n_200),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_204),
.B(n_205),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_213),
.C(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_212),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_213),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_218),
.B(n_219),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_224),
.B(n_225),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_245),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_226),
.Y(n_245)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_235),
.B2(n_236),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_236),
.C(n_245),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_239),
.C(n_244),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_244),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_242),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_243),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_248),
.B(n_249),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_269),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_262),
.B2(n_263),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_263),
.C(n_269),
.Y(n_272)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_255),
.C(n_259),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_257),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_261),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_268),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_264),
.A2(n_265),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_266),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_265),
.A2(n_283),
.B1(n_286),
.B2(n_333),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_266),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_272),
.B(n_273),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_289),
.B2(n_290),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_282),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_276),
.B(n_282),
.C(n_290),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B(n_281),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_280),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_294),
.C(n_305),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_281),
.A2(n_294),
.B1(n_295),
.B2(n_320),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_281),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_288),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_289),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_307),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_307),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.Y(n_295)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_296),
.Y(n_303)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_300),
.C(n_301),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_301),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_301),
.A2(n_304),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_309),
.C(n_314),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_305),
.A2(n_306),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_314),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_316),
.B(n_317),
.Y(n_321)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_326),
.Y(n_328)
);


endmodule