module real_aes_7708_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_635;
wire n_357;
wire n_503;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_577;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_1064;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_1034;
wire n_376;
wire n_549;
wire n_694;
wire n_491;
wire n_923;
wire n_571;
wire n_894;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_884;
wire n_537;
wire n_551;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_1021;
wire n_399;
wire n_700;
wire n_948;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_774;
wire n_992;
wire n_813;
wire n_981;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_369;
wire n_726;
wire n_517;
wire n_931;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_973;
wire n_455;
wire n_725;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_1006;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_769;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_869;
wire n_613;
wire n_642;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_756;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_997;
wire n_569;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1003;
wire n_1000;
wire n_1028;
wire n_366;
wire n_727;
wire n_1014;
wire n_397;
wire n_358;
wire n_385;
wire n_1056;
wire n_663;
wire n_749;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_354;
wire n_972;
wire n_435;
wire n_710;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_831;
wire n_487;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_922;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_968;
wire n_646;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g664 ( .A1(n_0), .A2(n_158), .B1(n_665), .B2(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_1), .B(n_438), .Y(n_551) );
XOR2x2_ASAP7_75t_L g512 ( .A(n_2), .B(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g984 ( .A(n_3), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_4), .A2(n_272), .B1(n_630), .B2(n_631), .Y(n_629) );
OA22x2_ASAP7_75t_L g608 ( .A1(n_5), .A2(n_609), .B1(n_610), .B2(n_639), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_5), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_6), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_7), .A2(n_77), .B1(n_634), .B2(n_635), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g856 ( .A1(n_8), .A2(n_261), .B1(n_580), .B2(n_662), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_9), .A2(n_319), .B1(n_966), .B2(n_973), .Y(n_1027) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_10), .Y(n_488) );
AO22x2_ASAP7_75t_L g376 ( .A1(n_11), .A2(n_196), .B1(n_377), .B2(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g1017 ( .A(n_11), .Y(n_1017) );
AOI22xp33_ASAP7_75t_SL g787 ( .A1(n_12), .A2(n_182), .B1(n_518), .B2(n_788), .Y(n_787) );
AOI22xp5_ASAP7_75t_SL g890 ( .A1(n_13), .A2(n_346), .B1(n_502), .B2(n_666), .Y(n_890) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_14), .A2(n_274), .B1(n_463), .B2(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_15), .A2(n_57), .B1(n_621), .B2(n_833), .Y(n_832) );
AOI22xp5_ASAP7_75t_SL g886 ( .A1(n_16), .A2(n_222), .B1(n_494), .B2(n_697), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_17), .A2(n_101), .B1(n_492), .B2(n_783), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_18), .A2(n_23), .B1(n_662), .B2(n_1032), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_19), .A2(n_349), .B1(n_504), .B2(n_709), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_20), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_21), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_22), .A2(n_338), .B1(n_425), .B2(n_506), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_24), .A2(n_237), .B1(n_557), .B2(n_559), .Y(n_863) );
INVx1_ASAP7_75t_L g533 ( .A(n_25), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_26), .A2(n_333), .B1(n_425), .B2(n_637), .Y(n_636) );
AOI22xp33_ASAP7_75t_SL g883 ( .A1(n_27), .A2(n_160), .B1(n_527), .B2(n_884), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_28), .A2(n_307), .B1(n_566), .B2(n_567), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_29), .A2(n_89), .B1(n_464), .B2(n_535), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_30), .A2(n_366), .B1(n_466), .B2(n_467), .Y(n_365) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_30), .Y(n_466) );
AOI22xp33_ASAP7_75t_SL g844 ( .A1(n_31), .A2(n_49), .B1(n_722), .B2(n_845), .Y(n_844) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_32), .Y(n_623) );
AO22x2_ASAP7_75t_L g381 ( .A1(n_33), .A2(n_106), .B1(n_377), .B2(n_382), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g755 ( .A1(n_34), .A2(n_232), .B1(n_590), .B2(n_756), .Y(n_755) );
AOI22xp33_ASAP7_75t_SL g686 ( .A1(n_35), .A2(n_97), .B1(n_621), .B2(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_36), .A2(n_248), .B1(n_516), .B2(n_783), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g962 ( .A(n_37), .Y(n_962) );
AOI22xp5_ASAP7_75t_L g1050 ( .A1(n_38), .A2(n_54), .B1(n_421), .B2(n_785), .Y(n_1050) );
AOI22xp33_ASAP7_75t_SL g667 ( .A1(n_39), .A2(n_296), .B1(n_595), .B2(n_668), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_40), .A2(n_201), .B1(n_816), .B2(n_931), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_41), .B(n_655), .Y(n_836) );
AOI22xp33_ASAP7_75t_SL g851 ( .A1(n_42), .A2(n_244), .B1(n_421), .B2(n_759), .Y(n_851) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_43), .A2(n_134), .B1(n_267), .B2(n_454), .C1(n_458), .C2(n_462), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_44), .A2(n_240), .B1(n_484), .B2(n_579), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g912 ( .A(n_45), .Y(n_912) );
AOI22xp33_ASAP7_75t_SL g650 ( .A1(n_46), .A2(n_176), .B1(n_579), .B2(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_47), .A2(n_130), .B1(n_494), .B2(n_499), .Y(n_846) );
AOI22xp5_ASAP7_75t_SL g1049 ( .A1(n_48), .A2(n_193), .B1(n_502), .B2(n_722), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_50), .B(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_51), .Y(n_739) );
AOI22xp33_ASAP7_75t_SL g991 ( .A1(n_52), .A2(n_301), .B1(n_635), .B2(n_672), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_53), .A2(n_190), .B1(n_504), .B2(n_637), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_55), .A2(n_170), .B1(n_902), .B2(n_903), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g954 ( .A(n_56), .Y(n_954) );
CKINVDCx20_ASAP7_75t_R g916 ( .A(n_58), .Y(n_916) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_59), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_60), .A2(n_334), .B1(n_559), .B2(n_560), .Y(n_558) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_61), .A2(n_269), .B1(n_556), .B2(n_557), .Y(n_555) );
AOI22xp5_ASAP7_75t_SL g977 ( .A1(n_62), .A2(n_978), .B1(n_997), .B2(n_998), .Y(n_977) );
CKINVDCx16_ASAP7_75t_R g998 ( .A(n_62), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_63), .A2(n_183), .B1(n_410), .B2(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g892 ( .A(n_64), .Y(n_892) );
AOI222xp33_ASAP7_75t_L g940 ( .A1(n_65), .A2(n_181), .B1(n_215), .B2(n_648), .C1(n_807), .C2(n_808), .Y(n_940) );
CKINVDCx20_ASAP7_75t_R g956 ( .A(n_66), .Y(n_956) );
CKINVDCx20_ASAP7_75t_R g988 ( .A(n_67), .Y(n_988) );
AOI22xp33_ASAP7_75t_SL g674 ( .A1(n_68), .A2(n_242), .B1(n_506), .B2(n_675), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_69), .A2(n_251), .B1(n_410), .B2(n_845), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_70), .A2(n_133), .B1(n_419), .B2(n_556), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_71), .A2(n_227), .B1(n_459), .B2(n_528), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_72), .A2(n_209), .B1(n_492), .B2(n_816), .Y(n_815) );
AOI22xp5_ASAP7_75t_SL g887 ( .A1(n_73), .A2(n_225), .B1(n_499), .B2(n_888), .Y(n_887) );
AOI22xp33_ASAP7_75t_SL g837 ( .A1(n_74), .A2(n_202), .B1(n_535), .B2(n_838), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_75), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_76), .A2(n_223), .B1(n_506), .B2(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g996 ( .A1(n_78), .A2(n_122), .B1(n_499), .B2(n_722), .Y(n_996) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_79), .A2(n_250), .B1(n_556), .B2(n_600), .Y(n_599) );
AOI22xp5_ASAP7_75t_SL g1052 ( .A1(n_80), .A2(n_91), .B1(n_506), .B2(n_931), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_81), .A2(n_276), .B1(n_504), .B2(n_785), .Y(n_784) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_82), .A2(n_192), .B1(n_595), .B2(n_597), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_83), .A2(n_111), .B1(n_494), .B2(n_845), .Y(n_938) );
CKINVDCx20_ASAP7_75t_R g855 ( .A(n_84), .Y(n_855) );
AO22x2_ASAP7_75t_L g384 ( .A1(n_85), .A2(n_231), .B1(n_377), .B2(n_378), .Y(n_384) );
INVx1_ASAP7_75t_L g1014 ( .A(n_85), .Y(n_1014) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_86), .A2(n_351), .B(n_359), .C(n_1019), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_87), .A2(n_93), .B1(n_590), .B2(n_592), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g695 ( .A1(n_88), .A2(n_288), .B1(n_371), .B2(n_600), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_90), .Y(n_408) );
AOI22xp33_ASAP7_75t_SL g1053 ( .A1(n_92), .A2(n_180), .B1(n_566), .B2(n_567), .Y(n_1053) );
INVx1_ASAP7_75t_L g1043 ( .A(n_94), .Y(n_1043) );
AOI22xp5_ASAP7_75t_SL g891 ( .A1(n_95), .A2(n_187), .B1(n_410), .B2(n_675), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_96), .A2(n_271), .B1(n_722), .B2(n_790), .Y(n_939) );
AOI211xp5_ASAP7_75t_L g696 ( .A1(n_98), .A2(n_697), .B(n_698), .C(n_701), .Y(n_696) );
AOI22xp33_ASAP7_75t_SL g689 ( .A1(n_99), .A2(n_257), .B1(n_547), .B2(n_690), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g1020 ( .A1(n_100), .A2(n_1021), .B1(n_1022), .B2(n_1034), .Y(n_1020) );
CKINVDCx20_ASAP7_75t_R g1034 ( .A(n_100), .Y(n_1034) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_102), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g896 ( .A1(n_103), .A2(n_897), .B1(n_922), .B2(n_923), .Y(n_896) );
INVx1_ASAP7_75t_L g922 ( .A(n_103), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_104), .A2(n_110), .B1(n_807), .B2(n_808), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_105), .A2(n_162), .B1(n_458), .B2(n_528), .Y(n_717) );
INVx1_ASAP7_75t_L g1018 ( .A(n_106), .Y(n_1018) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_107), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_108), .B(n_918), .Y(n_917) );
CKINVDCx20_ASAP7_75t_R g951 ( .A(n_109), .Y(n_951) );
AOI22xp33_ASAP7_75t_SL g936 ( .A1(n_112), .A2(n_303), .B1(n_528), .B2(n_662), .Y(n_936) );
AOI22xp33_ASAP7_75t_SL g670 ( .A1(n_113), .A2(n_179), .B1(n_671), .B2(n_672), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_114), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_115), .B(n_433), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g1056 ( .A(n_116), .Y(n_1056) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_117), .A2(n_185), .B1(n_658), .B2(n_660), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_118), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_119), .A2(n_128), .B1(n_463), .B2(n_484), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g1060 ( .A1(n_120), .A2(n_229), .B1(n_580), .B2(n_662), .Y(n_1060) );
AOI22xp33_ASAP7_75t_SL g841 ( .A1(n_121), .A2(n_167), .B1(n_516), .B2(n_756), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_123), .A2(n_304), .B1(n_631), .B2(n_722), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_124), .A2(n_217), .B1(n_528), .B2(n_535), .Y(n_552) );
AOI22xp33_ASAP7_75t_SL g878 ( .A1(n_125), .A2(n_314), .B1(n_463), .B2(n_651), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_126), .A2(n_171), .B1(n_433), .B2(n_436), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_127), .A2(n_331), .B1(n_762), .B2(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g568 ( .A(n_129), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_131), .B(n_438), .Y(n_859) );
AND2x6_ASAP7_75t_L g353 ( .A(n_132), .B(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g1011 ( .A(n_132), .Y(n_1011) );
AOI22xp33_ASAP7_75t_SL g501 ( .A1(n_135), .A2(n_337), .B1(n_502), .B2(n_504), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_136), .A2(n_169), .B1(n_564), .B2(n_672), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g1062 ( .A(n_137), .Y(n_1062) );
CKINVDCx20_ASAP7_75t_R g981 ( .A(n_138), .Y(n_981) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_139), .B(n_432), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_140), .A2(n_320), .B1(n_506), .B2(n_507), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_141), .A2(n_172), .B1(n_419), .B2(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_142), .B(n_655), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_143), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g934 ( .A(n_144), .Y(n_934) );
AOI22xp33_ASAP7_75t_SL g719 ( .A1(n_145), .A2(n_163), .B1(n_564), .B2(n_720), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_146), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_147), .B(n_550), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_148), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g417 ( .A(n_149), .Y(n_417) );
AOI222xp33_ASAP7_75t_L g1033 ( .A1(n_150), .A2(n_184), .B1(n_308), .B2(n_462), .C1(n_486), .C2(n_778), .Y(n_1033) );
AOI22xp33_ASAP7_75t_SL g691 ( .A1(n_151), .A2(n_210), .B1(n_433), .B2(n_655), .Y(n_691) );
AO22x2_ASAP7_75t_L g386 ( .A1(n_152), .A2(n_224), .B1(n_377), .B2(n_382), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g1015 ( .A(n_152), .B(n_1016), .Y(n_1015) );
CKINVDCx20_ASAP7_75t_R g946 ( .A(n_153), .Y(n_946) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_154), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g862 ( .A1(n_155), .A2(n_263), .B1(n_412), .B2(n_673), .Y(n_862) );
AOI22xp33_ASAP7_75t_SL g965 ( .A1(n_156), .A2(n_165), .B1(n_603), .B2(n_966), .Y(n_965) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_157), .A2(n_239), .B1(n_507), .B2(n_694), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_159), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_161), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_164), .A2(n_233), .B1(n_559), .B2(n_722), .Y(n_721) );
AOI22xp33_ASAP7_75t_SL g967 ( .A1(n_166), .A2(n_295), .B1(n_668), .B2(n_968), .Y(n_967) );
CKINVDCx20_ASAP7_75t_R g921 ( .A(n_168), .Y(n_921) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_173), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_174), .Y(n_616) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_175), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_177), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_178), .A2(n_275), .B1(n_372), .B2(n_790), .Y(n_789) );
XNOR2xp5_ASAP7_75t_L g681 ( .A(n_186), .B(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_SL g491 ( .A1(n_188), .A2(n_216), .B1(n_492), .B2(n_494), .Y(n_491) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_189), .A2(n_208), .B1(n_496), .B2(n_499), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_191), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_194), .A2(n_214), .B1(n_372), .B2(n_504), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_195), .A2(n_309), .B1(n_907), .B2(n_908), .Y(n_906) );
NAND2xp5_ASAP7_75t_SL g882 ( .A(n_197), .B(n_432), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_198), .A2(n_325), .B1(n_463), .B2(n_618), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_199), .A2(n_236), .B1(n_566), .B2(n_567), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_200), .A2(n_243), .B1(n_618), .B2(n_619), .Y(n_617) );
AOI22xp33_ASAP7_75t_SL g757 ( .A1(n_203), .A2(n_278), .B1(n_631), .B2(n_758), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_204), .B(n_668), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_205), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_206), .A2(n_330), .B1(n_419), .B2(n_993), .Y(n_992) );
OA22x2_ASAP7_75t_L g469 ( .A1(n_207), .A2(n_470), .B1(n_471), .B2(n_472), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_207), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_211), .A2(n_226), .B1(n_556), .B2(n_785), .Y(n_932) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_212), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_213), .A2(n_298), .B1(n_592), .B2(n_931), .Y(n_1024) );
CKINVDCx20_ASAP7_75t_R g961 ( .A(n_218), .Y(n_961) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_219), .Y(n_877) );
AOI22xp33_ASAP7_75t_SL g707 ( .A1(n_220), .A2(n_268), .B1(n_556), .B2(n_567), .Y(n_707) );
AND2x2_ASAP7_75t_L g357 ( .A(n_221), .B(n_358), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_228), .Y(n_479) );
XNOR2x1_ASAP7_75t_L g827 ( .A(n_230), .B(n_828), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_234), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_235), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_238), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_241), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_245), .Y(n_825) );
AOI22xp33_ASAP7_75t_SL g971 ( .A1(n_246), .A2(n_266), .B1(n_560), .B2(n_635), .Y(n_971) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_247), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_249), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_252), .Y(n_749) );
OA22x2_ASAP7_75t_L g794 ( .A1(n_253), .A2(n_795), .B1(n_796), .B2(n_797), .Y(n_794) );
CKINVDCx16_ASAP7_75t_R g795 ( .A(n_253), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_254), .B(n_432), .Y(n_935) );
CKINVDCx20_ASAP7_75t_R g1057 ( .A(n_255), .Y(n_1057) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_256), .A2(n_322), .B1(n_499), .B2(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g377 ( .A(n_258), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_258), .Y(n_379) );
CKINVDCx20_ASAP7_75t_R g958 ( .A(n_259), .Y(n_958) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_260), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_262), .A2(n_306), .B1(n_758), .B2(n_790), .Y(n_817) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_264), .A2(n_347), .B1(n_432), .B2(n_436), .C(n_439), .Y(n_431) );
AOI22xp33_ASAP7_75t_SL g563 ( .A1(n_265), .A2(n_299), .B1(n_496), .B2(n_564), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_270), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g1064 ( .A(n_273), .Y(n_1064) );
CKINVDCx20_ASAP7_75t_R g911 ( .A(n_277), .Y(n_911) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_279), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_280), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_281), .A2(n_643), .B1(n_644), .B2(n_676), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_281), .Y(n_643) );
XNOR2x1_ASAP7_75t_L g765 ( .A(n_282), .B(n_766), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g987 ( .A(n_283), .Y(n_987) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_284), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_285), .A2(n_328), .B1(n_527), .B2(n_530), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_286), .Y(n_920) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_287), .Y(n_723) );
INVx1_ASAP7_75t_L g358 ( .A(n_289), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_290), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_291), .Y(n_743) );
INVx1_ASAP7_75t_L g354 ( .A(n_292), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_293), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_294), .Y(n_573) );
AOI22xp33_ASAP7_75t_SL g995 ( .A1(n_297), .A2(n_336), .B1(n_425), .B2(n_566), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_300), .A2(n_343), .B1(n_464), .B2(n_547), .Y(n_774) );
XOR2x2_ASAP7_75t_L g732 ( .A(n_302), .B(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_305), .B(n_524), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_310), .A2(n_342), .B1(n_580), .B2(n_662), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g1059 ( .A(n_311), .Y(n_1059) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_312), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_313), .Y(n_423) );
CKINVDCx20_ASAP7_75t_R g831 ( .A(n_315), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_316), .B(n_550), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_317), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_318), .A2(n_348), .B1(n_524), .B2(n_525), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g982 ( .A(n_321), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_323), .A2(n_332), .B1(n_675), .B2(n_783), .Y(n_1028) );
XNOR2x1_ASAP7_75t_L g569 ( .A(n_324), .B(n_570), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_326), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_327), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_329), .B(n_438), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_335), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_339), .B(n_484), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_340), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g950 ( .A(n_341), .Y(n_950) );
CKINVDCx20_ASAP7_75t_R g941 ( .A(n_344), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_345), .B(n_881), .Y(n_880) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
HB1xp67_ASAP7_75t_L g1010 ( .A(n_354), .Y(n_1010) );
OAI21xp5_ASAP7_75t_L g1041 ( .A1(n_355), .A2(n_1009), .B(n_1042), .Y(n_1041) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_870), .B1(n_1004), .B2(n_1005), .C(n_1006), .Y(n_359) );
INVx1_ASAP7_75t_L g1004 ( .A(n_360), .Y(n_1004) );
XNOR2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_605), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_363), .B1(n_508), .B2(n_604), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_468), .B2(n_469), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g467 ( .A(n_366), .Y(n_467) );
AND4x1_ASAP7_75t_L g366 ( .A(n_367), .B(n_406), .C(n_431), .D(n_453), .Y(n_366) );
NOR2xp33_ASAP7_75t_SL g367 ( .A(n_368), .B(n_393), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B1(n_387), .B2(n_388), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx3_ASAP7_75t_L g494 ( .A(n_373), .Y(n_494) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_373), .Y(n_566) );
INVx2_ASAP7_75t_L g638 ( .A(n_373), .Y(n_638) );
BUFx3_ASAP7_75t_L g709 ( .A(n_373), .Y(n_709) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_383), .Y(n_373) );
AND2x4_ASAP7_75t_L g390 ( .A(n_374), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g426 ( .A(n_374), .B(n_415), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_374), .B(n_398), .Y(n_430) );
AND2x2_ASAP7_75t_L g503 ( .A(n_374), .B(n_398), .Y(n_503) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_380), .Y(n_374) );
AND2x2_ASAP7_75t_L g397 ( .A(n_375), .B(n_381), .Y(n_397) );
OR2x2_ASAP7_75t_L g414 ( .A(n_375), .B(n_381), .Y(n_414) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g444 ( .A(n_376), .B(n_386), .Y(n_444) );
AND2x2_ASAP7_75t_L g450 ( .A(n_376), .B(n_381), .Y(n_450) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g382 ( .A(n_379), .Y(n_382) );
INVx1_ASAP7_75t_L g445 ( .A(n_380), .Y(n_445) );
AND2x2_ASAP7_75t_L g460 ( .A(n_380), .B(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g405 ( .A(n_381), .Y(n_405) );
AND2x4_ASAP7_75t_L g435 ( .A(n_383), .B(n_413), .Y(n_435) );
AND2x6_ASAP7_75t_L g438 ( .A(n_383), .B(n_397), .Y(n_438) );
INVx1_ASAP7_75t_L g478 ( .A(n_383), .Y(n_478) );
NAND2x1p5_ASAP7_75t_L g481 ( .A(n_383), .B(n_397), .Y(n_481) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_384), .B(n_386), .Y(n_392) );
INVx1_ASAP7_75t_L g399 ( .A(n_384), .Y(n_399) );
INVx1_ASAP7_75t_L g416 ( .A(n_384), .Y(n_416) );
INVx1_ASAP7_75t_L g461 ( .A(n_384), .Y(n_461) );
AND2x2_ASAP7_75t_L g415 ( .A(n_385), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g398 ( .A(n_386), .B(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx3_ASAP7_75t_L g504 ( .A(n_390), .Y(n_504) );
BUFx3_ASAP7_75t_L g557 ( .A(n_390), .Y(n_557) );
INVx1_ASAP7_75t_L g601 ( .A(n_390), .Y(n_601) );
BUFx2_ASAP7_75t_SL g635 ( .A(n_390), .Y(n_635) );
BUFx2_ASAP7_75t_L g666 ( .A(n_390), .Y(n_666) );
BUFx2_ASAP7_75t_SL g756 ( .A(n_390), .Y(n_756) );
BUFx3_ASAP7_75t_L g931 ( .A(n_390), .Y(n_931) );
AND2x2_ASAP7_75t_L g567 ( .A(n_391), .B(n_445), .Y(n_567) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OR2x6_ASAP7_75t_L g404 ( .A(n_392), .B(n_405), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B1(n_400), .B2(n_401), .Y(n_393) );
OAI21xp33_ASAP7_75t_L g698 ( .A1(n_395), .A2(n_699), .B(n_700), .Y(n_698) );
BUFx2_ASAP7_75t_R g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_397), .B(n_398), .Y(n_396) );
AND2x4_ASAP7_75t_L g421 ( .A(n_397), .B(n_415), .Y(n_421) );
AND2x2_ASAP7_75t_L g498 ( .A(n_397), .B(n_398), .Y(n_498) );
INVx1_ASAP7_75t_L g452 ( .A(n_399), .Y(n_452) );
INVxp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx2_ASAP7_75t_L g499 ( .A(n_403), .Y(n_499) );
BUFx2_ASAP7_75t_L g790 ( .A(n_403), .Y(n_790) );
BUFx4f_ASAP7_75t_SL g908 ( .A(n_403), .Y(n_908) );
INVx6_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g597 ( .A(n_404), .Y(n_597) );
INVx1_ASAP7_75t_L g631 ( .A(n_404), .Y(n_631) );
INVx1_ASAP7_75t_SL g668 ( .A(n_404), .Y(n_668) );
INVx1_ASAP7_75t_L g529 ( .A(n_405), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_422), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_417), .B2(n_418), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVx4_ASAP7_75t_L g506 ( .A(n_411), .Y(n_506) );
INVx4_ASAP7_75t_L g634 ( .A(n_411), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_411), .B(n_702), .Y(n_701) );
INVx3_ASAP7_75t_L g993 ( .A(n_411), .Y(n_993) );
INVx11_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx11_ASAP7_75t_L g561 ( .A(n_412), .Y(n_561) );
AND2x6_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g477 ( .A(n_414), .B(n_478), .Y(n_477) );
AND2x6_ASAP7_75t_L g457 ( .A(n_415), .B(n_450), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_418), .A2(n_819), .B1(n_820), .B2(n_821), .Y(n_818) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g675 ( .A(n_420), .Y(n_675) );
INVx2_ASAP7_75t_L g788 ( .A(n_420), .Y(n_788) );
INVx3_ASAP7_75t_L g845 ( .A(n_420), .Y(n_845) );
INVx6_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx3_ASAP7_75t_L g507 ( .A(n_421), .Y(n_507) );
BUFx3_ASAP7_75t_L g564 ( .A(n_421), .Y(n_564) );
BUFx3_ASAP7_75t_L g603 ( .A(n_421), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B1(n_427), .B2(n_428), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx2_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g493 ( .A(n_426), .Y(n_493) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_426), .Y(n_559) );
BUFx2_ASAP7_75t_SL g697 ( .A(n_426), .Y(n_697) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g821 ( .A(n_429), .Y(n_821) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx5_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g524 ( .A(n_434), .Y(n_524) );
INVx2_ASAP7_75t_L g550 ( .A(n_434), .Y(n_550) );
INVx4_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g881 ( .A(n_437), .Y(n_881) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
BUFx4f_ASAP7_75t_L g525 ( .A(n_438), .Y(n_525) );
BUFx2_ASAP7_75t_L g655 ( .A(n_438), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B1(n_446), .B2(n_447), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_441), .A2(n_776), .B1(n_777), .B2(n_779), .Y(n_775) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx3_ASAP7_75t_SL g583 ( .A(n_442), .Y(n_583) );
INVx4_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_443), .A2(n_448), .B1(n_488), .B2(n_489), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_443), .A2(n_585), .B1(n_613), .B2(n_614), .Y(n_612) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_443), .Y(n_750) );
OAI22xp33_ASAP7_75t_SL g810 ( .A1(n_443), .A2(n_752), .B1(n_811), .B2(n_812), .Y(n_810) );
BUFx3_ASAP7_75t_L g960 ( .A(n_443), .Y(n_960) );
NAND2x1p5_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
AND2x4_ASAP7_75t_L g459 ( .A(n_444), .B(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g464 ( .A(n_444), .B(n_465), .Y(n_464) );
AND2x4_ASAP7_75t_L g528 ( .A(n_444), .B(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
CKINVDCx16_ASAP7_75t_R g586 ( .A(n_448), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_448), .A2(n_583), .B1(n_987), .B2(n_988), .Y(n_986) );
OR2x6_ASAP7_75t_L g448 ( .A(n_449), .B(n_451), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g530 ( .A(n_450), .B(n_452), .Y(n_530) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g913 ( .A1(n_455), .A2(n_914), .B1(n_915), .B2(n_916), .C(n_917), .Y(n_913) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_456), .A2(n_712), .B(n_713), .Y(n_711) );
OAI21xp5_ASAP7_75t_SL g830 ( .A1(n_456), .A2(n_831), .B(n_832), .Y(n_830) );
OAI21xp5_ASAP7_75t_L g854 ( .A1(n_456), .A2(n_855), .B(n_856), .Y(n_854) );
OAI21xp5_ASAP7_75t_SL g876 ( .A1(n_456), .A2(n_877), .B(n_878), .Y(n_876) );
OAI22xp5_ASAP7_75t_SL g1061 ( .A1(n_456), .A2(n_1062), .B1(n_1063), .B2(n_1064), .Y(n_1061) );
INVx4_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g486 ( .A(n_457), .Y(n_486) );
INVx2_ASAP7_75t_L g545 ( .A(n_457), .Y(n_545) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_457), .Y(n_648) );
INVx2_ASAP7_75t_SL g955 ( .A(n_457), .Y(n_955) );
BUFx4f_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_459), .Y(n_484) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_459), .Y(n_535) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_459), .Y(n_618) );
BUFx2_ASAP7_75t_L g778 ( .A(n_459), .Y(n_778) );
INVx1_ASAP7_75t_L g465 ( .A(n_461), .Y(n_465) );
BUFx4f_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g809 ( .A(n_463), .Y(n_809) );
BUFx12f_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_464), .Y(n_580) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_464), .Y(n_621) );
INVx2_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND3x1_ASAP7_75t_L g472 ( .A(n_473), .B(n_490), .C(n_500), .Y(n_472) );
NOR3xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_482), .C(n_487), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B1(n_479), .B2(n_480), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_476), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_476), .A2(n_771), .B1(n_911), .B2(n_912), .Y(n_910) );
BUFx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_477), .Y(n_624) );
INVx2_ASAP7_75t_L g738 ( .A(n_477), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_477), .A2(n_769), .B1(n_770), .B2(n_771), .Y(n_768) );
BUFx3_ASAP7_75t_L g575 ( .A(n_480), .Y(n_575) );
INVx2_ASAP7_75t_L g741 ( .A(n_480), .Y(n_741) );
OAI22xp5_ASAP7_75t_SL g949 ( .A1(n_480), .A2(n_624), .B1(n_950), .B2(n_951), .Y(n_949) );
BUFx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g627 ( .A(n_481), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
INVx4_ASAP7_75t_L g652 ( .A(n_484), .Y(n_652) );
BUFx2_ASAP7_75t_L g807 ( .A(n_484), .Y(n_807) );
INVx2_ASAP7_75t_L g1063 ( .A(n_484), .Y(n_1063) );
INVx3_ASAP7_75t_L g532 ( .A(n_486), .Y(n_532) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_495), .Y(n_490) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx3_ASAP7_75t_L g785 ( .A(n_493), .Y(n_785) );
INVx1_ASAP7_75t_L g824 ( .A(n_494), .Y(n_824) );
BUFx2_ASAP7_75t_L g630 ( .A(n_496), .Y(n_630) );
BUFx6f_ASAP7_75t_L g907 ( .A(n_496), .Y(n_907) );
INVx5_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g518 ( .A(n_497), .Y(n_518) );
BUFx3_ASAP7_75t_L g596 ( .A(n_497), .Y(n_596) );
INVx3_ASAP7_75t_L g722 ( .A(n_497), .Y(n_722) );
INVx4_ASAP7_75t_L g759 ( .A(n_497), .Y(n_759) );
INVx8_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_505), .Y(n_500) );
BUFx2_ASAP7_75t_L g694 ( .A(n_502), .Y(n_694) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx3_ASAP7_75t_L g516 ( .A(n_503), .Y(n_516) );
BUFx3_ASAP7_75t_L g556 ( .A(n_503), .Y(n_556) );
BUFx3_ASAP7_75t_L g673 ( .A(n_503), .Y(n_673) );
INVx1_ASAP7_75t_L g604 ( .A(n_508), .Y(n_604) );
BUFx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AO22x1_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_536), .B2(n_537), .Y(n_510) );
INVx1_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
NOR4xp75_ASAP7_75t_L g513 ( .A(n_514), .B(n_519), .C(n_522), .D(n_531), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_515), .B(n_517), .Y(n_514) );
BUFx3_ASAP7_75t_L g903 ( .A(n_516), .Y(n_903) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_520), .B(n_521), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_523), .B(n_526), .Y(n_522) );
BUFx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g659 ( .A(n_528), .Y(n_659) );
BUFx2_ASAP7_75t_L g690 ( .A(n_528), .Y(n_690) );
BUFx2_ASAP7_75t_L g838 ( .A(n_528), .Y(n_838) );
BUFx3_ASAP7_75t_L g547 ( .A(n_530), .Y(n_547) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_530), .Y(n_662) );
BUFx2_ASAP7_75t_SL g833 ( .A(n_530), .Y(n_833) );
BUFx2_ASAP7_75t_SL g884 ( .A(n_530), .Y(n_884) );
OAI21xp5_ASAP7_75t_SL g531 ( .A1(n_532), .A2(n_533), .B(n_534), .Y(n_531) );
OAI21xp33_ASAP7_75t_L g772 ( .A1(n_532), .A2(n_773), .B(n_774), .Y(n_772) );
OAI21xp33_ASAP7_75t_SL g804 ( .A1(n_532), .A2(n_805), .B(n_806), .Y(n_804) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_535), .Y(n_687) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
XNOR2x1_ASAP7_75t_SL g537 ( .A(n_538), .B(n_569), .Y(n_537) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
XOR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_568), .Y(n_540) );
NAND2x1p5_ASAP7_75t_L g541 ( .A(n_542), .B(n_553), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_548), .Y(n_542) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_545), .B(n_546), .Y(n_543) );
OAI21xp33_ASAP7_75t_SL g576 ( .A1(n_545), .A2(n_577), .B(n_578), .Y(n_576) );
OAI21xp33_ASAP7_75t_L g615 ( .A1(n_545), .A2(n_616), .B(n_617), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g742 ( .A1(n_545), .A2(n_743), .B1(n_744), .B2(n_746), .C(n_747), .Y(n_742) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_551), .C(n_552), .Y(n_548) );
NOR2x1_ASAP7_75t_L g553 ( .A(n_554), .B(n_562), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_558), .Y(n_554) );
INVx3_ASAP7_75t_L g591 ( .A(n_559), .Y(n_591) );
BUFx6f_ASAP7_75t_L g671 ( .A(n_559), .Y(n_671) );
BUFx3_ASAP7_75t_L g902 ( .A(n_559), .Y(n_902) );
BUFx3_ASAP7_75t_L g966 ( .A(n_559), .Y(n_966) );
INVx5_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_SL g720 ( .A(n_561), .Y(n_720) );
INVx4_ASAP7_75t_L g783 ( .A(n_561), .Y(n_783) );
INVx2_ASAP7_75t_L g816 ( .A(n_561), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx4_ASAP7_75t_L g593 ( .A(n_566), .Y(n_593) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_587), .Y(n_570) );
NOR3xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_576), .C(n_581), .Y(n_571) );
OAI22xp5_ASAP7_75t_SL g799 ( .A1(n_575), .A2(n_800), .B1(n_802), .B2(n_803), .Y(n_799) );
INVx1_ASAP7_75t_L g957 ( .A(n_579), .Y(n_957) );
BUFx4f_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .B1(n_584), .B2(n_585), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_583), .A2(n_752), .B1(n_920), .B2(n_921), .Y(n_919) );
OAI22xp5_ASAP7_75t_SL g1055 ( .A1(n_583), .A2(n_626), .B1(n_1056), .B2(n_1057), .Y(n_1055) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g752 ( .A(n_586), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_598), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_594), .Y(n_588) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx4_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx3_ASAP7_75t_L g665 ( .A(n_593), .Y(n_665) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_601), .A2(n_823), .B1(n_824), .B2(n_825), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_728), .B1(n_868), .B2(n_869), .Y(n_605) );
INVx1_ASAP7_75t_L g868 ( .A(n_606), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_679), .B1(n_726), .B2(n_727), .Y(n_606) );
INVx1_ASAP7_75t_L g726 ( .A(n_607), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_640), .B1(n_677), .B2(n_678), .Y(n_607) );
INVx1_ASAP7_75t_L g677 ( .A(n_608), .Y(n_677) );
INVx2_ASAP7_75t_L g639 ( .A(n_610), .Y(n_639) );
NAND2x1_ASAP7_75t_L g610 ( .A(n_611), .B(n_628), .Y(n_610) );
NOR3xp33_ASAP7_75t_SL g611 ( .A(n_612), .B(n_615), .C(n_622), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g915 ( .A(n_618), .Y(n_915) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
BUFx3_ASAP7_75t_L g745 ( .A(n_621), .Y(n_745) );
BUFx2_ASAP7_75t_L g918 ( .A(n_621), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B1(n_625), .B2(n_626), .Y(n_622) );
INVx1_ASAP7_75t_L g801 ( .A(n_624), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_624), .A2(n_626), .B1(n_981), .B2(n_982), .Y(n_980) );
OAI21xp5_ASAP7_75t_SL g1058 ( .A1(n_624), .A2(n_1059), .B(n_1060), .Y(n_1058) );
OA211x2_ASAP7_75t_L g933 ( .A1(n_626), .A2(n_934), .B(n_935), .C(n_936), .Y(n_933) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g771 ( .A(n_627), .Y(n_771) );
AND4x1_ASAP7_75t_L g628 ( .A(n_629), .B(n_632), .C(n_633), .D(n_636), .Y(n_628) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g678 ( .A(n_640), .Y(n_678) );
BUFx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g676 ( .A(n_644), .Y(n_676) );
NAND3x1_ASAP7_75t_L g644 ( .A(n_645), .B(n_663), .C(n_669), .Y(n_644) );
NOR2x1_ASAP7_75t_L g645 ( .A(n_646), .B(n_653), .Y(n_645) );
OAI21xp5_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_649), .B(n_650), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g684 ( .A1(n_647), .A2(n_685), .B(n_686), .Y(n_684) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx3_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .C(n_657), .Y(n_653) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g1032 ( .A(n_659), .Y(n_1032) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_667), .Y(n_663) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_674), .Y(n_669) );
BUFx4f_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g974 ( .A(n_673), .Y(n_974) );
INVx1_ASAP7_75t_L g727 ( .A(n_679), .Y(n_727) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
OAI22x1_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_703), .B1(n_724), .B2(n_725), .Y(n_680) );
INVx1_ASAP7_75t_L g724 ( .A(n_681), .Y(n_724) );
NAND3x1_ASAP7_75t_L g682 ( .A(n_683), .B(n_692), .C(n_696), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_688), .Y(n_683) );
INVx2_ASAP7_75t_SL g953 ( .A(n_687), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g725 ( .A(n_703), .Y(n_725) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
XOR2x2_ASAP7_75t_L g764 ( .A(n_704), .B(n_765), .Y(n_764) );
XOR2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_723), .Y(n_704) );
NAND3x1_ASAP7_75t_L g705 ( .A(n_706), .B(n_710), .C(n_718), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
BUFx2_ASAP7_75t_L g762 ( .A(n_709), .Y(n_762) );
NOR2x1_ASAP7_75t_L g710 ( .A(n_711), .B(n_714), .Y(n_710) );
NAND3xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .C(n_717), .Y(n_714) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_721), .Y(n_718) );
INVx1_ASAP7_75t_L g869 ( .A(n_728), .Y(n_869) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_793), .B1(n_866), .B2(n_867), .Y(n_730) );
INVx2_ASAP7_75t_L g866 ( .A(n_731), .Y(n_866) );
OA22x2_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_764), .B1(n_791), .B2(n_792), .Y(n_731) );
INVx2_ASAP7_75t_L g791 ( .A(n_732), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_753), .Y(n_733) );
NOR3xp33_ASAP7_75t_L g734 ( .A(n_735), .B(n_742), .C(n_748), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B1(n_739), .B2(n_740), .Y(n_735) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B1(n_751), .B2(n_752), .Y(n_748) );
OAI22xp5_ASAP7_75t_SL g959 ( .A1(n_752), .A2(n_960), .B1(n_961), .B2(n_962), .Y(n_959) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_760), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_757), .Y(n_754) );
BUFx6f_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
BUFx2_ASAP7_75t_L g888 ( .A(n_759), .Y(n_888) );
INVx2_ASAP7_75t_L g969 ( .A(n_759), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_763), .Y(n_760) );
INVx2_ASAP7_75t_L g792 ( .A(n_764), .Y(n_792) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_780), .Y(n_766) );
NOR3xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_772), .C(n_775), .Y(n_767) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_786), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_784), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_789), .Y(n_786) );
INVx1_ASAP7_75t_L g867 ( .A(n_793), .Y(n_867) );
XNOR2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_826), .Y(n_793) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_813), .Y(n_797) );
NOR3xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_804), .C(n_810), .Y(n_798) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx3_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
NOR3xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_818), .C(n_822), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_817), .Y(n_814) );
OAI22x1_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_847), .B1(n_848), .B2(n_865), .Y(n_826) );
INVx2_ASAP7_75t_L g865 ( .A(n_827), .Y(n_865) );
AND2x4_ASAP7_75t_L g828 ( .A(n_829), .B(n_839), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_834), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g834 ( .A(n_835), .B(n_836), .C(n_837), .Y(n_834) );
NOR2x1_ASAP7_75t_L g839 ( .A(n_840), .B(n_843), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_841), .B(n_842), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_844), .B(n_846), .Y(n_843) );
INVx3_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
XOR2x2_ASAP7_75t_L g848 ( .A(n_849), .B(n_864), .Y(n_848) );
NAND3x1_ASAP7_75t_SL g849 ( .A(n_850), .B(n_853), .C(n_861), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
NOR2x1_ASAP7_75t_L g853 ( .A(n_854), .B(n_857), .Y(n_853) );
NAND3xp33_ASAP7_75t_L g857 ( .A(n_858), .B(n_859), .C(n_860), .Y(n_857) );
AND2x2_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
INVx1_ASAP7_75t_L g1005 ( .A(n_870), .Y(n_1005) );
AOI22xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B1(n_893), .B2(n_1003), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
XOR2x2_ASAP7_75t_L g873 ( .A(n_874), .B(n_892), .Y(n_873) );
NAND3x1_ASAP7_75t_L g874 ( .A(n_875), .B(n_885), .C(n_889), .Y(n_874) );
NOR2x1_ASAP7_75t_L g875 ( .A(n_876), .B(n_879), .Y(n_875) );
NAND3xp33_ASAP7_75t_L g879 ( .A(n_880), .B(n_882), .C(n_883), .Y(n_879) );
AND2x2_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
AND2x2_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
INVx1_ASAP7_75t_L g1003 ( .A(n_893), .Y(n_1003) );
AOI22xp5_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_943), .B1(n_1001), .B2(n_1002), .Y(n_893) );
INVx1_ASAP7_75t_L g1001 ( .A(n_894), .Y(n_1001) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g895 ( .A1(n_896), .A2(n_924), .B1(n_925), .B2(n_942), .Y(n_895) );
INVx1_ASAP7_75t_L g942 ( .A(n_896), .Y(n_942) );
INVx1_ASAP7_75t_SL g923 ( .A(n_897), .Y(n_923) );
AND2x2_ASAP7_75t_SL g897 ( .A(n_898), .B(n_909), .Y(n_897) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_904), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_905), .B(n_906), .Y(n_904) );
NOR3xp33_ASAP7_75t_L g909 ( .A(n_910), .B(n_913), .C(n_919), .Y(n_909) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
AO22x1_ASAP7_75t_L g976 ( .A1(n_926), .A2(n_927), .B1(n_977), .B2(n_999), .Y(n_976) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
XOR2x2_ASAP7_75t_L g927 ( .A(n_928), .B(n_941), .Y(n_927) );
NAND4xp75_ASAP7_75t_L g928 ( .A(n_929), .B(n_933), .C(n_937), .D(n_940), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_930), .B(n_932), .Y(n_929) );
AND2x2_ASAP7_75t_L g937 ( .A(n_938), .B(n_939), .Y(n_937) );
INVx2_ASAP7_75t_L g1002 ( .A(n_943), .Y(n_1002) );
BUFx2_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
AOI22xp5_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_975), .B1(n_976), .B2(n_1000), .Y(n_944) );
INVx2_ASAP7_75t_L g1000 ( .A(n_945), .Y(n_1000) );
XNOR2x2_ASAP7_75t_L g945 ( .A(n_946), .B(n_947), .Y(n_945) );
AND2x2_ASAP7_75t_L g947 ( .A(n_948), .B(n_963), .Y(n_947) );
NOR3xp33_ASAP7_75t_L g948 ( .A(n_949), .B(n_952), .C(n_959), .Y(n_948) );
OAI222xp33_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_954), .B1(n_955), .B2(n_956), .C1(n_957), .C2(n_958), .Y(n_952) );
OAI21xp5_ASAP7_75t_SL g983 ( .A1(n_955), .A2(n_984), .B(n_985), .Y(n_983) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_964), .B(n_970), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_965), .B(n_967), .Y(n_964) );
INVx3_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_971), .B(n_972), .Y(n_970) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
INVx1_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g999 ( .A(n_977), .Y(n_999) );
INVx2_ASAP7_75t_L g997 ( .A(n_978), .Y(n_997) );
AND2x2_ASAP7_75t_L g978 ( .A(n_979), .B(n_989), .Y(n_978) );
NOR3xp33_ASAP7_75t_L g979 ( .A(n_980), .B(n_983), .C(n_986), .Y(n_979) );
NOR2xp33_ASAP7_75t_L g989 ( .A(n_990), .B(n_994), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_991), .B(n_992), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_995), .B(n_996), .Y(n_994) );
INVx1_ASAP7_75t_SL g1006 ( .A(n_1007), .Y(n_1006) );
NOR2x1_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1012), .Y(n_1007) );
OR2x2_ASAP7_75t_SL g1067 ( .A(n_1008), .B(n_1013), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1011), .Y(n_1008) );
CKINVDCx20_ASAP7_75t_R g1037 ( .A(n_1009), .Y(n_1037) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_1010), .B(n_1039), .Y(n_1042) );
CKINVDCx16_ASAP7_75t_R g1039 ( .A(n_1011), .Y(n_1039) );
CKINVDCx20_ASAP7_75t_R g1012 ( .A(n_1013), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1015), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_1017), .B(n_1018), .Y(n_1016) );
OAI322xp33_ASAP7_75t_L g1019 ( .A1(n_1020), .A2(n_1035), .A3(n_1038), .B1(n_1040), .B2(n_1043), .C1(n_1044), .C2(n_1065), .Y(n_1019) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
NAND4xp75_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1026), .C(n_1029), .D(n_1033), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1025), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1028), .Y(n_1026) );
AND2x2_ASAP7_75t_SL g1029 ( .A(n_1030), .B(n_1031), .Y(n_1029) );
HB1xp67_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
HB1xp67_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
CKINVDCx16_ASAP7_75t_R g1040 ( .A(n_1041), .Y(n_1040) );
XNOR2xp5_ASAP7_75t_L g1046 ( .A(n_1043), .B(n_1047), .Y(n_1046) );
INVx1_ASAP7_75t_SL g1044 ( .A(n_1045), .Y(n_1044) );
HB1xp67_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
NAND3x1_ASAP7_75t_SL g1047 ( .A(n_1048), .B(n_1051), .C(n_1054), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1050), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1053), .Y(n_1051) );
NOR3xp33_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1058), .C(n_1061), .Y(n_1054) );
CKINVDCx20_ASAP7_75t_R g1065 ( .A(n_1066), .Y(n_1065) );
CKINVDCx20_ASAP7_75t_R g1066 ( .A(n_1067), .Y(n_1066) );
endmodule